module mux_aoi_ready_valid_const_21_17 (
	I,
	S,
	ready_in,
	ready_out,
	valid_in,
	valid_out,
	out_sel,
	O
);
	input wire [356:0] I;
	input wire [4:0] S;
	input wire ready_in;
	output wire ready_out;
	input wire [20:0] valid_in;
	output wire valid_out;
	output wire [31:0] out_sel;
	output wire [16:0] O;
	wire [16:0] O_int0;
	wire [16:0] O_int1;
	wire [16:0] O_int2;
	wire [16:0] O_int3;
	wire [16:0] O_int4;
	wire [16:0] O_int5;
	wire [16:0] O_int6;
	wire [16:0] O_int7;
	wire [16:0] O_int8;
	wire [16:0] O_int9;
	wire [16:0] O_int10;
	wire [10:0] valid_out_temp;
	precoder_17_21 u_precoder(
		.S(S),
		.out_sel(out_sel)
	);
	mux_logic_17_21 u_mux_logic(
		.I0(I[0+:17]),
		.I1(I[17+:17]),
		.I2(I[34+:17]),
		.I3(I[51+:17]),
		.I4(I[68+:17]),
		.I5(I[85+:17]),
		.I6(I[102+:17]),
		.I7(I[119+:17]),
		.I8(I[136+:17]),
		.I9(I[153+:17]),
		.I10(I[170+:17]),
		.I11(I[187+:17]),
		.I12(I[204+:17]),
		.I13(I[221+:17]),
		.I14(I[238+:17]),
		.I15(I[255+:17]),
		.I16(I[272+:17]),
		.I17(I[289+:17]),
		.I18(I[306+:17]),
		.I19(I[323+:17]),
		.I20(I[340+:17]),
		.out_sel(out_sel),
		.valid_in(valid_in),
		.valid_out(valid_out_temp),
		.O0(O_int0),
		.O1(O_int1),
		.O2(O_int2),
		.O3(O_int3),
		.O4(O_int4),
		.O5(O_int5),
		.O6(O_int6),
		.O7(O_int7),
		.O8(O_int8),
		.O9(O_int9),
		.O10(O_int10)
	);
	assign O = (((((((((O_int0 | O_int1) | O_int2) | O_int3) | O_int4) | O_int5) | O_int6) | O_int7) | O_int8) | O_int9) | O_int10;
	assign ready_out = ready_in;
	assign valid_out = |valid_out_temp;
endmodule
module precoder_17_21 (
	S,
	out_sel
);
	input wire [4:0] S;
	output reg [31:0] out_sel;
	always @(*) begin : mux_sel
		case (S)
			5'd0: out_sel = 32'b00000000000000000000000000000001;
			5'd1: out_sel = 32'b00000000000000000000000000000010;
			5'd2: out_sel = 32'b00000000000000000000000000000100;
			5'd3: out_sel = 32'b00000000000000000000000000001000;
			5'd4: out_sel = 32'b00000000000000000000000000010000;
			5'd5: out_sel = 32'b00000000000000000000000000100000;
			5'd6: out_sel = 32'b00000000000000000000000001000000;
			5'd7: out_sel = 32'b00000000000000000000000010000000;
			5'd8: out_sel = 32'b00000000000000000000000100000000;
			5'd9: out_sel = 32'b00000000000000000000001000000000;
			5'd10: out_sel = 32'b00000000000000000000010000000000;
			5'd11: out_sel = 32'b00000000000000000000100000000000;
			5'd12: out_sel = 32'b00000000000000000001000000000000;
			5'd13: out_sel = 32'b00000000000000000010000000000000;
			5'd14: out_sel = 32'b00000000000000000100000000000000;
			5'd15: out_sel = 32'b00000000000000001000000000000000;
			5'd16: out_sel = 32'b00000000000000010000000000000000;
			5'd17: out_sel = 32'b00000000000000100000000000000000;
			5'd18: out_sel = 32'b00000000000001000000000000000000;
			5'd19: out_sel = 32'b00000000000010000000000000000000;
			5'd20: out_sel = 32'b00000000000100000000000000000000;
			5'd21: out_sel = 32'b00000000001000000000000000000000;
			default: out_sel = 32'b00000000000000000000000000000000;
		endcase
	end
endmodule
module mux_logic_17_21 (
	out_sel,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	I9,
	I10,
	I11,
	I12,
	I13,
	I14,
	I15,
	I16,
	I17,
	I18,
	I19,
	I20,
	valid_in,
	valid_out,
	O0,
	O1,
	O2,
	O3,
	O4,
	O5,
	O6,
	O7,
	O8,
	O9,
	O10
);
	input wire [31:0] out_sel;
	input wire [16:0] I0;
	input wire [16:0] I1;
	input wire [16:0] I2;
	input wire [16:0] I3;
	input wire [16:0] I4;
	input wire [16:0] I5;
	input wire [16:0] I6;
	input wire [16:0] I7;
	input wire [16:0] I8;
	input wire [16:0] I9;
	input wire [16:0] I10;
	input wire [16:0] I11;
	input wire [16:0] I12;
	input wire [16:0] I13;
	input wire [16:0] I14;
	input wire [16:0] I15;
	input wire [16:0] I16;
	input wire [16:0] I17;
	input wire [16:0] I18;
	input wire [16:0] I19;
	input wire [16:0] I20;
	input wire [20:0] valid_in;
	output wire [10:0] valid_out;
	output wire [16:0] O0;
	output wire [16:0] O1;
	output wire [16:0] O2;
	output wire [16:0] O3;
	output wire [16:0] O4;
	output wire [16:0] O5;
	output wire [16:0] O6;
	output wire [16:0] O7;
	output wire [16:0] O8;
	output wire [16:0] O9;
	output wire [16:0] O10;
	AO_CELL inst_0_0(
		.A1(out_sel[0]),
		.A2(I0[0]),
		.B1(out_sel[1]),
		.B2(I1[0]),
		.Z(O0[0])
	);
	AO_CELL inst_1_0(
		.A1(out_sel[2]),
		.A2(I2[0]),
		.B1(out_sel[3]),
		.B2(I3[0]),
		.Z(O1[0])
	);
	AO_CELL inst_2_0(
		.A1(out_sel[4]),
		.A2(I4[0]),
		.B1(out_sel[5]),
		.B2(I5[0]),
		.Z(O2[0])
	);
	AO_CELL inst_3_0(
		.A1(out_sel[6]),
		.A2(I6[0]),
		.B1(out_sel[7]),
		.B2(I7[0]),
		.Z(O3[0])
	);
	AO_CELL inst_4_0(
		.A1(out_sel[8]),
		.A2(I8[0]),
		.B1(out_sel[9]),
		.B2(I9[0]),
		.Z(O4[0])
	);
	AO_CELL inst_5_0(
		.A1(out_sel[10]),
		.A2(I10[0]),
		.B1(out_sel[11]),
		.B2(I11[0]),
		.Z(O5[0])
	);
	AO_CELL inst_6_0(
		.A1(out_sel[12]),
		.A2(I12[0]),
		.B1(out_sel[13]),
		.B2(I13[0]),
		.Z(O6[0])
	);
	AO_CELL inst_7_0(
		.A1(out_sel[14]),
		.A2(I14[0]),
		.B1(out_sel[15]),
		.B2(I15[0]),
		.Z(O7[0])
	);
	AO_CELL inst_8_0(
		.A1(out_sel[16]),
		.A2(I16[0]),
		.B1(out_sel[17]),
		.B2(I17[0]),
		.Z(O8[0])
	);
	AO_CELL inst_9_0(
		.A1(out_sel[18]),
		.A2(I18[0]),
		.B1(out_sel[19]),
		.B2(I19[0]),
		.Z(O9[0])
	);
	AO_CELL inst_10_0(
		.A1(out_sel[20]),
		.A2(I20[0]),
		.B1(out_sel[21]),
		.B2(1'b0),
		.Z(O10[0])
	);
	AO_CELL inst_0_1(
		.A1(out_sel[0]),
		.A2(I0[1]),
		.B1(out_sel[1]),
		.B2(I1[1]),
		.Z(O0[1])
	);
	AO_CELL inst_1_1(
		.A1(out_sel[2]),
		.A2(I2[1]),
		.B1(out_sel[3]),
		.B2(I3[1]),
		.Z(O1[1])
	);
	AO_CELL inst_2_1(
		.A1(out_sel[4]),
		.A2(I4[1]),
		.B1(out_sel[5]),
		.B2(I5[1]),
		.Z(O2[1])
	);
	AO_CELL inst_3_1(
		.A1(out_sel[6]),
		.A2(I6[1]),
		.B1(out_sel[7]),
		.B2(I7[1]),
		.Z(O3[1])
	);
	AO_CELL inst_4_1(
		.A1(out_sel[8]),
		.A2(I8[1]),
		.B1(out_sel[9]),
		.B2(I9[1]),
		.Z(O4[1])
	);
	AO_CELL inst_5_1(
		.A1(out_sel[10]),
		.A2(I10[1]),
		.B1(out_sel[11]),
		.B2(I11[1]),
		.Z(O5[1])
	);
	AO_CELL inst_6_1(
		.A1(out_sel[12]),
		.A2(I12[1]),
		.B1(out_sel[13]),
		.B2(I13[1]),
		.Z(O6[1])
	);
	AO_CELL inst_7_1(
		.A1(out_sel[14]),
		.A2(I14[1]),
		.B1(out_sel[15]),
		.B2(I15[1]),
		.Z(O7[1])
	);
	AO_CELL inst_8_1(
		.A1(out_sel[16]),
		.A2(I16[1]),
		.B1(out_sel[17]),
		.B2(I17[1]),
		.Z(O8[1])
	);
	AO_CELL inst_9_1(
		.A1(out_sel[18]),
		.A2(I18[1]),
		.B1(out_sel[19]),
		.B2(I19[1]),
		.Z(O9[1])
	);
	AO_CELL inst_10_1(
		.A1(out_sel[20]),
		.A2(I20[1]),
		.B1(out_sel[21]),
		.B2(1'b0),
		.Z(O10[1])
	);
	AO_CELL inst_0_2(
		.A1(out_sel[0]),
		.A2(I0[2]),
		.B1(out_sel[1]),
		.B2(I1[2]),
		.Z(O0[2])
	);
	AO_CELL inst_1_2(
		.A1(out_sel[2]),
		.A2(I2[2]),
		.B1(out_sel[3]),
		.B2(I3[2]),
		.Z(O1[2])
	);
	AO_CELL inst_2_2(
		.A1(out_sel[4]),
		.A2(I4[2]),
		.B1(out_sel[5]),
		.B2(I5[2]),
		.Z(O2[2])
	);
	AO_CELL inst_3_2(
		.A1(out_sel[6]),
		.A2(I6[2]),
		.B1(out_sel[7]),
		.B2(I7[2]),
		.Z(O3[2])
	);
	AO_CELL inst_4_2(
		.A1(out_sel[8]),
		.A2(I8[2]),
		.B1(out_sel[9]),
		.B2(I9[2]),
		.Z(O4[2])
	);
	AO_CELL inst_5_2(
		.A1(out_sel[10]),
		.A2(I10[2]),
		.B1(out_sel[11]),
		.B2(I11[2]),
		.Z(O5[2])
	);
	AO_CELL inst_6_2(
		.A1(out_sel[12]),
		.A2(I12[2]),
		.B1(out_sel[13]),
		.B2(I13[2]),
		.Z(O6[2])
	);
	AO_CELL inst_7_2(
		.A1(out_sel[14]),
		.A2(I14[2]),
		.B1(out_sel[15]),
		.B2(I15[2]),
		.Z(O7[2])
	);
	AO_CELL inst_8_2(
		.A1(out_sel[16]),
		.A2(I16[2]),
		.B1(out_sel[17]),
		.B2(I17[2]),
		.Z(O8[2])
	);
	AO_CELL inst_9_2(
		.A1(out_sel[18]),
		.A2(I18[2]),
		.B1(out_sel[19]),
		.B2(I19[2]),
		.Z(O9[2])
	);
	AO_CELL inst_10_2(
		.A1(out_sel[20]),
		.A2(I20[2]),
		.B1(out_sel[21]),
		.B2(1'b0),
		.Z(O10[2])
	);
	AO_CELL inst_0_3(
		.A1(out_sel[0]),
		.A2(I0[3]),
		.B1(out_sel[1]),
		.B2(I1[3]),
		.Z(O0[3])
	);
	AO_CELL inst_1_3(
		.A1(out_sel[2]),
		.A2(I2[3]),
		.B1(out_sel[3]),
		.B2(I3[3]),
		.Z(O1[3])
	);
	AO_CELL inst_2_3(
		.A1(out_sel[4]),
		.A2(I4[3]),
		.B1(out_sel[5]),
		.B2(I5[3]),
		.Z(O2[3])
	);
	AO_CELL inst_3_3(
		.A1(out_sel[6]),
		.A2(I6[3]),
		.B1(out_sel[7]),
		.B2(I7[3]),
		.Z(O3[3])
	);
	AO_CELL inst_4_3(
		.A1(out_sel[8]),
		.A2(I8[3]),
		.B1(out_sel[9]),
		.B2(I9[3]),
		.Z(O4[3])
	);
	AO_CELL inst_5_3(
		.A1(out_sel[10]),
		.A2(I10[3]),
		.B1(out_sel[11]),
		.B2(I11[3]),
		.Z(O5[3])
	);
	AO_CELL inst_6_3(
		.A1(out_sel[12]),
		.A2(I12[3]),
		.B1(out_sel[13]),
		.B2(I13[3]),
		.Z(O6[3])
	);
	AO_CELL inst_7_3(
		.A1(out_sel[14]),
		.A2(I14[3]),
		.B1(out_sel[15]),
		.B2(I15[3]),
		.Z(O7[3])
	);
	AO_CELL inst_8_3(
		.A1(out_sel[16]),
		.A2(I16[3]),
		.B1(out_sel[17]),
		.B2(I17[3]),
		.Z(O8[3])
	);
	AO_CELL inst_9_3(
		.A1(out_sel[18]),
		.A2(I18[3]),
		.B1(out_sel[19]),
		.B2(I19[3]),
		.Z(O9[3])
	);
	AO_CELL inst_10_3(
		.A1(out_sel[20]),
		.A2(I20[3]),
		.B1(out_sel[21]),
		.B2(1'b0),
		.Z(O10[3])
	);
	AO_CELL inst_0_4(
		.A1(out_sel[0]),
		.A2(I0[4]),
		.B1(out_sel[1]),
		.B2(I1[4]),
		.Z(O0[4])
	);
	AO_CELL inst_1_4(
		.A1(out_sel[2]),
		.A2(I2[4]),
		.B1(out_sel[3]),
		.B2(I3[4]),
		.Z(O1[4])
	);
	AO_CELL inst_2_4(
		.A1(out_sel[4]),
		.A2(I4[4]),
		.B1(out_sel[5]),
		.B2(I5[4]),
		.Z(O2[4])
	);
	AO_CELL inst_3_4(
		.A1(out_sel[6]),
		.A2(I6[4]),
		.B1(out_sel[7]),
		.B2(I7[4]),
		.Z(O3[4])
	);
	AO_CELL inst_4_4(
		.A1(out_sel[8]),
		.A2(I8[4]),
		.B1(out_sel[9]),
		.B2(I9[4]),
		.Z(O4[4])
	);
	AO_CELL inst_5_4(
		.A1(out_sel[10]),
		.A2(I10[4]),
		.B1(out_sel[11]),
		.B2(I11[4]),
		.Z(O5[4])
	);
	AO_CELL inst_6_4(
		.A1(out_sel[12]),
		.A2(I12[4]),
		.B1(out_sel[13]),
		.B2(I13[4]),
		.Z(O6[4])
	);
	AO_CELL inst_7_4(
		.A1(out_sel[14]),
		.A2(I14[4]),
		.B1(out_sel[15]),
		.B2(I15[4]),
		.Z(O7[4])
	);
	AO_CELL inst_8_4(
		.A1(out_sel[16]),
		.A2(I16[4]),
		.B1(out_sel[17]),
		.B2(I17[4]),
		.Z(O8[4])
	);
	AO_CELL inst_9_4(
		.A1(out_sel[18]),
		.A2(I18[4]),
		.B1(out_sel[19]),
		.B2(I19[4]),
		.Z(O9[4])
	);
	AO_CELL inst_10_4(
		.A1(out_sel[20]),
		.A2(I20[4]),
		.B1(out_sel[21]),
		.B2(1'b0),
		.Z(O10[4])
	);
	AO_CELL inst_0_5(
		.A1(out_sel[0]),
		.A2(I0[5]),
		.B1(out_sel[1]),
		.B2(I1[5]),
		.Z(O0[5])
	);
	AO_CELL inst_1_5(
		.A1(out_sel[2]),
		.A2(I2[5]),
		.B1(out_sel[3]),
		.B2(I3[5]),
		.Z(O1[5])
	);
	AO_CELL inst_2_5(
		.A1(out_sel[4]),
		.A2(I4[5]),
		.B1(out_sel[5]),
		.B2(I5[5]),
		.Z(O2[5])
	);
	AO_CELL inst_3_5(
		.A1(out_sel[6]),
		.A2(I6[5]),
		.B1(out_sel[7]),
		.B2(I7[5]),
		.Z(O3[5])
	);
	AO_CELL inst_4_5(
		.A1(out_sel[8]),
		.A2(I8[5]),
		.B1(out_sel[9]),
		.B2(I9[5]),
		.Z(O4[5])
	);
	AO_CELL inst_5_5(
		.A1(out_sel[10]),
		.A2(I10[5]),
		.B1(out_sel[11]),
		.B2(I11[5]),
		.Z(O5[5])
	);
	AO_CELL inst_6_5(
		.A1(out_sel[12]),
		.A2(I12[5]),
		.B1(out_sel[13]),
		.B2(I13[5]),
		.Z(O6[5])
	);
	AO_CELL inst_7_5(
		.A1(out_sel[14]),
		.A2(I14[5]),
		.B1(out_sel[15]),
		.B2(I15[5]),
		.Z(O7[5])
	);
	AO_CELL inst_8_5(
		.A1(out_sel[16]),
		.A2(I16[5]),
		.B1(out_sel[17]),
		.B2(I17[5]),
		.Z(O8[5])
	);
	AO_CELL inst_9_5(
		.A1(out_sel[18]),
		.A2(I18[5]),
		.B1(out_sel[19]),
		.B2(I19[5]),
		.Z(O9[5])
	);
	AO_CELL inst_10_5(
		.A1(out_sel[20]),
		.A2(I20[5]),
		.B1(out_sel[21]),
		.B2(1'b0),
		.Z(O10[5])
	);
	AO_CELL inst_0_6(
		.A1(out_sel[0]),
		.A2(I0[6]),
		.B1(out_sel[1]),
		.B2(I1[6]),
		.Z(O0[6])
	);
	AO_CELL inst_1_6(
		.A1(out_sel[2]),
		.A2(I2[6]),
		.B1(out_sel[3]),
		.B2(I3[6]),
		.Z(O1[6])
	);
	AO_CELL inst_2_6(
		.A1(out_sel[4]),
		.A2(I4[6]),
		.B1(out_sel[5]),
		.B2(I5[6]),
		.Z(O2[6])
	);
	AO_CELL inst_3_6(
		.A1(out_sel[6]),
		.A2(I6[6]),
		.B1(out_sel[7]),
		.B2(I7[6]),
		.Z(O3[6])
	);
	AO_CELL inst_4_6(
		.A1(out_sel[8]),
		.A2(I8[6]),
		.B1(out_sel[9]),
		.B2(I9[6]),
		.Z(O4[6])
	);
	AO_CELL inst_5_6(
		.A1(out_sel[10]),
		.A2(I10[6]),
		.B1(out_sel[11]),
		.B2(I11[6]),
		.Z(O5[6])
	);
	AO_CELL inst_6_6(
		.A1(out_sel[12]),
		.A2(I12[6]),
		.B1(out_sel[13]),
		.B2(I13[6]),
		.Z(O6[6])
	);
	AO_CELL inst_7_6(
		.A1(out_sel[14]),
		.A2(I14[6]),
		.B1(out_sel[15]),
		.B2(I15[6]),
		.Z(O7[6])
	);
	AO_CELL inst_8_6(
		.A1(out_sel[16]),
		.A2(I16[6]),
		.B1(out_sel[17]),
		.B2(I17[6]),
		.Z(O8[6])
	);
	AO_CELL inst_9_6(
		.A1(out_sel[18]),
		.A2(I18[6]),
		.B1(out_sel[19]),
		.B2(I19[6]),
		.Z(O9[6])
	);
	AO_CELL inst_10_6(
		.A1(out_sel[20]),
		.A2(I20[6]),
		.B1(out_sel[21]),
		.B2(1'b0),
		.Z(O10[6])
	);
	AO_CELL inst_0_7(
		.A1(out_sel[0]),
		.A2(I0[7]),
		.B1(out_sel[1]),
		.B2(I1[7]),
		.Z(O0[7])
	);
	AO_CELL inst_1_7(
		.A1(out_sel[2]),
		.A2(I2[7]),
		.B1(out_sel[3]),
		.B2(I3[7]),
		.Z(O1[7])
	);
	AO_CELL inst_2_7(
		.A1(out_sel[4]),
		.A2(I4[7]),
		.B1(out_sel[5]),
		.B2(I5[7]),
		.Z(O2[7])
	);
	AO_CELL inst_3_7(
		.A1(out_sel[6]),
		.A2(I6[7]),
		.B1(out_sel[7]),
		.B2(I7[7]),
		.Z(O3[7])
	);
	AO_CELL inst_4_7(
		.A1(out_sel[8]),
		.A2(I8[7]),
		.B1(out_sel[9]),
		.B2(I9[7]),
		.Z(O4[7])
	);
	AO_CELL inst_5_7(
		.A1(out_sel[10]),
		.A2(I10[7]),
		.B1(out_sel[11]),
		.B2(I11[7]),
		.Z(O5[7])
	);
	AO_CELL inst_6_7(
		.A1(out_sel[12]),
		.A2(I12[7]),
		.B1(out_sel[13]),
		.B2(I13[7]),
		.Z(O6[7])
	);
	AO_CELL inst_7_7(
		.A1(out_sel[14]),
		.A2(I14[7]),
		.B1(out_sel[15]),
		.B2(I15[7]),
		.Z(O7[7])
	);
	AO_CELL inst_8_7(
		.A1(out_sel[16]),
		.A2(I16[7]),
		.B1(out_sel[17]),
		.B2(I17[7]),
		.Z(O8[7])
	);
	AO_CELL inst_9_7(
		.A1(out_sel[18]),
		.A2(I18[7]),
		.B1(out_sel[19]),
		.B2(I19[7]),
		.Z(O9[7])
	);
	AO_CELL inst_10_7(
		.A1(out_sel[20]),
		.A2(I20[7]),
		.B1(out_sel[21]),
		.B2(1'b0),
		.Z(O10[7])
	);
	AO_CELL inst_0_8(
		.A1(out_sel[0]),
		.A2(I0[8]),
		.B1(out_sel[1]),
		.B2(I1[8]),
		.Z(O0[8])
	);
	AO_CELL inst_1_8(
		.A1(out_sel[2]),
		.A2(I2[8]),
		.B1(out_sel[3]),
		.B2(I3[8]),
		.Z(O1[8])
	);
	AO_CELL inst_2_8(
		.A1(out_sel[4]),
		.A2(I4[8]),
		.B1(out_sel[5]),
		.B2(I5[8]),
		.Z(O2[8])
	);
	AO_CELL inst_3_8(
		.A1(out_sel[6]),
		.A2(I6[8]),
		.B1(out_sel[7]),
		.B2(I7[8]),
		.Z(O3[8])
	);
	AO_CELL inst_4_8(
		.A1(out_sel[8]),
		.A2(I8[8]),
		.B1(out_sel[9]),
		.B2(I9[8]),
		.Z(O4[8])
	);
	AO_CELL inst_5_8(
		.A1(out_sel[10]),
		.A2(I10[8]),
		.B1(out_sel[11]),
		.B2(I11[8]),
		.Z(O5[8])
	);
	AO_CELL inst_6_8(
		.A1(out_sel[12]),
		.A2(I12[8]),
		.B1(out_sel[13]),
		.B2(I13[8]),
		.Z(O6[8])
	);
	AO_CELL inst_7_8(
		.A1(out_sel[14]),
		.A2(I14[8]),
		.B1(out_sel[15]),
		.B2(I15[8]),
		.Z(O7[8])
	);
	AO_CELL inst_8_8(
		.A1(out_sel[16]),
		.A2(I16[8]),
		.B1(out_sel[17]),
		.B2(I17[8]),
		.Z(O8[8])
	);
	AO_CELL inst_9_8(
		.A1(out_sel[18]),
		.A2(I18[8]),
		.B1(out_sel[19]),
		.B2(I19[8]),
		.Z(O9[8])
	);
	AO_CELL inst_10_8(
		.A1(out_sel[20]),
		.A2(I20[8]),
		.B1(out_sel[21]),
		.B2(1'b0),
		.Z(O10[8])
	);
	AO_CELL inst_0_9(
		.A1(out_sel[0]),
		.A2(I0[9]),
		.B1(out_sel[1]),
		.B2(I1[9]),
		.Z(O0[9])
	);
	AO_CELL inst_1_9(
		.A1(out_sel[2]),
		.A2(I2[9]),
		.B1(out_sel[3]),
		.B2(I3[9]),
		.Z(O1[9])
	);
	AO_CELL inst_2_9(
		.A1(out_sel[4]),
		.A2(I4[9]),
		.B1(out_sel[5]),
		.B2(I5[9]),
		.Z(O2[9])
	);
	AO_CELL inst_3_9(
		.A1(out_sel[6]),
		.A2(I6[9]),
		.B1(out_sel[7]),
		.B2(I7[9]),
		.Z(O3[9])
	);
	AO_CELL inst_4_9(
		.A1(out_sel[8]),
		.A2(I8[9]),
		.B1(out_sel[9]),
		.B2(I9[9]),
		.Z(O4[9])
	);
	AO_CELL inst_5_9(
		.A1(out_sel[10]),
		.A2(I10[9]),
		.B1(out_sel[11]),
		.B2(I11[9]),
		.Z(O5[9])
	);
	AO_CELL inst_6_9(
		.A1(out_sel[12]),
		.A2(I12[9]),
		.B1(out_sel[13]),
		.B2(I13[9]),
		.Z(O6[9])
	);
	AO_CELL inst_7_9(
		.A1(out_sel[14]),
		.A2(I14[9]),
		.B1(out_sel[15]),
		.B2(I15[9]),
		.Z(O7[9])
	);
	AO_CELL inst_8_9(
		.A1(out_sel[16]),
		.A2(I16[9]),
		.B1(out_sel[17]),
		.B2(I17[9]),
		.Z(O8[9])
	);
	AO_CELL inst_9_9(
		.A1(out_sel[18]),
		.A2(I18[9]),
		.B1(out_sel[19]),
		.B2(I19[9]),
		.Z(O9[9])
	);
	AO_CELL inst_10_9(
		.A1(out_sel[20]),
		.A2(I20[9]),
		.B1(out_sel[21]),
		.B2(1'b0),
		.Z(O10[9])
	);
	AO_CELL inst_0_10(
		.A1(out_sel[0]),
		.A2(I0[10]),
		.B1(out_sel[1]),
		.B2(I1[10]),
		.Z(O0[10])
	);
	AO_CELL inst_1_10(
		.A1(out_sel[2]),
		.A2(I2[10]),
		.B1(out_sel[3]),
		.B2(I3[10]),
		.Z(O1[10])
	);
	AO_CELL inst_2_10(
		.A1(out_sel[4]),
		.A2(I4[10]),
		.B1(out_sel[5]),
		.B2(I5[10]),
		.Z(O2[10])
	);
	AO_CELL inst_3_10(
		.A1(out_sel[6]),
		.A2(I6[10]),
		.B1(out_sel[7]),
		.B2(I7[10]),
		.Z(O3[10])
	);
	AO_CELL inst_4_10(
		.A1(out_sel[8]),
		.A2(I8[10]),
		.B1(out_sel[9]),
		.B2(I9[10]),
		.Z(O4[10])
	);
	AO_CELL inst_5_10(
		.A1(out_sel[10]),
		.A2(I10[10]),
		.B1(out_sel[11]),
		.B2(I11[10]),
		.Z(O5[10])
	);
	AO_CELL inst_6_10(
		.A1(out_sel[12]),
		.A2(I12[10]),
		.B1(out_sel[13]),
		.B2(I13[10]),
		.Z(O6[10])
	);
	AO_CELL inst_7_10(
		.A1(out_sel[14]),
		.A2(I14[10]),
		.B1(out_sel[15]),
		.B2(I15[10]),
		.Z(O7[10])
	);
	AO_CELL inst_8_10(
		.A1(out_sel[16]),
		.A2(I16[10]),
		.B1(out_sel[17]),
		.B2(I17[10]),
		.Z(O8[10])
	);
	AO_CELL inst_9_10(
		.A1(out_sel[18]),
		.A2(I18[10]),
		.B1(out_sel[19]),
		.B2(I19[10]),
		.Z(O9[10])
	);
	AO_CELL inst_10_10(
		.A1(out_sel[20]),
		.A2(I20[10]),
		.B1(out_sel[21]),
		.B2(1'b0),
		.Z(O10[10])
	);
	AO_CELL inst_0_11(
		.A1(out_sel[0]),
		.A2(I0[11]),
		.B1(out_sel[1]),
		.B2(I1[11]),
		.Z(O0[11])
	);
	AO_CELL inst_1_11(
		.A1(out_sel[2]),
		.A2(I2[11]),
		.B1(out_sel[3]),
		.B2(I3[11]),
		.Z(O1[11])
	);
	AO_CELL inst_2_11(
		.A1(out_sel[4]),
		.A2(I4[11]),
		.B1(out_sel[5]),
		.B2(I5[11]),
		.Z(O2[11])
	);
	AO_CELL inst_3_11(
		.A1(out_sel[6]),
		.A2(I6[11]),
		.B1(out_sel[7]),
		.B2(I7[11]),
		.Z(O3[11])
	);
	AO_CELL inst_4_11(
		.A1(out_sel[8]),
		.A2(I8[11]),
		.B1(out_sel[9]),
		.B2(I9[11]),
		.Z(O4[11])
	);
	AO_CELL inst_5_11(
		.A1(out_sel[10]),
		.A2(I10[11]),
		.B1(out_sel[11]),
		.B2(I11[11]),
		.Z(O5[11])
	);
	AO_CELL inst_6_11(
		.A1(out_sel[12]),
		.A2(I12[11]),
		.B1(out_sel[13]),
		.B2(I13[11]),
		.Z(O6[11])
	);
	AO_CELL inst_7_11(
		.A1(out_sel[14]),
		.A2(I14[11]),
		.B1(out_sel[15]),
		.B2(I15[11]),
		.Z(O7[11])
	);
	AO_CELL inst_8_11(
		.A1(out_sel[16]),
		.A2(I16[11]),
		.B1(out_sel[17]),
		.B2(I17[11]),
		.Z(O8[11])
	);
	AO_CELL inst_9_11(
		.A1(out_sel[18]),
		.A2(I18[11]),
		.B1(out_sel[19]),
		.B2(I19[11]),
		.Z(O9[11])
	);
	AO_CELL inst_10_11(
		.A1(out_sel[20]),
		.A2(I20[11]),
		.B1(out_sel[21]),
		.B2(1'b0),
		.Z(O10[11])
	);
	AO_CELL inst_0_12(
		.A1(out_sel[0]),
		.A2(I0[12]),
		.B1(out_sel[1]),
		.B2(I1[12]),
		.Z(O0[12])
	);
	AO_CELL inst_1_12(
		.A1(out_sel[2]),
		.A2(I2[12]),
		.B1(out_sel[3]),
		.B2(I3[12]),
		.Z(O1[12])
	);
	AO_CELL inst_2_12(
		.A1(out_sel[4]),
		.A2(I4[12]),
		.B1(out_sel[5]),
		.B2(I5[12]),
		.Z(O2[12])
	);
	AO_CELL inst_3_12(
		.A1(out_sel[6]),
		.A2(I6[12]),
		.B1(out_sel[7]),
		.B2(I7[12]),
		.Z(O3[12])
	);
	AO_CELL inst_4_12(
		.A1(out_sel[8]),
		.A2(I8[12]),
		.B1(out_sel[9]),
		.B2(I9[12]),
		.Z(O4[12])
	);
	AO_CELL inst_5_12(
		.A1(out_sel[10]),
		.A2(I10[12]),
		.B1(out_sel[11]),
		.B2(I11[12]),
		.Z(O5[12])
	);
	AO_CELL inst_6_12(
		.A1(out_sel[12]),
		.A2(I12[12]),
		.B1(out_sel[13]),
		.B2(I13[12]),
		.Z(O6[12])
	);
	AO_CELL inst_7_12(
		.A1(out_sel[14]),
		.A2(I14[12]),
		.B1(out_sel[15]),
		.B2(I15[12]),
		.Z(O7[12])
	);
	AO_CELL inst_8_12(
		.A1(out_sel[16]),
		.A2(I16[12]),
		.B1(out_sel[17]),
		.B2(I17[12]),
		.Z(O8[12])
	);
	AO_CELL inst_9_12(
		.A1(out_sel[18]),
		.A2(I18[12]),
		.B1(out_sel[19]),
		.B2(I19[12]),
		.Z(O9[12])
	);
	AO_CELL inst_10_12(
		.A1(out_sel[20]),
		.A2(I20[12]),
		.B1(out_sel[21]),
		.B2(1'b0),
		.Z(O10[12])
	);
	AO_CELL inst_0_13(
		.A1(out_sel[0]),
		.A2(I0[13]),
		.B1(out_sel[1]),
		.B2(I1[13]),
		.Z(O0[13])
	);
	AO_CELL inst_1_13(
		.A1(out_sel[2]),
		.A2(I2[13]),
		.B1(out_sel[3]),
		.B2(I3[13]),
		.Z(O1[13])
	);
	AO_CELL inst_2_13(
		.A1(out_sel[4]),
		.A2(I4[13]),
		.B1(out_sel[5]),
		.B2(I5[13]),
		.Z(O2[13])
	);
	AO_CELL inst_3_13(
		.A1(out_sel[6]),
		.A2(I6[13]),
		.B1(out_sel[7]),
		.B2(I7[13]),
		.Z(O3[13])
	);
	AO_CELL inst_4_13(
		.A1(out_sel[8]),
		.A2(I8[13]),
		.B1(out_sel[9]),
		.B2(I9[13]),
		.Z(O4[13])
	);
	AO_CELL inst_5_13(
		.A1(out_sel[10]),
		.A2(I10[13]),
		.B1(out_sel[11]),
		.B2(I11[13]),
		.Z(O5[13])
	);
	AO_CELL inst_6_13(
		.A1(out_sel[12]),
		.A2(I12[13]),
		.B1(out_sel[13]),
		.B2(I13[13]),
		.Z(O6[13])
	);
	AO_CELL inst_7_13(
		.A1(out_sel[14]),
		.A2(I14[13]),
		.B1(out_sel[15]),
		.B2(I15[13]),
		.Z(O7[13])
	);
	AO_CELL inst_8_13(
		.A1(out_sel[16]),
		.A2(I16[13]),
		.B1(out_sel[17]),
		.B2(I17[13]),
		.Z(O8[13])
	);
	AO_CELL inst_9_13(
		.A1(out_sel[18]),
		.A2(I18[13]),
		.B1(out_sel[19]),
		.B2(I19[13]),
		.Z(O9[13])
	);
	AO_CELL inst_10_13(
		.A1(out_sel[20]),
		.A2(I20[13]),
		.B1(out_sel[21]),
		.B2(1'b0),
		.Z(O10[13])
	);
	AO_CELL inst_0_14(
		.A1(out_sel[0]),
		.A2(I0[14]),
		.B1(out_sel[1]),
		.B2(I1[14]),
		.Z(O0[14])
	);
	AO_CELL inst_1_14(
		.A1(out_sel[2]),
		.A2(I2[14]),
		.B1(out_sel[3]),
		.B2(I3[14]),
		.Z(O1[14])
	);
	AO_CELL inst_2_14(
		.A1(out_sel[4]),
		.A2(I4[14]),
		.B1(out_sel[5]),
		.B2(I5[14]),
		.Z(O2[14])
	);
	AO_CELL inst_3_14(
		.A1(out_sel[6]),
		.A2(I6[14]),
		.B1(out_sel[7]),
		.B2(I7[14]),
		.Z(O3[14])
	);
	AO_CELL inst_4_14(
		.A1(out_sel[8]),
		.A2(I8[14]),
		.B1(out_sel[9]),
		.B2(I9[14]),
		.Z(O4[14])
	);
	AO_CELL inst_5_14(
		.A1(out_sel[10]),
		.A2(I10[14]),
		.B1(out_sel[11]),
		.B2(I11[14]),
		.Z(O5[14])
	);
	AO_CELL inst_6_14(
		.A1(out_sel[12]),
		.A2(I12[14]),
		.B1(out_sel[13]),
		.B2(I13[14]),
		.Z(O6[14])
	);
	AO_CELL inst_7_14(
		.A1(out_sel[14]),
		.A2(I14[14]),
		.B1(out_sel[15]),
		.B2(I15[14]),
		.Z(O7[14])
	);
	AO_CELL inst_8_14(
		.A1(out_sel[16]),
		.A2(I16[14]),
		.B1(out_sel[17]),
		.B2(I17[14]),
		.Z(O8[14])
	);
	AO_CELL inst_9_14(
		.A1(out_sel[18]),
		.A2(I18[14]),
		.B1(out_sel[19]),
		.B2(I19[14]),
		.Z(O9[14])
	);
	AO_CELL inst_10_14(
		.A1(out_sel[20]),
		.A2(I20[14]),
		.B1(out_sel[21]),
		.B2(1'b0),
		.Z(O10[14])
	);
	AO_CELL inst_0_15(
		.A1(out_sel[0]),
		.A2(I0[15]),
		.B1(out_sel[1]),
		.B2(I1[15]),
		.Z(O0[15])
	);
	AO_CELL inst_1_15(
		.A1(out_sel[2]),
		.A2(I2[15]),
		.B1(out_sel[3]),
		.B2(I3[15]),
		.Z(O1[15])
	);
	AO_CELL inst_2_15(
		.A1(out_sel[4]),
		.A2(I4[15]),
		.B1(out_sel[5]),
		.B2(I5[15]),
		.Z(O2[15])
	);
	AO_CELL inst_3_15(
		.A1(out_sel[6]),
		.A2(I6[15]),
		.B1(out_sel[7]),
		.B2(I7[15]),
		.Z(O3[15])
	);
	AO_CELL inst_4_15(
		.A1(out_sel[8]),
		.A2(I8[15]),
		.B1(out_sel[9]),
		.B2(I9[15]),
		.Z(O4[15])
	);
	AO_CELL inst_5_15(
		.A1(out_sel[10]),
		.A2(I10[15]),
		.B1(out_sel[11]),
		.B2(I11[15]),
		.Z(O5[15])
	);
	AO_CELL inst_6_15(
		.A1(out_sel[12]),
		.A2(I12[15]),
		.B1(out_sel[13]),
		.B2(I13[15]),
		.Z(O6[15])
	);
	AO_CELL inst_7_15(
		.A1(out_sel[14]),
		.A2(I14[15]),
		.B1(out_sel[15]),
		.B2(I15[15]),
		.Z(O7[15])
	);
	AO_CELL inst_8_15(
		.A1(out_sel[16]),
		.A2(I16[15]),
		.B1(out_sel[17]),
		.B2(I17[15]),
		.Z(O8[15])
	);
	AO_CELL inst_9_15(
		.A1(out_sel[18]),
		.A2(I18[15]),
		.B1(out_sel[19]),
		.B2(I19[15]),
		.Z(O9[15])
	);
	AO_CELL inst_10_15(
		.A1(out_sel[20]),
		.A2(I20[15]),
		.B1(out_sel[21]),
		.B2(1'b0),
		.Z(O10[15])
	);
	AO_CELL inst_0_16(
		.A1(out_sel[0]),
		.A2(I0[16]),
		.B1(out_sel[1]),
		.B2(I1[16]),
		.Z(O0[16])
	);
	AO_CELL inst_1_16(
		.A1(out_sel[2]),
		.A2(I2[16]),
		.B1(out_sel[3]),
		.B2(I3[16]),
		.Z(O1[16])
	);
	AO_CELL inst_2_16(
		.A1(out_sel[4]),
		.A2(I4[16]),
		.B1(out_sel[5]),
		.B2(I5[16]),
		.Z(O2[16])
	);
	AO_CELL inst_3_16(
		.A1(out_sel[6]),
		.A2(I6[16]),
		.B1(out_sel[7]),
		.B2(I7[16]),
		.Z(O3[16])
	);
	AO_CELL inst_4_16(
		.A1(out_sel[8]),
		.A2(I8[16]),
		.B1(out_sel[9]),
		.B2(I9[16]),
		.Z(O4[16])
	);
	AO_CELL inst_5_16(
		.A1(out_sel[10]),
		.A2(I10[16]),
		.B1(out_sel[11]),
		.B2(I11[16]),
		.Z(O5[16])
	);
	AO_CELL inst_6_16(
		.A1(out_sel[12]),
		.A2(I12[16]),
		.B1(out_sel[13]),
		.B2(I13[16]),
		.Z(O6[16])
	);
	AO_CELL inst_7_16(
		.A1(out_sel[14]),
		.A2(I14[16]),
		.B1(out_sel[15]),
		.B2(I15[16]),
		.Z(O7[16])
	);
	AO_CELL inst_8_16(
		.A1(out_sel[16]),
		.A2(I16[16]),
		.B1(out_sel[17]),
		.B2(I17[16]),
		.Z(O8[16])
	);
	AO_CELL inst_9_16(
		.A1(out_sel[18]),
		.A2(I18[16]),
		.B1(out_sel[19]),
		.B2(I19[16]),
		.Z(O9[16])
	);
	AO_CELL inst_10_16(
		.A1(out_sel[20]),
		.A2(I20[16]),
		.B1(out_sel[21]),
		.B2(1'b0),
		.Z(O10[16])
	);
	AO_CELL inst_0_valid(
		.A1(out_sel[0]),
		.A2(valid_in[0]),
		.B1(out_sel[1]),
		.B2(valid_in[1]),
		.Z(valid_out[0])
	);
	AO_CELL inst_1_valid(
		.A1(out_sel[2]),
		.A2(valid_in[2]),
		.B1(out_sel[3]),
		.B2(valid_in[3]),
		.Z(valid_out[1])
	);
	AO_CELL inst_2_valid(
		.A1(out_sel[4]),
		.A2(valid_in[4]),
		.B1(out_sel[5]),
		.B2(valid_in[5]),
		.Z(valid_out[2])
	);
	AO_CELL inst_3_valid(
		.A1(out_sel[6]),
		.A2(valid_in[6]),
		.B1(out_sel[7]),
		.B2(valid_in[7]),
		.Z(valid_out[3])
	);
	AO_CELL inst_4_valid(
		.A1(out_sel[8]),
		.A2(valid_in[8]),
		.B1(out_sel[9]),
		.B2(valid_in[9]),
		.Z(valid_out[4])
	);
	AO_CELL inst_5_valid(
		.A1(out_sel[10]),
		.A2(valid_in[10]),
		.B1(out_sel[11]),
		.B2(valid_in[11]),
		.Z(valid_out[5])
	);
	AO_CELL inst_6_valid(
		.A1(out_sel[12]),
		.A2(valid_in[12]),
		.B1(out_sel[13]),
		.B2(valid_in[13]),
		.Z(valid_out[6])
	);
	AO_CELL inst_7_valid(
		.A1(out_sel[14]),
		.A2(valid_in[14]),
		.B1(out_sel[15]),
		.B2(valid_in[15]),
		.Z(valid_out[7])
	);
	AO_CELL inst_8_valid(
		.A1(out_sel[16]),
		.A2(valid_in[16]),
		.B1(out_sel[17]),
		.B2(valid_in[17]),
		.Z(valid_out[8])
	);
	AO_CELL inst_9_valid(
		.A1(out_sel[18]),
		.A2(valid_in[18]),
		.B1(out_sel[19]),
		.B2(valid_in[19]),
		.Z(valid_out[9])
	);
	AO_CELL inst_10_valid(
		.A1(out_sel[20]),
		.A2(valid_in[20]),
		.B1(out_sel[21]),
		.B2(1'b0),
		.Z(valid_out[10])
	);
endmodule
module mux_aoi_ready_valid_const_21_1 (
	I,
	S,
	ready_in,
	ready_out,
	valid_in,
	valid_out,
	out_sel,
	O
);
	input wire [20:0] I;
	input wire [4:0] S;
	input wire ready_in;
	output wire ready_out;
	input wire [20:0] valid_in;
	output wire valid_out;
	output wire [31:0] out_sel;
	output wire [0:0] O;
	wire [0:0] O_int0;
	wire [0:0] O_int1;
	wire [0:0] O_int2;
	wire [0:0] O_int3;
	wire [0:0] O_int4;
	wire [0:0] O_int5;
	wire [0:0] O_int6;
	wire [0:0] O_int7;
	wire [0:0] O_int8;
	wire [0:0] O_int9;
	wire [0:0] O_int10;
	wire [10:0] valid_out_temp;
	precoder_1_21 u_precoder(
		.S(S),
		.out_sel(out_sel)
	);
	mux_logic_1_21 u_mux_logic(
		.I0(I[0+:1]),
		.I1(I[1+:1]),
		.I2(I[2+:1]),
		.I3(I[3+:1]),
		.I4(I[4+:1]),
		.I5(I[5+:1]),
		.I6(I[6+:1]),
		.I7(I[7+:1]),
		.I8(I[8+:1]),
		.I9(I[9+:1]),
		.I10(I[10+:1]),
		.I11(I[11+:1]),
		.I12(I[12+:1]),
		.I13(I[13+:1]),
		.I14(I[14+:1]),
		.I15(I[15+:1]),
		.I16(I[16+:1]),
		.I17(I[17+:1]),
		.I18(I[18+:1]),
		.I19(I[19+:1]),
		.I20(I[20+:1]),
		.out_sel(out_sel),
		.valid_in(valid_in),
		.valid_out(valid_out_temp),
		.O0(O_int0),
		.O1(O_int1),
		.O2(O_int2),
		.O3(O_int3),
		.O4(O_int4),
		.O5(O_int5),
		.O6(O_int6),
		.O7(O_int7),
		.O8(O_int8),
		.O9(O_int9),
		.O10(O_int10)
	);
	assign O = (((((((((O_int0 | O_int1) | O_int2) | O_int3) | O_int4) | O_int5) | O_int6) | O_int7) | O_int8) | O_int9) | O_int10;
	assign ready_out = ready_in;
	assign valid_out = |valid_out_temp;
endmodule
module precoder_1_21 (
	S,
	out_sel
);
	input wire [4:0] S;
	output reg [31:0] out_sel;
	always @(*) begin : mux_sel
		case (S)
			5'd0: out_sel = 32'b00000000000000000000000000000001;
			5'd1: out_sel = 32'b00000000000000000000000000000010;
			5'd2: out_sel = 32'b00000000000000000000000000000100;
			5'd3: out_sel = 32'b00000000000000000000000000001000;
			5'd4: out_sel = 32'b00000000000000000000000000010000;
			5'd5: out_sel = 32'b00000000000000000000000000100000;
			5'd6: out_sel = 32'b00000000000000000000000001000000;
			5'd7: out_sel = 32'b00000000000000000000000010000000;
			5'd8: out_sel = 32'b00000000000000000000000100000000;
			5'd9: out_sel = 32'b00000000000000000000001000000000;
			5'd10: out_sel = 32'b00000000000000000000010000000000;
			5'd11: out_sel = 32'b00000000000000000000100000000000;
			5'd12: out_sel = 32'b00000000000000000001000000000000;
			5'd13: out_sel = 32'b00000000000000000010000000000000;
			5'd14: out_sel = 32'b00000000000000000100000000000000;
			5'd15: out_sel = 32'b00000000000000001000000000000000;
			5'd16: out_sel = 32'b00000000000000010000000000000000;
			5'd17: out_sel = 32'b00000000000000100000000000000000;
			5'd18: out_sel = 32'b00000000000001000000000000000000;
			5'd19: out_sel = 32'b00000000000010000000000000000000;
			5'd20: out_sel = 32'b00000000000100000000000000000000;
			5'd21: out_sel = 32'b00000000001000000000000000000000;
			default: out_sel = 32'b00000000000000000000000000000000;
		endcase
	end
endmodule
module mux_logic_1_21 (
	out_sel,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	I9,
	I10,
	I11,
	I12,
	I13,
	I14,
	I15,
	I16,
	I17,
	I18,
	I19,
	I20,
	valid_in,
	valid_out,
	O0,
	O1,
	O2,
	O3,
	O4,
	O5,
	O6,
	O7,
	O8,
	O9,
	O10
);
	input wire [31:0] out_sel;
	input wire [0:0] I0;
	input wire [0:0] I1;
	input wire [0:0] I2;
	input wire [0:0] I3;
	input wire [0:0] I4;
	input wire [0:0] I5;
	input wire [0:0] I6;
	input wire [0:0] I7;
	input wire [0:0] I8;
	input wire [0:0] I9;
	input wire [0:0] I10;
	input wire [0:0] I11;
	input wire [0:0] I12;
	input wire [0:0] I13;
	input wire [0:0] I14;
	input wire [0:0] I15;
	input wire [0:0] I16;
	input wire [0:0] I17;
	input wire [0:0] I18;
	input wire [0:0] I19;
	input wire [0:0] I20;
	input wire [20:0] valid_in;
	output wire [10:0] valid_out;
	output wire [0:0] O0;
	output wire [0:0] O1;
	output wire [0:0] O2;
	output wire [0:0] O3;
	output wire [0:0] O4;
	output wire [0:0] O5;
	output wire [0:0] O6;
	output wire [0:0] O7;
	output wire [0:0] O8;
	output wire [0:0] O9;
	output wire [0:0] O10;
	AO_CELL inst_0_0(
		.A1(out_sel[0]),
		.A2(I0[0]),
		.B1(out_sel[1]),
		.B2(I1[0]),
		.Z(O0[0])
	);
	AO_CELL inst_1_0(
		.A1(out_sel[2]),
		.A2(I2[0]),
		.B1(out_sel[3]),
		.B2(I3[0]),
		.Z(O1[0])
	);
	AO_CELL inst_2_0(
		.A1(out_sel[4]),
		.A2(I4[0]),
		.B1(out_sel[5]),
		.B2(I5[0]),
		.Z(O2[0])
	);
	AO_CELL inst_3_0(
		.A1(out_sel[6]),
		.A2(I6[0]),
		.B1(out_sel[7]),
		.B2(I7[0]),
		.Z(O3[0])
	);
	AO_CELL inst_4_0(
		.A1(out_sel[8]),
		.A2(I8[0]),
		.B1(out_sel[9]),
		.B2(I9[0]),
		.Z(O4[0])
	);
	AO_CELL inst_5_0(
		.A1(out_sel[10]),
		.A2(I10[0]),
		.B1(out_sel[11]),
		.B2(I11[0]),
		.Z(O5[0])
	);
	AO_CELL inst_6_0(
		.A1(out_sel[12]),
		.A2(I12[0]),
		.B1(out_sel[13]),
		.B2(I13[0]),
		.Z(O6[0])
	);
	AO_CELL inst_7_0(
		.A1(out_sel[14]),
		.A2(I14[0]),
		.B1(out_sel[15]),
		.B2(I15[0]),
		.Z(O7[0])
	);
	AO_CELL inst_8_0(
		.A1(out_sel[16]),
		.A2(I16[0]),
		.B1(out_sel[17]),
		.B2(I17[0]),
		.Z(O8[0])
	);
	AO_CELL inst_9_0(
		.A1(out_sel[18]),
		.A2(I18[0]),
		.B1(out_sel[19]),
		.B2(I19[0]),
		.Z(O9[0])
	);
	AO_CELL inst_10_0(
		.A1(out_sel[20]),
		.A2(I20[0]),
		.B1(out_sel[21]),
		.B2(1'b0),
		.Z(O10[0])
	);
	AO_CELL inst_0_valid(
		.A1(out_sel[0]),
		.A2(valid_in[0]),
		.B1(out_sel[1]),
		.B2(valid_in[1]),
		.Z(valid_out[0])
	);
	AO_CELL inst_1_valid(
		.A1(out_sel[2]),
		.A2(valid_in[2]),
		.B1(out_sel[3]),
		.B2(valid_in[3]),
		.Z(valid_out[1])
	);
	AO_CELL inst_2_valid(
		.A1(out_sel[4]),
		.A2(valid_in[4]),
		.B1(out_sel[5]),
		.B2(valid_in[5]),
		.Z(valid_out[2])
	);
	AO_CELL inst_3_valid(
		.A1(out_sel[6]),
		.A2(valid_in[6]),
		.B1(out_sel[7]),
		.B2(valid_in[7]),
		.Z(valid_out[3])
	);
	AO_CELL inst_4_valid(
		.A1(out_sel[8]),
		.A2(valid_in[8]),
		.B1(out_sel[9]),
		.B2(valid_in[9]),
		.Z(valid_out[4])
	);
	AO_CELL inst_5_valid(
		.A1(out_sel[10]),
		.A2(valid_in[10]),
		.B1(out_sel[11]),
		.B2(valid_in[11]),
		.Z(valid_out[5])
	);
	AO_CELL inst_6_valid(
		.A1(out_sel[12]),
		.A2(valid_in[12]),
		.B1(out_sel[13]),
		.B2(valid_in[13]),
		.Z(valid_out[6])
	);
	AO_CELL inst_7_valid(
		.A1(out_sel[14]),
		.A2(valid_in[14]),
		.B1(out_sel[15]),
		.B2(valid_in[15]),
		.Z(valid_out[7])
	);
	AO_CELL inst_8_valid(
		.A1(out_sel[16]),
		.A2(valid_in[16]),
		.B1(out_sel[17]),
		.B2(valid_in[17]),
		.Z(valid_out[8])
	);
	AO_CELL inst_9_valid(
		.A1(out_sel[18]),
		.A2(valid_in[18]),
		.B1(out_sel[19]),
		.B2(valid_in[19]),
		.Z(valid_out[9])
	);
	AO_CELL inst_10_valid(
		.A1(out_sel[20]),
		.A2(valid_in[20]),
		.B1(out_sel[21]),
		.B2(1'b0),
		.Z(valid_out[10])
	);
endmodule
module mux_aoi_ready_valid_const_20_17 (
	I,
	S,
	ready_in,
	ready_out,
	valid_in,
	valid_out,
	out_sel,
	O
);
	input wire [339:0] I;
	input wire [4:0] S;
	input wire ready_in;
	output wire ready_out;
	input wire [19:0] valid_in;
	output wire valid_out;
	output wire [31:0] out_sel;
	output wire [16:0] O;
	wire [16:0] O_int0;
	wire [16:0] O_int1;
	wire [16:0] O_int2;
	wire [16:0] O_int3;
	wire [16:0] O_int4;
	wire [16:0] O_int5;
	wire [16:0] O_int6;
	wire [16:0] O_int7;
	wire [16:0] O_int8;
	wire [16:0] O_int9;
	wire [16:0] O_int10;
	wire [10:0] valid_out_temp;
	precoder_17_20 u_precoder(
		.S(S),
		.out_sel(out_sel)
	);
	mux_logic_17_20 u_mux_logic(
		.I0(I[0+:17]),
		.I1(I[17+:17]),
		.I2(I[34+:17]),
		.I3(I[51+:17]),
		.I4(I[68+:17]),
		.I5(I[85+:17]),
		.I6(I[102+:17]),
		.I7(I[119+:17]),
		.I8(I[136+:17]),
		.I9(I[153+:17]),
		.I10(I[170+:17]),
		.I11(I[187+:17]),
		.I12(I[204+:17]),
		.I13(I[221+:17]),
		.I14(I[238+:17]),
		.I15(I[255+:17]),
		.I16(I[272+:17]),
		.I17(I[289+:17]),
		.I18(I[306+:17]),
		.I19(I[323+:17]),
		.out_sel(out_sel),
		.valid_in(valid_in),
		.valid_out(valid_out_temp),
		.O0(O_int0),
		.O1(O_int1),
		.O2(O_int2),
		.O3(O_int3),
		.O4(O_int4),
		.O5(O_int5),
		.O6(O_int6),
		.O7(O_int7),
		.O8(O_int8),
		.O9(O_int9),
		.O10(O_int10)
	);
	assign O = (((((((((O_int0 | O_int1) | O_int2) | O_int3) | O_int4) | O_int5) | O_int6) | O_int7) | O_int8) | O_int9) | O_int10;
	assign ready_out = ready_in;
	assign valid_out = |valid_out_temp;
endmodule
module precoder_17_20 (
	S,
	out_sel
);
	input wire [4:0] S;
	output reg [31:0] out_sel;
	always @(*) begin : mux_sel
		case (S)
			5'd0: out_sel = 32'b00000000000000000000000000000001;
			5'd1: out_sel = 32'b00000000000000000000000000000010;
			5'd2: out_sel = 32'b00000000000000000000000000000100;
			5'd3: out_sel = 32'b00000000000000000000000000001000;
			5'd4: out_sel = 32'b00000000000000000000000000010000;
			5'd5: out_sel = 32'b00000000000000000000000000100000;
			5'd6: out_sel = 32'b00000000000000000000000001000000;
			5'd7: out_sel = 32'b00000000000000000000000010000000;
			5'd8: out_sel = 32'b00000000000000000000000100000000;
			5'd9: out_sel = 32'b00000000000000000000001000000000;
			5'd10: out_sel = 32'b00000000000000000000010000000000;
			5'd11: out_sel = 32'b00000000000000000000100000000000;
			5'd12: out_sel = 32'b00000000000000000001000000000000;
			5'd13: out_sel = 32'b00000000000000000010000000000000;
			5'd14: out_sel = 32'b00000000000000000100000000000000;
			5'd15: out_sel = 32'b00000000000000001000000000000000;
			5'd16: out_sel = 32'b00000000000000010000000000000000;
			5'd17: out_sel = 32'b00000000000000100000000000000000;
			5'd18: out_sel = 32'b00000000000001000000000000000000;
			5'd19: out_sel = 32'b00000000000010000000000000000000;
			5'd20: out_sel = 32'b00000000000100000000000000000000;
			default: out_sel = 32'b00000000000000000000000000000000;
		endcase
	end
endmodule
module mux_logic_17_20 (
	out_sel,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	I9,
	I10,
	I11,
	I12,
	I13,
	I14,
	I15,
	I16,
	I17,
	I18,
	I19,
	valid_in,
	valid_out,
	O0,
	O1,
	O2,
	O3,
	O4,
	O5,
	O6,
	O7,
	O8,
	O9,
	O10
);
	input wire [31:0] out_sel;
	input wire [16:0] I0;
	input wire [16:0] I1;
	input wire [16:0] I2;
	input wire [16:0] I3;
	input wire [16:0] I4;
	input wire [16:0] I5;
	input wire [16:0] I6;
	input wire [16:0] I7;
	input wire [16:0] I8;
	input wire [16:0] I9;
	input wire [16:0] I10;
	input wire [16:0] I11;
	input wire [16:0] I12;
	input wire [16:0] I13;
	input wire [16:0] I14;
	input wire [16:0] I15;
	input wire [16:0] I16;
	input wire [16:0] I17;
	input wire [16:0] I18;
	input wire [16:0] I19;
	input wire [19:0] valid_in;
	output wire [10:0] valid_out;
	output wire [16:0] O0;
	output wire [16:0] O1;
	output wire [16:0] O2;
	output wire [16:0] O3;
	output wire [16:0] O4;
	output wire [16:0] O5;
	output wire [16:0] O6;
	output wire [16:0] O7;
	output wire [16:0] O8;
	output wire [16:0] O9;
	output wire [16:0] O10;
	AO_CELL inst_0_0(
		.A1(out_sel[0]),
		.A2(I0[0]),
		.B1(out_sel[1]),
		.B2(I1[0]),
		.Z(O0[0])
	);
	AO_CELL inst_1_0(
		.A1(out_sel[2]),
		.A2(I2[0]),
		.B1(out_sel[3]),
		.B2(I3[0]),
		.Z(O1[0])
	);
	AO_CELL inst_2_0(
		.A1(out_sel[4]),
		.A2(I4[0]),
		.B1(out_sel[5]),
		.B2(I5[0]),
		.Z(O2[0])
	);
	AO_CELL inst_3_0(
		.A1(out_sel[6]),
		.A2(I6[0]),
		.B1(out_sel[7]),
		.B2(I7[0]),
		.Z(O3[0])
	);
	AO_CELL inst_4_0(
		.A1(out_sel[8]),
		.A2(I8[0]),
		.B1(out_sel[9]),
		.B2(I9[0]),
		.Z(O4[0])
	);
	AO_CELL inst_5_0(
		.A1(out_sel[10]),
		.A2(I10[0]),
		.B1(out_sel[11]),
		.B2(I11[0]),
		.Z(O5[0])
	);
	AO_CELL inst_6_0(
		.A1(out_sel[12]),
		.A2(I12[0]),
		.B1(out_sel[13]),
		.B2(I13[0]),
		.Z(O6[0])
	);
	AO_CELL inst_7_0(
		.A1(out_sel[14]),
		.A2(I14[0]),
		.B1(out_sel[15]),
		.B2(I15[0]),
		.Z(O7[0])
	);
	AO_CELL inst_8_0(
		.A1(out_sel[16]),
		.A2(I16[0]),
		.B1(out_sel[17]),
		.B2(I17[0]),
		.Z(O8[0])
	);
	AO_CELL inst_9_0(
		.A1(out_sel[18]),
		.A2(I18[0]),
		.B1(out_sel[19]),
		.B2(I19[0]),
		.Z(O9[0])
	);
	AN_CELL inst_and_0(
		.A1(out_sel[20]),
		.A2(1'b0),
		.Z(O10[0])
	);
	AO_CELL inst_0_1(
		.A1(out_sel[0]),
		.A2(I0[1]),
		.B1(out_sel[1]),
		.B2(I1[1]),
		.Z(O0[1])
	);
	AO_CELL inst_1_1(
		.A1(out_sel[2]),
		.A2(I2[1]),
		.B1(out_sel[3]),
		.B2(I3[1]),
		.Z(O1[1])
	);
	AO_CELL inst_2_1(
		.A1(out_sel[4]),
		.A2(I4[1]),
		.B1(out_sel[5]),
		.B2(I5[1]),
		.Z(O2[1])
	);
	AO_CELL inst_3_1(
		.A1(out_sel[6]),
		.A2(I6[1]),
		.B1(out_sel[7]),
		.B2(I7[1]),
		.Z(O3[1])
	);
	AO_CELL inst_4_1(
		.A1(out_sel[8]),
		.A2(I8[1]),
		.B1(out_sel[9]),
		.B2(I9[1]),
		.Z(O4[1])
	);
	AO_CELL inst_5_1(
		.A1(out_sel[10]),
		.A2(I10[1]),
		.B1(out_sel[11]),
		.B2(I11[1]),
		.Z(O5[1])
	);
	AO_CELL inst_6_1(
		.A1(out_sel[12]),
		.A2(I12[1]),
		.B1(out_sel[13]),
		.B2(I13[1]),
		.Z(O6[1])
	);
	AO_CELL inst_7_1(
		.A1(out_sel[14]),
		.A2(I14[1]),
		.B1(out_sel[15]),
		.B2(I15[1]),
		.Z(O7[1])
	);
	AO_CELL inst_8_1(
		.A1(out_sel[16]),
		.A2(I16[1]),
		.B1(out_sel[17]),
		.B2(I17[1]),
		.Z(O8[1])
	);
	AO_CELL inst_9_1(
		.A1(out_sel[18]),
		.A2(I18[1]),
		.B1(out_sel[19]),
		.B2(I19[1]),
		.Z(O9[1])
	);
	AN_CELL inst_and_1(
		.A1(out_sel[20]),
		.A2(1'b0),
		.Z(O10[1])
	);
	AO_CELL inst_0_2(
		.A1(out_sel[0]),
		.A2(I0[2]),
		.B1(out_sel[1]),
		.B2(I1[2]),
		.Z(O0[2])
	);
	AO_CELL inst_1_2(
		.A1(out_sel[2]),
		.A2(I2[2]),
		.B1(out_sel[3]),
		.B2(I3[2]),
		.Z(O1[2])
	);
	AO_CELL inst_2_2(
		.A1(out_sel[4]),
		.A2(I4[2]),
		.B1(out_sel[5]),
		.B2(I5[2]),
		.Z(O2[2])
	);
	AO_CELL inst_3_2(
		.A1(out_sel[6]),
		.A2(I6[2]),
		.B1(out_sel[7]),
		.B2(I7[2]),
		.Z(O3[2])
	);
	AO_CELL inst_4_2(
		.A1(out_sel[8]),
		.A2(I8[2]),
		.B1(out_sel[9]),
		.B2(I9[2]),
		.Z(O4[2])
	);
	AO_CELL inst_5_2(
		.A1(out_sel[10]),
		.A2(I10[2]),
		.B1(out_sel[11]),
		.B2(I11[2]),
		.Z(O5[2])
	);
	AO_CELL inst_6_2(
		.A1(out_sel[12]),
		.A2(I12[2]),
		.B1(out_sel[13]),
		.B2(I13[2]),
		.Z(O6[2])
	);
	AO_CELL inst_7_2(
		.A1(out_sel[14]),
		.A2(I14[2]),
		.B1(out_sel[15]),
		.B2(I15[2]),
		.Z(O7[2])
	);
	AO_CELL inst_8_2(
		.A1(out_sel[16]),
		.A2(I16[2]),
		.B1(out_sel[17]),
		.B2(I17[2]),
		.Z(O8[2])
	);
	AO_CELL inst_9_2(
		.A1(out_sel[18]),
		.A2(I18[2]),
		.B1(out_sel[19]),
		.B2(I19[2]),
		.Z(O9[2])
	);
	AN_CELL inst_and_2(
		.A1(out_sel[20]),
		.A2(1'b0),
		.Z(O10[2])
	);
	AO_CELL inst_0_3(
		.A1(out_sel[0]),
		.A2(I0[3]),
		.B1(out_sel[1]),
		.B2(I1[3]),
		.Z(O0[3])
	);
	AO_CELL inst_1_3(
		.A1(out_sel[2]),
		.A2(I2[3]),
		.B1(out_sel[3]),
		.B2(I3[3]),
		.Z(O1[3])
	);
	AO_CELL inst_2_3(
		.A1(out_sel[4]),
		.A2(I4[3]),
		.B1(out_sel[5]),
		.B2(I5[3]),
		.Z(O2[3])
	);
	AO_CELL inst_3_3(
		.A1(out_sel[6]),
		.A2(I6[3]),
		.B1(out_sel[7]),
		.B2(I7[3]),
		.Z(O3[3])
	);
	AO_CELL inst_4_3(
		.A1(out_sel[8]),
		.A2(I8[3]),
		.B1(out_sel[9]),
		.B2(I9[3]),
		.Z(O4[3])
	);
	AO_CELL inst_5_3(
		.A1(out_sel[10]),
		.A2(I10[3]),
		.B1(out_sel[11]),
		.B2(I11[3]),
		.Z(O5[3])
	);
	AO_CELL inst_6_3(
		.A1(out_sel[12]),
		.A2(I12[3]),
		.B1(out_sel[13]),
		.B2(I13[3]),
		.Z(O6[3])
	);
	AO_CELL inst_7_3(
		.A1(out_sel[14]),
		.A2(I14[3]),
		.B1(out_sel[15]),
		.B2(I15[3]),
		.Z(O7[3])
	);
	AO_CELL inst_8_3(
		.A1(out_sel[16]),
		.A2(I16[3]),
		.B1(out_sel[17]),
		.B2(I17[3]),
		.Z(O8[3])
	);
	AO_CELL inst_9_3(
		.A1(out_sel[18]),
		.A2(I18[3]),
		.B1(out_sel[19]),
		.B2(I19[3]),
		.Z(O9[3])
	);
	AN_CELL inst_and_3(
		.A1(out_sel[20]),
		.A2(1'b0),
		.Z(O10[3])
	);
	AO_CELL inst_0_4(
		.A1(out_sel[0]),
		.A2(I0[4]),
		.B1(out_sel[1]),
		.B2(I1[4]),
		.Z(O0[4])
	);
	AO_CELL inst_1_4(
		.A1(out_sel[2]),
		.A2(I2[4]),
		.B1(out_sel[3]),
		.B2(I3[4]),
		.Z(O1[4])
	);
	AO_CELL inst_2_4(
		.A1(out_sel[4]),
		.A2(I4[4]),
		.B1(out_sel[5]),
		.B2(I5[4]),
		.Z(O2[4])
	);
	AO_CELL inst_3_4(
		.A1(out_sel[6]),
		.A2(I6[4]),
		.B1(out_sel[7]),
		.B2(I7[4]),
		.Z(O3[4])
	);
	AO_CELL inst_4_4(
		.A1(out_sel[8]),
		.A2(I8[4]),
		.B1(out_sel[9]),
		.B2(I9[4]),
		.Z(O4[4])
	);
	AO_CELL inst_5_4(
		.A1(out_sel[10]),
		.A2(I10[4]),
		.B1(out_sel[11]),
		.B2(I11[4]),
		.Z(O5[4])
	);
	AO_CELL inst_6_4(
		.A1(out_sel[12]),
		.A2(I12[4]),
		.B1(out_sel[13]),
		.B2(I13[4]),
		.Z(O6[4])
	);
	AO_CELL inst_7_4(
		.A1(out_sel[14]),
		.A2(I14[4]),
		.B1(out_sel[15]),
		.B2(I15[4]),
		.Z(O7[4])
	);
	AO_CELL inst_8_4(
		.A1(out_sel[16]),
		.A2(I16[4]),
		.B1(out_sel[17]),
		.B2(I17[4]),
		.Z(O8[4])
	);
	AO_CELL inst_9_4(
		.A1(out_sel[18]),
		.A2(I18[4]),
		.B1(out_sel[19]),
		.B2(I19[4]),
		.Z(O9[4])
	);
	AN_CELL inst_and_4(
		.A1(out_sel[20]),
		.A2(1'b0),
		.Z(O10[4])
	);
	AO_CELL inst_0_5(
		.A1(out_sel[0]),
		.A2(I0[5]),
		.B1(out_sel[1]),
		.B2(I1[5]),
		.Z(O0[5])
	);
	AO_CELL inst_1_5(
		.A1(out_sel[2]),
		.A2(I2[5]),
		.B1(out_sel[3]),
		.B2(I3[5]),
		.Z(O1[5])
	);
	AO_CELL inst_2_5(
		.A1(out_sel[4]),
		.A2(I4[5]),
		.B1(out_sel[5]),
		.B2(I5[5]),
		.Z(O2[5])
	);
	AO_CELL inst_3_5(
		.A1(out_sel[6]),
		.A2(I6[5]),
		.B1(out_sel[7]),
		.B2(I7[5]),
		.Z(O3[5])
	);
	AO_CELL inst_4_5(
		.A1(out_sel[8]),
		.A2(I8[5]),
		.B1(out_sel[9]),
		.B2(I9[5]),
		.Z(O4[5])
	);
	AO_CELL inst_5_5(
		.A1(out_sel[10]),
		.A2(I10[5]),
		.B1(out_sel[11]),
		.B2(I11[5]),
		.Z(O5[5])
	);
	AO_CELL inst_6_5(
		.A1(out_sel[12]),
		.A2(I12[5]),
		.B1(out_sel[13]),
		.B2(I13[5]),
		.Z(O6[5])
	);
	AO_CELL inst_7_5(
		.A1(out_sel[14]),
		.A2(I14[5]),
		.B1(out_sel[15]),
		.B2(I15[5]),
		.Z(O7[5])
	);
	AO_CELL inst_8_5(
		.A1(out_sel[16]),
		.A2(I16[5]),
		.B1(out_sel[17]),
		.B2(I17[5]),
		.Z(O8[5])
	);
	AO_CELL inst_9_5(
		.A1(out_sel[18]),
		.A2(I18[5]),
		.B1(out_sel[19]),
		.B2(I19[5]),
		.Z(O9[5])
	);
	AN_CELL inst_and_5(
		.A1(out_sel[20]),
		.A2(1'b0),
		.Z(O10[5])
	);
	AO_CELL inst_0_6(
		.A1(out_sel[0]),
		.A2(I0[6]),
		.B1(out_sel[1]),
		.B2(I1[6]),
		.Z(O0[6])
	);
	AO_CELL inst_1_6(
		.A1(out_sel[2]),
		.A2(I2[6]),
		.B1(out_sel[3]),
		.B2(I3[6]),
		.Z(O1[6])
	);
	AO_CELL inst_2_6(
		.A1(out_sel[4]),
		.A2(I4[6]),
		.B1(out_sel[5]),
		.B2(I5[6]),
		.Z(O2[6])
	);
	AO_CELL inst_3_6(
		.A1(out_sel[6]),
		.A2(I6[6]),
		.B1(out_sel[7]),
		.B2(I7[6]),
		.Z(O3[6])
	);
	AO_CELL inst_4_6(
		.A1(out_sel[8]),
		.A2(I8[6]),
		.B1(out_sel[9]),
		.B2(I9[6]),
		.Z(O4[6])
	);
	AO_CELL inst_5_6(
		.A1(out_sel[10]),
		.A2(I10[6]),
		.B1(out_sel[11]),
		.B2(I11[6]),
		.Z(O5[6])
	);
	AO_CELL inst_6_6(
		.A1(out_sel[12]),
		.A2(I12[6]),
		.B1(out_sel[13]),
		.B2(I13[6]),
		.Z(O6[6])
	);
	AO_CELL inst_7_6(
		.A1(out_sel[14]),
		.A2(I14[6]),
		.B1(out_sel[15]),
		.B2(I15[6]),
		.Z(O7[6])
	);
	AO_CELL inst_8_6(
		.A1(out_sel[16]),
		.A2(I16[6]),
		.B1(out_sel[17]),
		.B2(I17[6]),
		.Z(O8[6])
	);
	AO_CELL inst_9_6(
		.A1(out_sel[18]),
		.A2(I18[6]),
		.B1(out_sel[19]),
		.B2(I19[6]),
		.Z(O9[6])
	);
	AN_CELL inst_and_6(
		.A1(out_sel[20]),
		.A2(1'b0),
		.Z(O10[6])
	);
	AO_CELL inst_0_7(
		.A1(out_sel[0]),
		.A2(I0[7]),
		.B1(out_sel[1]),
		.B2(I1[7]),
		.Z(O0[7])
	);
	AO_CELL inst_1_7(
		.A1(out_sel[2]),
		.A2(I2[7]),
		.B1(out_sel[3]),
		.B2(I3[7]),
		.Z(O1[7])
	);
	AO_CELL inst_2_7(
		.A1(out_sel[4]),
		.A2(I4[7]),
		.B1(out_sel[5]),
		.B2(I5[7]),
		.Z(O2[7])
	);
	AO_CELL inst_3_7(
		.A1(out_sel[6]),
		.A2(I6[7]),
		.B1(out_sel[7]),
		.B2(I7[7]),
		.Z(O3[7])
	);
	AO_CELL inst_4_7(
		.A1(out_sel[8]),
		.A2(I8[7]),
		.B1(out_sel[9]),
		.B2(I9[7]),
		.Z(O4[7])
	);
	AO_CELL inst_5_7(
		.A1(out_sel[10]),
		.A2(I10[7]),
		.B1(out_sel[11]),
		.B2(I11[7]),
		.Z(O5[7])
	);
	AO_CELL inst_6_7(
		.A1(out_sel[12]),
		.A2(I12[7]),
		.B1(out_sel[13]),
		.B2(I13[7]),
		.Z(O6[7])
	);
	AO_CELL inst_7_7(
		.A1(out_sel[14]),
		.A2(I14[7]),
		.B1(out_sel[15]),
		.B2(I15[7]),
		.Z(O7[7])
	);
	AO_CELL inst_8_7(
		.A1(out_sel[16]),
		.A2(I16[7]),
		.B1(out_sel[17]),
		.B2(I17[7]),
		.Z(O8[7])
	);
	AO_CELL inst_9_7(
		.A1(out_sel[18]),
		.A2(I18[7]),
		.B1(out_sel[19]),
		.B2(I19[7]),
		.Z(O9[7])
	);
	AN_CELL inst_and_7(
		.A1(out_sel[20]),
		.A2(1'b0),
		.Z(O10[7])
	);
	AO_CELL inst_0_8(
		.A1(out_sel[0]),
		.A2(I0[8]),
		.B1(out_sel[1]),
		.B2(I1[8]),
		.Z(O0[8])
	);
	AO_CELL inst_1_8(
		.A1(out_sel[2]),
		.A2(I2[8]),
		.B1(out_sel[3]),
		.B2(I3[8]),
		.Z(O1[8])
	);
	AO_CELL inst_2_8(
		.A1(out_sel[4]),
		.A2(I4[8]),
		.B1(out_sel[5]),
		.B2(I5[8]),
		.Z(O2[8])
	);
	AO_CELL inst_3_8(
		.A1(out_sel[6]),
		.A2(I6[8]),
		.B1(out_sel[7]),
		.B2(I7[8]),
		.Z(O3[8])
	);
	AO_CELL inst_4_8(
		.A1(out_sel[8]),
		.A2(I8[8]),
		.B1(out_sel[9]),
		.B2(I9[8]),
		.Z(O4[8])
	);
	AO_CELL inst_5_8(
		.A1(out_sel[10]),
		.A2(I10[8]),
		.B1(out_sel[11]),
		.B2(I11[8]),
		.Z(O5[8])
	);
	AO_CELL inst_6_8(
		.A1(out_sel[12]),
		.A2(I12[8]),
		.B1(out_sel[13]),
		.B2(I13[8]),
		.Z(O6[8])
	);
	AO_CELL inst_7_8(
		.A1(out_sel[14]),
		.A2(I14[8]),
		.B1(out_sel[15]),
		.B2(I15[8]),
		.Z(O7[8])
	);
	AO_CELL inst_8_8(
		.A1(out_sel[16]),
		.A2(I16[8]),
		.B1(out_sel[17]),
		.B2(I17[8]),
		.Z(O8[8])
	);
	AO_CELL inst_9_8(
		.A1(out_sel[18]),
		.A2(I18[8]),
		.B1(out_sel[19]),
		.B2(I19[8]),
		.Z(O9[8])
	);
	AN_CELL inst_and_8(
		.A1(out_sel[20]),
		.A2(1'b0),
		.Z(O10[8])
	);
	AO_CELL inst_0_9(
		.A1(out_sel[0]),
		.A2(I0[9]),
		.B1(out_sel[1]),
		.B2(I1[9]),
		.Z(O0[9])
	);
	AO_CELL inst_1_9(
		.A1(out_sel[2]),
		.A2(I2[9]),
		.B1(out_sel[3]),
		.B2(I3[9]),
		.Z(O1[9])
	);
	AO_CELL inst_2_9(
		.A1(out_sel[4]),
		.A2(I4[9]),
		.B1(out_sel[5]),
		.B2(I5[9]),
		.Z(O2[9])
	);
	AO_CELL inst_3_9(
		.A1(out_sel[6]),
		.A2(I6[9]),
		.B1(out_sel[7]),
		.B2(I7[9]),
		.Z(O3[9])
	);
	AO_CELL inst_4_9(
		.A1(out_sel[8]),
		.A2(I8[9]),
		.B1(out_sel[9]),
		.B2(I9[9]),
		.Z(O4[9])
	);
	AO_CELL inst_5_9(
		.A1(out_sel[10]),
		.A2(I10[9]),
		.B1(out_sel[11]),
		.B2(I11[9]),
		.Z(O5[9])
	);
	AO_CELL inst_6_9(
		.A1(out_sel[12]),
		.A2(I12[9]),
		.B1(out_sel[13]),
		.B2(I13[9]),
		.Z(O6[9])
	);
	AO_CELL inst_7_9(
		.A1(out_sel[14]),
		.A2(I14[9]),
		.B1(out_sel[15]),
		.B2(I15[9]),
		.Z(O7[9])
	);
	AO_CELL inst_8_9(
		.A1(out_sel[16]),
		.A2(I16[9]),
		.B1(out_sel[17]),
		.B2(I17[9]),
		.Z(O8[9])
	);
	AO_CELL inst_9_9(
		.A1(out_sel[18]),
		.A2(I18[9]),
		.B1(out_sel[19]),
		.B2(I19[9]),
		.Z(O9[9])
	);
	AN_CELL inst_and_9(
		.A1(out_sel[20]),
		.A2(1'b0),
		.Z(O10[9])
	);
	AO_CELL inst_0_10(
		.A1(out_sel[0]),
		.A2(I0[10]),
		.B1(out_sel[1]),
		.B2(I1[10]),
		.Z(O0[10])
	);
	AO_CELL inst_1_10(
		.A1(out_sel[2]),
		.A2(I2[10]),
		.B1(out_sel[3]),
		.B2(I3[10]),
		.Z(O1[10])
	);
	AO_CELL inst_2_10(
		.A1(out_sel[4]),
		.A2(I4[10]),
		.B1(out_sel[5]),
		.B2(I5[10]),
		.Z(O2[10])
	);
	AO_CELL inst_3_10(
		.A1(out_sel[6]),
		.A2(I6[10]),
		.B1(out_sel[7]),
		.B2(I7[10]),
		.Z(O3[10])
	);
	AO_CELL inst_4_10(
		.A1(out_sel[8]),
		.A2(I8[10]),
		.B1(out_sel[9]),
		.B2(I9[10]),
		.Z(O4[10])
	);
	AO_CELL inst_5_10(
		.A1(out_sel[10]),
		.A2(I10[10]),
		.B1(out_sel[11]),
		.B2(I11[10]),
		.Z(O5[10])
	);
	AO_CELL inst_6_10(
		.A1(out_sel[12]),
		.A2(I12[10]),
		.B1(out_sel[13]),
		.B2(I13[10]),
		.Z(O6[10])
	);
	AO_CELL inst_7_10(
		.A1(out_sel[14]),
		.A2(I14[10]),
		.B1(out_sel[15]),
		.B2(I15[10]),
		.Z(O7[10])
	);
	AO_CELL inst_8_10(
		.A1(out_sel[16]),
		.A2(I16[10]),
		.B1(out_sel[17]),
		.B2(I17[10]),
		.Z(O8[10])
	);
	AO_CELL inst_9_10(
		.A1(out_sel[18]),
		.A2(I18[10]),
		.B1(out_sel[19]),
		.B2(I19[10]),
		.Z(O9[10])
	);
	AN_CELL inst_and_10(
		.A1(out_sel[20]),
		.A2(1'b0),
		.Z(O10[10])
	);
	AO_CELL inst_0_11(
		.A1(out_sel[0]),
		.A2(I0[11]),
		.B1(out_sel[1]),
		.B2(I1[11]),
		.Z(O0[11])
	);
	AO_CELL inst_1_11(
		.A1(out_sel[2]),
		.A2(I2[11]),
		.B1(out_sel[3]),
		.B2(I3[11]),
		.Z(O1[11])
	);
	AO_CELL inst_2_11(
		.A1(out_sel[4]),
		.A2(I4[11]),
		.B1(out_sel[5]),
		.B2(I5[11]),
		.Z(O2[11])
	);
	AO_CELL inst_3_11(
		.A1(out_sel[6]),
		.A2(I6[11]),
		.B1(out_sel[7]),
		.B2(I7[11]),
		.Z(O3[11])
	);
	AO_CELL inst_4_11(
		.A1(out_sel[8]),
		.A2(I8[11]),
		.B1(out_sel[9]),
		.B2(I9[11]),
		.Z(O4[11])
	);
	AO_CELL inst_5_11(
		.A1(out_sel[10]),
		.A2(I10[11]),
		.B1(out_sel[11]),
		.B2(I11[11]),
		.Z(O5[11])
	);
	AO_CELL inst_6_11(
		.A1(out_sel[12]),
		.A2(I12[11]),
		.B1(out_sel[13]),
		.B2(I13[11]),
		.Z(O6[11])
	);
	AO_CELL inst_7_11(
		.A1(out_sel[14]),
		.A2(I14[11]),
		.B1(out_sel[15]),
		.B2(I15[11]),
		.Z(O7[11])
	);
	AO_CELL inst_8_11(
		.A1(out_sel[16]),
		.A2(I16[11]),
		.B1(out_sel[17]),
		.B2(I17[11]),
		.Z(O8[11])
	);
	AO_CELL inst_9_11(
		.A1(out_sel[18]),
		.A2(I18[11]),
		.B1(out_sel[19]),
		.B2(I19[11]),
		.Z(O9[11])
	);
	AN_CELL inst_and_11(
		.A1(out_sel[20]),
		.A2(1'b0),
		.Z(O10[11])
	);
	AO_CELL inst_0_12(
		.A1(out_sel[0]),
		.A2(I0[12]),
		.B1(out_sel[1]),
		.B2(I1[12]),
		.Z(O0[12])
	);
	AO_CELL inst_1_12(
		.A1(out_sel[2]),
		.A2(I2[12]),
		.B1(out_sel[3]),
		.B2(I3[12]),
		.Z(O1[12])
	);
	AO_CELL inst_2_12(
		.A1(out_sel[4]),
		.A2(I4[12]),
		.B1(out_sel[5]),
		.B2(I5[12]),
		.Z(O2[12])
	);
	AO_CELL inst_3_12(
		.A1(out_sel[6]),
		.A2(I6[12]),
		.B1(out_sel[7]),
		.B2(I7[12]),
		.Z(O3[12])
	);
	AO_CELL inst_4_12(
		.A1(out_sel[8]),
		.A2(I8[12]),
		.B1(out_sel[9]),
		.B2(I9[12]),
		.Z(O4[12])
	);
	AO_CELL inst_5_12(
		.A1(out_sel[10]),
		.A2(I10[12]),
		.B1(out_sel[11]),
		.B2(I11[12]),
		.Z(O5[12])
	);
	AO_CELL inst_6_12(
		.A1(out_sel[12]),
		.A2(I12[12]),
		.B1(out_sel[13]),
		.B2(I13[12]),
		.Z(O6[12])
	);
	AO_CELL inst_7_12(
		.A1(out_sel[14]),
		.A2(I14[12]),
		.B1(out_sel[15]),
		.B2(I15[12]),
		.Z(O7[12])
	);
	AO_CELL inst_8_12(
		.A1(out_sel[16]),
		.A2(I16[12]),
		.B1(out_sel[17]),
		.B2(I17[12]),
		.Z(O8[12])
	);
	AO_CELL inst_9_12(
		.A1(out_sel[18]),
		.A2(I18[12]),
		.B1(out_sel[19]),
		.B2(I19[12]),
		.Z(O9[12])
	);
	AN_CELL inst_and_12(
		.A1(out_sel[20]),
		.A2(1'b0),
		.Z(O10[12])
	);
	AO_CELL inst_0_13(
		.A1(out_sel[0]),
		.A2(I0[13]),
		.B1(out_sel[1]),
		.B2(I1[13]),
		.Z(O0[13])
	);
	AO_CELL inst_1_13(
		.A1(out_sel[2]),
		.A2(I2[13]),
		.B1(out_sel[3]),
		.B2(I3[13]),
		.Z(O1[13])
	);
	AO_CELL inst_2_13(
		.A1(out_sel[4]),
		.A2(I4[13]),
		.B1(out_sel[5]),
		.B2(I5[13]),
		.Z(O2[13])
	);
	AO_CELL inst_3_13(
		.A1(out_sel[6]),
		.A2(I6[13]),
		.B1(out_sel[7]),
		.B2(I7[13]),
		.Z(O3[13])
	);
	AO_CELL inst_4_13(
		.A1(out_sel[8]),
		.A2(I8[13]),
		.B1(out_sel[9]),
		.B2(I9[13]),
		.Z(O4[13])
	);
	AO_CELL inst_5_13(
		.A1(out_sel[10]),
		.A2(I10[13]),
		.B1(out_sel[11]),
		.B2(I11[13]),
		.Z(O5[13])
	);
	AO_CELL inst_6_13(
		.A1(out_sel[12]),
		.A2(I12[13]),
		.B1(out_sel[13]),
		.B2(I13[13]),
		.Z(O6[13])
	);
	AO_CELL inst_7_13(
		.A1(out_sel[14]),
		.A2(I14[13]),
		.B1(out_sel[15]),
		.B2(I15[13]),
		.Z(O7[13])
	);
	AO_CELL inst_8_13(
		.A1(out_sel[16]),
		.A2(I16[13]),
		.B1(out_sel[17]),
		.B2(I17[13]),
		.Z(O8[13])
	);
	AO_CELL inst_9_13(
		.A1(out_sel[18]),
		.A2(I18[13]),
		.B1(out_sel[19]),
		.B2(I19[13]),
		.Z(O9[13])
	);
	AN_CELL inst_and_13(
		.A1(out_sel[20]),
		.A2(1'b0),
		.Z(O10[13])
	);
	AO_CELL inst_0_14(
		.A1(out_sel[0]),
		.A2(I0[14]),
		.B1(out_sel[1]),
		.B2(I1[14]),
		.Z(O0[14])
	);
	AO_CELL inst_1_14(
		.A1(out_sel[2]),
		.A2(I2[14]),
		.B1(out_sel[3]),
		.B2(I3[14]),
		.Z(O1[14])
	);
	AO_CELL inst_2_14(
		.A1(out_sel[4]),
		.A2(I4[14]),
		.B1(out_sel[5]),
		.B2(I5[14]),
		.Z(O2[14])
	);
	AO_CELL inst_3_14(
		.A1(out_sel[6]),
		.A2(I6[14]),
		.B1(out_sel[7]),
		.B2(I7[14]),
		.Z(O3[14])
	);
	AO_CELL inst_4_14(
		.A1(out_sel[8]),
		.A2(I8[14]),
		.B1(out_sel[9]),
		.B2(I9[14]),
		.Z(O4[14])
	);
	AO_CELL inst_5_14(
		.A1(out_sel[10]),
		.A2(I10[14]),
		.B1(out_sel[11]),
		.B2(I11[14]),
		.Z(O5[14])
	);
	AO_CELL inst_6_14(
		.A1(out_sel[12]),
		.A2(I12[14]),
		.B1(out_sel[13]),
		.B2(I13[14]),
		.Z(O6[14])
	);
	AO_CELL inst_7_14(
		.A1(out_sel[14]),
		.A2(I14[14]),
		.B1(out_sel[15]),
		.B2(I15[14]),
		.Z(O7[14])
	);
	AO_CELL inst_8_14(
		.A1(out_sel[16]),
		.A2(I16[14]),
		.B1(out_sel[17]),
		.B2(I17[14]),
		.Z(O8[14])
	);
	AO_CELL inst_9_14(
		.A1(out_sel[18]),
		.A2(I18[14]),
		.B1(out_sel[19]),
		.B2(I19[14]),
		.Z(O9[14])
	);
	AN_CELL inst_and_14(
		.A1(out_sel[20]),
		.A2(1'b0),
		.Z(O10[14])
	);
	AO_CELL inst_0_15(
		.A1(out_sel[0]),
		.A2(I0[15]),
		.B1(out_sel[1]),
		.B2(I1[15]),
		.Z(O0[15])
	);
	AO_CELL inst_1_15(
		.A1(out_sel[2]),
		.A2(I2[15]),
		.B1(out_sel[3]),
		.B2(I3[15]),
		.Z(O1[15])
	);
	AO_CELL inst_2_15(
		.A1(out_sel[4]),
		.A2(I4[15]),
		.B1(out_sel[5]),
		.B2(I5[15]),
		.Z(O2[15])
	);
	AO_CELL inst_3_15(
		.A1(out_sel[6]),
		.A2(I6[15]),
		.B1(out_sel[7]),
		.B2(I7[15]),
		.Z(O3[15])
	);
	AO_CELL inst_4_15(
		.A1(out_sel[8]),
		.A2(I8[15]),
		.B1(out_sel[9]),
		.B2(I9[15]),
		.Z(O4[15])
	);
	AO_CELL inst_5_15(
		.A1(out_sel[10]),
		.A2(I10[15]),
		.B1(out_sel[11]),
		.B2(I11[15]),
		.Z(O5[15])
	);
	AO_CELL inst_6_15(
		.A1(out_sel[12]),
		.A2(I12[15]),
		.B1(out_sel[13]),
		.B2(I13[15]),
		.Z(O6[15])
	);
	AO_CELL inst_7_15(
		.A1(out_sel[14]),
		.A2(I14[15]),
		.B1(out_sel[15]),
		.B2(I15[15]),
		.Z(O7[15])
	);
	AO_CELL inst_8_15(
		.A1(out_sel[16]),
		.A2(I16[15]),
		.B1(out_sel[17]),
		.B2(I17[15]),
		.Z(O8[15])
	);
	AO_CELL inst_9_15(
		.A1(out_sel[18]),
		.A2(I18[15]),
		.B1(out_sel[19]),
		.B2(I19[15]),
		.Z(O9[15])
	);
	AN_CELL inst_and_15(
		.A1(out_sel[20]),
		.A2(1'b0),
		.Z(O10[15])
	);
	AO_CELL inst_0_16(
		.A1(out_sel[0]),
		.A2(I0[16]),
		.B1(out_sel[1]),
		.B2(I1[16]),
		.Z(O0[16])
	);
	AO_CELL inst_1_16(
		.A1(out_sel[2]),
		.A2(I2[16]),
		.B1(out_sel[3]),
		.B2(I3[16]),
		.Z(O1[16])
	);
	AO_CELL inst_2_16(
		.A1(out_sel[4]),
		.A2(I4[16]),
		.B1(out_sel[5]),
		.B2(I5[16]),
		.Z(O2[16])
	);
	AO_CELL inst_3_16(
		.A1(out_sel[6]),
		.A2(I6[16]),
		.B1(out_sel[7]),
		.B2(I7[16]),
		.Z(O3[16])
	);
	AO_CELL inst_4_16(
		.A1(out_sel[8]),
		.A2(I8[16]),
		.B1(out_sel[9]),
		.B2(I9[16]),
		.Z(O4[16])
	);
	AO_CELL inst_5_16(
		.A1(out_sel[10]),
		.A2(I10[16]),
		.B1(out_sel[11]),
		.B2(I11[16]),
		.Z(O5[16])
	);
	AO_CELL inst_6_16(
		.A1(out_sel[12]),
		.A2(I12[16]),
		.B1(out_sel[13]),
		.B2(I13[16]),
		.Z(O6[16])
	);
	AO_CELL inst_7_16(
		.A1(out_sel[14]),
		.A2(I14[16]),
		.B1(out_sel[15]),
		.B2(I15[16]),
		.Z(O7[16])
	);
	AO_CELL inst_8_16(
		.A1(out_sel[16]),
		.A2(I16[16]),
		.B1(out_sel[17]),
		.B2(I17[16]),
		.Z(O8[16])
	);
	AO_CELL inst_9_16(
		.A1(out_sel[18]),
		.A2(I18[16]),
		.B1(out_sel[19]),
		.B2(I19[16]),
		.Z(O9[16])
	);
	AN_CELL inst_and_16(
		.A1(out_sel[20]),
		.A2(1'b0),
		.Z(O10[16])
	);
	AO_CELL inst_0_valid(
		.A1(out_sel[0]),
		.A2(valid_in[0]),
		.B1(out_sel[1]),
		.B2(valid_in[1]),
		.Z(valid_out[0])
	);
	AO_CELL inst_1_valid(
		.A1(out_sel[2]),
		.A2(valid_in[2]),
		.B1(out_sel[3]),
		.B2(valid_in[3]),
		.Z(valid_out[1])
	);
	AO_CELL inst_2_valid(
		.A1(out_sel[4]),
		.A2(valid_in[4]),
		.B1(out_sel[5]),
		.B2(valid_in[5]),
		.Z(valid_out[2])
	);
	AO_CELL inst_3_valid(
		.A1(out_sel[6]),
		.A2(valid_in[6]),
		.B1(out_sel[7]),
		.B2(valid_in[7]),
		.Z(valid_out[3])
	);
	AO_CELL inst_4_valid(
		.A1(out_sel[8]),
		.A2(valid_in[8]),
		.B1(out_sel[9]),
		.B2(valid_in[9]),
		.Z(valid_out[4])
	);
	AO_CELL inst_5_valid(
		.A1(out_sel[10]),
		.A2(valid_in[10]),
		.B1(out_sel[11]),
		.B2(valid_in[11]),
		.Z(valid_out[5])
	);
	AO_CELL inst_6_valid(
		.A1(out_sel[12]),
		.A2(valid_in[12]),
		.B1(out_sel[13]),
		.B2(valid_in[13]),
		.Z(valid_out[6])
	);
	AO_CELL inst_7_valid(
		.A1(out_sel[14]),
		.A2(valid_in[14]),
		.B1(out_sel[15]),
		.B2(valid_in[15]),
		.Z(valid_out[7])
	);
	AO_CELL inst_8_valid(
		.A1(out_sel[16]),
		.A2(valid_in[16]),
		.B1(out_sel[17]),
		.B2(valid_in[17]),
		.Z(valid_out[8])
	);
	AO_CELL inst_9_valid(
		.A1(out_sel[18]),
		.A2(valid_in[18]),
		.B1(out_sel[19]),
		.B2(valid_in[19]),
		.Z(valid_out[9])
	);
	AN_CELL inst_and_10_valid(
		.A1(out_sel[20]),
		.A2(1'b0),
		.Z(valid_out[10])
	);
endmodule
module mux_aoi_ready_valid_const_20_1 (
	I,
	S,
	ready_in,
	ready_out,
	valid_in,
	valid_out,
	out_sel,
	O
);
	input wire [19:0] I;
	input wire [4:0] S;
	input wire ready_in;
	output wire ready_out;
	input wire [19:0] valid_in;
	output wire valid_out;
	output wire [31:0] out_sel;
	output wire [0:0] O;
	wire [0:0] O_int0;
	wire [0:0] O_int1;
	wire [0:0] O_int2;
	wire [0:0] O_int3;
	wire [0:0] O_int4;
	wire [0:0] O_int5;
	wire [0:0] O_int6;
	wire [0:0] O_int7;
	wire [0:0] O_int8;
	wire [0:0] O_int9;
	wire [0:0] O_int10;
	wire [10:0] valid_out_temp;
	precoder_1_20 u_precoder(
		.S(S),
		.out_sel(out_sel)
	);
	mux_logic_1_20 u_mux_logic(
		.I0(I[0+:1]),
		.I1(I[1+:1]),
		.I2(I[2+:1]),
		.I3(I[3+:1]),
		.I4(I[4+:1]),
		.I5(I[5+:1]),
		.I6(I[6+:1]),
		.I7(I[7+:1]),
		.I8(I[8+:1]),
		.I9(I[9+:1]),
		.I10(I[10+:1]),
		.I11(I[11+:1]),
		.I12(I[12+:1]),
		.I13(I[13+:1]),
		.I14(I[14+:1]),
		.I15(I[15+:1]),
		.I16(I[16+:1]),
		.I17(I[17+:1]),
		.I18(I[18+:1]),
		.I19(I[19+:1]),
		.out_sel(out_sel),
		.valid_in(valid_in),
		.valid_out(valid_out_temp),
		.O0(O_int0),
		.O1(O_int1),
		.O2(O_int2),
		.O3(O_int3),
		.O4(O_int4),
		.O5(O_int5),
		.O6(O_int6),
		.O7(O_int7),
		.O8(O_int8),
		.O9(O_int9),
		.O10(O_int10)
	);
	assign O = (((((((((O_int0 | O_int1) | O_int2) | O_int3) | O_int4) | O_int5) | O_int6) | O_int7) | O_int8) | O_int9) | O_int10;
	assign ready_out = ready_in;
	assign valid_out = |valid_out_temp;
endmodule
module precoder_1_20 (
	S,
	out_sel
);
	input wire [4:0] S;
	output reg [31:0] out_sel;
	always @(*) begin : mux_sel
		case (S)
			5'd0: out_sel = 32'b00000000000000000000000000000001;
			5'd1: out_sel = 32'b00000000000000000000000000000010;
			5'd2: out_sel = 32'b00000000000000000000000000000100;
			5'd3: out_sel = 32'b00000000000000000000000000001000;
			5'd4: out_sel = 32'b00000000000000000000000000010000;
			5'd5: out_sel = 32'b00000000000000000000000000100000;
			5'd6: out_sel = 32'b00000000000000000000000001000000;
			5'd7: out_sel = 32'b00000000000000000000000010000000;
			5'd8: out_sel = 32'b00000000000000000000000100000000;
			5'd9: out_sel = 32'b00000000000000000000001000000000;
			5'd10: out_sel = 32'b00000000000000000000010000000000;
			5'd11: out_sel = 32'b00000000000000000000100000000000;
			5'd12: out_sel = 32'b00000000000000000001000000000000;
			5'd13: out_sel = 32'b00000000000000000010000000000000;
			5'd14: out_sel = 32'b00000000000000000100000000000000;
			5'd15: out_sel = 32'b00000000000000001000000000000000;
			5'd16: out_sel = 32'b00000000000000010000000000000000;
			5'd17: out_sel = 32'b00000000000000100000000000000000;
			5'd18: out_sel = 32'b00000000000001000000000000000000;
			5'd19: out_sel = 32'b00000000000010000000000000000000;
			5'd20: out_sel = 32'b00000000000100000000000000000000;
			default: out_sel = 32'b00000000000000000000000000000000;
		endcase
	end
endmodule
module mux_logic_1_20 (
	out_sel,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	I9,
	I10,
	I11,
	I12,
	I13,
	I14,
	I15,
	I16,
	I17,
	I18,
	I19,
	valid_in,
	valid_out,
	O0,
	O1,
	O2,
	O3,
	O4,
	O5,
	O6,
	O7,
	O8,
	O9,
	O10
);
	input wire [31:0] out_sel;
	input wire [0:0] I0;
	input wire [0:0] I1;
	input wire [0:0] I2;
	input wire [0:0] I3;
	input wire [0:0] I4;
	input wire [0:0] I5;
	input wire [0:0] I6;
	input wire [0:0] I7;
	input wire [0:0] I8;
	input wire [0:0] I9;
	input wire [0:0] I10;
	input wire [0:0] I11;
	input wire [0:0] I12;
	input wire [0:0] I13;
	input wire [0:0] I14;
	input wire [0:0] I15;
	input wire [0:0] I16;
	input wire [0:0] I17;
	input wire [0:0] I18;
	input wire [0:0] I19;
	input wire [19:0] valid_in;
	output wire [10:0] valid_out;
	output wire [0:0] O0;
	output wire [0:0] O1;
	output wire [0:0] O2;
	output wire [0:0] O3;
	output wire [0:0] O4;
	output wire [0:0] O5;
	output wire [0:0] O6;
	output wire [0:0] O7;
	output wire [0:0] O8;
	output wire [0:0] O9;
	output wire [0:0] O10;
	AO_CELL inst_0_0(
		.A1(out_sel[0]),
		.A2(I0[0]),
		.B1(out_sel[1]),
		.B2(I1[0]),
		.Z(O0[0])
	);
	AO_CELL inst_1_0(
		.A1(out_sel[2]),
		.A2(I2[0]),
		.B1(out_sel[3]),
		.B2(I3[0]),
		.Z(O1[0])
	);
	AO_CELL inst_2_0(
		.A1(out_sel[4]),
		.A2(I4[0]),
		.B1(out_sel[5]),
		.B2(I5[0]),
		.Z(O2[0])
	);
	AO_CELL inst_3_0(
		.A1(out_sel[6]),
		.A2(I6[0]),
		.B1(out_sel[7]),
		.B2(I7[0]),
		.Z(O3[0])
	);
	AO_CELL inst_4_0(
		.A1(out_sel[8]),
		.A2(I8[0]),
		.B1(out_sel[9]),
		.B2(I9[0]),
		.Z(O4[0])
	);
	AO_CELL inst_5_0(
		.A1(out_sel[10]),
		.A2(I10[0]),
		.B1(out_sel[11]),
		.B2(I11[0]),
		.Z(O5[0])
	);
	AO_CELL inst_6_0(
		.A1(out_sel[12]),
		.A2(I12[0]),
		.B1(out_sel[13]),
		.B2(I13[0]),
		.Z(O6[0])
	);
	AO_CELL inst_7_0(
		.A1(out_sel[14]),
		.A2(I14[0]),
		.B1(out_sel[15]),
		.B2(I15[0]),
		.Z(O7[0])
	);
	AO_CELL inst_8_0(
		.A1(out_sel[16]),
		.A2(I16[0]),
		.B1(out_sel[17]),
		.B2(I17[0]),
		.Z(O8[0])
	);
	AO_CELL inst_9_0(
		.A1(out_sel[18]),
		.A2(I18[0]),
		.B1(out_sel[19]),
		.B2(I19[0]),
		.Z(O9[0])
	);
	AN_CELL inst_and_0(
		.A1(out_sel[20]),
		.A2(1'b0),
		.Z(O10[0])
	);
	AO_CELL inst_0_valid(
		.A1(out_sel[0]),
		.A2(valid_in[0]),
		.B1(out_sel[1]),
		.B2(valid_in[1]),
		.Z(valid_out[0])
	);
	AO_CELL inst_1_valid(
		.A1(out_sel[2]),
		.A2(valid_in[2]),
		.B1(out_sel[3]),
		.B2(valid_in[3]),
		.Z(valid_out[1])
	);
	AO_CELL inst_2_valid(
		.A1(out_sel[4]),
		.A2(valid_in[4]),
		.B1(out_sel[5]),
		.B2(valid_in[5]),
		.Z(valid_out[2])
	);
	AO_CELL inst_3_valid(
		.A1(out_sel[6]),
		.A2(valid_in[6]),
		.B1(out_sel[7]),
		.B2(valid_in[7]),
		.Z(valid_out[3])
	);
	AO_CELL inst_4_valid(
		.A1(out_sel[8]),
		.A2(valid_in[8]),
		.B1(out_sel[9]),
		.B2(valid_in[9]),
		.Z(valid_out[4])
	);
	AO_CELL inst_5_valid(
		.A1(out_sel[10]),
		.A2(valid_in[10]),
		.B1(out_sel[11]),
		.B2(valid_in[11]),
		.Z(valid_out[5])
	);
	AO_CELL inst_6_valid(
		.A1(out_sel[12]),
		.A2(valid_in[12]),
		.B1(out_sel[13]),
		.B2(valid_in[13]),
		.Z(valid_out[6])
	);
	AO_CELL inst_7_valid(
		.A1(out_sel[14]),
		.A2(valid_in[14]),
		.B1(out_sel[15]),
		.B2(valid_in[15]),
		.Z(valid_out[7])
	);
	AO_CELL inst_8_valid(
		.A1(out_sel[16]),
		.A2(valid_in[16]),
		.B1(out_sel[17]),
		.B2(valid_in[17]),
		.Z(valid_out[8])
	);
	AO_CELL inst_9_valid(
		.A1(out_sel[18]),
		.A2(valid_in[18]),
		.B1(out_sel[19]),
		.B2(valid_in[19]),
		.Z(valid_out[9])
	);
	AN_CELL inst_and_10_valid(
		.A1(out_sel[20]),
		.A2(1'b0),
		.Z(valid_out[10])
	);
endmodule
module mux_aoi_ready_valid_7_17 (
	I,
	S,
	ready_in,
	ready_out,
	valid_in,
	valid_out,
	out_sel,
	O
);
	input wire [118:0] I;
	input wire [2:0] S;
	input wire ready_in;
	output wire ready_out;
	input wire [6:0] valid_in;
	output wire valid_out;
	output wire [7:0] out_sel;
	output wire [16:0] O;
	wire [16:0] O_int0;
	wire [16:0] O_int1;
	wire [16:0] O_int2;
	wire [16:0] O_int3;
	wire [3:0] valid_out_temp;
	precoder_17_7 u_precoder(
		.S(S),
		.out_sel(out_sel)
	);
	mux_logic_17_7 u_mux_logic(
		.I0(I[0+:17]),
		.I1(I[17+:17]),
		.I2(I[34+:17]),
		.I3(I[51+:17]),
		.I4(I[68+:17]),
		.I5(I[85+:17]),
		.I6(I[102+:17]),
		.out_sel(out_sel),
		.valid_in(valid_in),
		.valid_out(valid_out_temp),
		.O0(O_int0),
		.O1(O_int1),
		.O2(O_int2),
		.O3(O_int3)
	);
	assign O = ((O_int0 | O_int1) | O_int2) | O_int3;
	assign ready_out = ready_in;
	assign valid_out = |valid_out_temp;
endmodule
module precoder_17_7 (
	S,
	out_sel
);
	input wire [2:0] S;
	output reg [7:0] out_sel;
	always @(*) begin : mux_sel
		case (S)
			3'd0: out_sel = 8'b00000001;
			3'd1: out_sel = 8'b00000010;
			3'd2: out_sel = 8'b00000100;
			3'd3: out_sel = 8'b00001000;
			3'd4: out_sel = 8'b00010000;
			3'd5: out_sel = 8'b00100000;
			3'd6: out_sel = 8'b01000000;
			default: out_sel = 8'b00000000;
		endcase
	end
endmodule
module mux_logic_17_7 (
	out_sel,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	valid_in,
	valid_out,
	O0,
	O1,
	O2,
	O3
);
	input wire [7:0] out_sel;
	input wire [16:0] I0;
	input wire [16:0] I1;
	input wire [16:0] I2;
	input wire [16:0] I3;
	input wire [16:0] I4;
	input wire [16:0] I5;
	input wire [16:0] I6;
	input wire [6:0] valid_in;
	output wire [3:0] valid_out;
	output wire [16:0] O0;
	output wire [16:0] O1;
	output wire [16:0] O2;
	output wire [16:0] O3;
	AO_CELL inst_0_0(
		.A1(out_sel[0]),
		.A2(I0[0]),
		.B1(out_sel[1]),
		.B2(I1[0]),
		.Z(O0[0])
	);
	AO_CELL inst_1_0(
		.A1(out_sel[2]),
		.A2(I2[0]),
		.B1(out_sel[3]),
		.B2(I3[0]),
		.Z(O1[0])
	);
	AO_CELL inst_2_0(
		.A1(out_sel[4]),
		.A2(I4[0]),
		.B1(out_sel[5]),
		.B2(I5[0]),
		.Z(O2[0])
	);
	AN_CELL inst_and_0(
		.A1(out_sel[6]),
		.A2(I6[0]),
		.Z(O3[0])
	);
	AO_CELL inst_0_1(
		.A1(out_sel[0]),
		.A2(I0[1]),
		.B1(out_sel[1]),
		.B2(I1[1]),
		.Z(O0[1])
	);
	AO_CELL inst_1_1(
		.A1(out_sel[2]),
		.A2(I2[1]),
		.B1(out_sel[3]),
		.B2(I3[1]),
		.Z(O1[1])
	);
	AO_CELL inst_2_1(
		.A1(out_sel[4]),
		.A2(I4[1]),
		.B1(out_sel[5]),
		.B2(I5[1]),
		.Z(O2[1])
	);
	AN_CELL inst_and_1(
		.A1(out_sel[6]),
		.A2(I6[1]),
		.Z(O3[1])
	);
	AO_CELL inst_0_2(
		.A1(out_sel[0]),
		.A2(I0[2]),
		.B1(out_sel[1]),
		.B2(I1[2]),
		.Z(O0[2])
	);
	AO_CELL inst_1_2(
		.A1(out_sel[2]),
		.A2(I2[2]),
		.B1(out_sel[3]),
		.B2(I3[2]),
		.Z(O1[2])
	);
	AO_CELL inst_2_2(
		.A1(out_sel[4]),
		.A2(I4[2]),
		.B1(out_sel[5]),
		.B2(I5[2]),
		.Z(O2[2])
	);
	AN_CELL inst_and_2(
		.A1(out_sel[6]),
		.A2(I6[2]),
		.Z(O3[2])
	);
	AO_CELL inst_0_3(
		.A1(out_sel[0]),
		.A2(I0[3]),
		.B1(out_sel[1]),
		.B2(I1[3]),
		.Z(O0[3])
	);
	AO_CELL inst_1_3(
		.A1(out_sel[2]),
		.A2(I2[3]),
		.B1(out_sel[3]),
		.B2(I3[3]),
		.Z(O1[3])
	);
	AO_CELL inst_2_3(
		.A1(out_sel[4]),
		.A2(I4[3]),
		.B1(out_sel[5]),
		.B2(I5[3]),
		.Z(O2[3])
	);
	AN_CELL inst_and_3(
		.A1(out_sel[6]),
		.A2(I6[3]),
		.Z(O3[3])
	);
	AO_CELL inst_0_4(
		.A1(out_sel[0]),
		.A2(I0[4]),
		.B1(out_sel[1]),
		.B2(I1[4]),
		.Z(O0[4])
	);
	AO_CELL inst_1_4(
		.A1(out_sel[2]),
		.A2(I2[4]),
		.B1(out_sel[3]),
		.B2(I3[4]),
		.Z(O1[4])
	);
	AO_CELL inst_2_4(
		.A1(out_sel[4]),
		.A2(I4[4]),
		.B1(out_sel[5]),
		.B2(I5[4]),
		.Z(O2[4])
	);
	AN_CELL inst_and_4(
		.A1(out_sel[6]),
		.A2(I6[4]),
		.Z(O3[4])
	);
	AO_CELL inst_0_5(
		.A1(out_sel[0]),
		.A2(I0[5]),
		.B1(out_sel[1]),
		.B2(I1[5]),
		.Z(O0[5])
	);
	AO_CELL inst_1_5(
		.A1(out_sel[2]),
		.A2(I2[5]),
		.B1(out_sel[3]),
		.B2(I3[5]),
		.Z(O1[5])
	);
	AO_CELL inst_2_5(
		.A1(out_sel[4]),
		.A2(I4[5]),
		.B1(out_sel[5]),
		.B2(I5[5]),
		.Z(O2[5])
	);
	AN_CELL inst_and_5(
		.A1(out_sel[6]),
		.A2(I6[5]),
		.Z(O3[5])
	);
	AO_CELL inst_0_6(
		.A1(out_sel[0]),
		.A2(I0[6]),
		.B1(out_sel[1]),
		.B2(I1[6]),
		.Z(O0[6])
	);
	AO_CELL inst_1_6(
		.A1(out_sel[2]),
		.A2(I2[6]),
		.B1(out_sel[3]),
		.B2(I3[6]),
		.Z(O1[6])
	);
	AO_CELL inst_2_6(
		.A1(out_sel[4]),
		.A2(I4[6]),
		.B1(out_sel[5]),
		.B2(I5[6]),
		.Z(O2[6])
	);
	AN_CELL inst_and_6(
		.A1(out_sel[6]),
		.A2(I6[6]),
		.Z(O3[6])
	);
	AO_CELL inst_0_7(
		.A1(out_sel[0]),
		.A2(I0[7]),
		.B1(out_sel[1]),
		.B2(I1[7]),
		.Z(O0[7])
	);
	AO_CELL inst_1_7(
		.A1(out_sel[2]),
		.A2(I2[7]),
		.B1(out_sel[3]),
		.B2(I3[7]),
		.Z(O1[7])
	);
	AO_CELL inst_2_7(
		.A1(out_sel[4]),
		.A2(I4[7]),
		.B1(out_sel[5]),
		.B2(I5[7]),
		.Z(O2[7])
	);
	AN_CELL inst_and_7(
		.A1(out_sel[6]),
		.A2(I6[7]),
		.Z(O3[7])
	);
	AO_CELL inst_0_8(
		.A1(out_sel[0]),
		.A2(I0[8]),
		.B1(out_sel[1]),
		.B2(I1[8]),
		.Z(O0[8])
	);
	AO_CELL inst_1_8(
		.A1(out_sel[2]),
		.A2(I2[8]),
		.B1(out_sel[3]),
		.B2(I3[8]),
		.Z(O1[8])
	);
	AO_CELL inst_2_8(
		.A1(out_sel[4]),
		.A2(I4[8]),
		.B1(out_sel[5]),
		.B2(I5[8]),
		.Z(O2[8])
	);
	AN_CELL inst_and_8(
		.A1(out_sel[6]),
		.A2(I6[8]),
		.Z(O3[8])
	);
	AO_CELL inst_0_9(
		.A1(out_sel[0]),
		.A2(I0[9]),
		.B1(out_sel[1]),
		.B2(I1[9]),
		.Z(O0[9])
	);
	AO_CELL inst_1_9(
		.A1(out_sel[2]),
		.A2(I2[9]),
		.B1(out_sel[3]),
		.B2(I3[9]),
		.Z(O1[9])
	);
	AO_CELL inst_2_9(
		.A1(out_sel[4]),
		.A2(I4[9]),
		.B1(out_sel[5]),
		.B2(I5[9]),
		.Z(O2[9])
	);
	AN_CELL inst_and_9(
		.A1(out_sel[6]),
		.A2(I6[9]),
		.Z(O3[9])
	);
	AO_CELL inst_0_10(
		.A1(out_sel[0]),
		.A2(I0[10]),
		.B1(out_sel[1]),
		.B2(I1[10]),
		.Z(O0[10])
	);
	AO_CELL inst_1_10(
		.A1(out_sel[2]),
		.A2(I2[10]),
		.B1(out_sel[3]),
		.B2(I3[10]),
		.Z(O1[10])
	);
	AO_CELL inst_2_10(
		.A1(out_sel[4]),
		.A2(I4[10]),
		.B1(out_sel[5]),
		.B2(I5[10]),
		.Z(O2[10])
	);
	AN_CELL inst_and_10(
		.A1(out_sel[6]),
		.A2(I6[10]),
		.Z(O3[10])
	);
	AO_CELL inst_0_11(
		.A1(out_sel[0]),
		.A2(I0[11]),
		.B1(out_sel[1]),
		.B2(I1[11]),
		.Z(O0[11])
	);
	AO_CELL inst_1_11(
		.A1(out_sel[2]),
		.A2(I2[11]),
		.B1(out_sel[3]),
		.B2(I3[11]),
		.Z(O1[11])
	);
	AO_CELL inst_2_11(
		.A1(out_sel[4]),
		.A2(I4[11]),
		.B1(out_sel[5]),
		.B2(I5[11]),
		.Z(O2[11])
	);
	AN_CELL inst_and_11(
		.A1(out_sel[6]),
		.A2(I6[11]),
		.Z(O3[11])
	);
	AO_CELL inst_0_12(
		.A1(out_sel[0]),
		.A2(I0[12]),
		.B1(out_sel[1]),
		.B2(I1[12]),
		.Z(O0[12])
	);
	AO_CELL inst_1_12(
		.A1(out_sel[2]),
		.A2(I2[12]),
		.B1(out_sel[3]),
		.B2(I3[12]),
		.Z(O1[12])
	);
	AO_CELL inst_2_12(
		.A1(out_sel[4]),
		.A2(I4[12]),
		.B1(out_sel[5]),
		.B2(I5[12]),
		.Z(O2[12])
	);
	AN_CELL inst_and_12(
		.A1(out_sel[6]),
		.A2(I6[12]),
		.Z(O3[12])
	);
	AO_CELL inst_0_13(
		.A1(out_sel[0]),
		.A2(I0[13]),
		.B1(out_sel[1]),
		.B2(I1[13]),
		.Z(O0[13])
	);
	AO_CELL inst_1_13(
		.A1(out_sel[2]),
		.A2(I2[13]),
		.B1(out_sel[3]),
		.B2(I3[13]),
		.Z(O1[13])
	);
	AO_CELL inst_2_13(
		.A1(out_sel[4]),
		.A2(I4[13]),
		.B1(out_sel[5]),
		.B2(I5[13]),
		.Z(O2[13])
	);
	AN_CELL inst_and_13(
		.A1(out_sel[6]),
		.A2(I6[13]),
		.Z(O3[13])
	);
	AO_CELL inst_0_14(
		.A1(out_sel[0]),
		.A2(I0[14]),
		.B1(out_sel[1]),
		.B2(I1[14]),
		.Z(O0[14])
	);
	AO_CELL inst_1_14(
		.A1(out_sel[2]),
		.A2(I2[14]),
		.B1(out_sel[3]),
		.B2(I3[14]),
		.Z(O1[14])
	);
	AO_CELL inst_2_14(
		.A1(out_sel[4]),
		.A2(I4[14]),
		.B1(out_sel[5]),
		.B2(I5[14]),
		.Z(O2[14])
	);
	AN_CELL inst_and_14(
		.A1(out_sel[6]),
		.A2(I6[14]),
		.Z(O3[14])
	);
	AO_CELL inst_0_15(
		.A1(out_sel[0]),
		.A2(I0[15]),
		.B1(out_sel[1]),
		.B2(I1[15]),
		.Z(O0[15])
	);
	AO_CELL inst_1_15(
		.A1(out_sel[2]),
		.A2(I2[15]),
		.B1(out_sel[3]),
		.B2(I3[15]),
		.Z(O1[15])
	);
	AO_CELL inst_2_15(
		.A1(out_sel[4]),
		.A2(I4[15]),
		.B1(out_sel[5]),
		.B2(I5[15]),
		.Z(O2[15])
	);
	AN_CELL inst_and_15(
		.A1(out_sel[6]),
		.A2(I6[15]),
		.Z(O3[15])
	);
	AO_CELL inst_0_16(
		.A1(out_sel[0]),
		.A2(I0[16]),
		.B1(out_sel[1]),
		.B2(I1[16]),
		.Z(O0[16])
	);
	AO_CELL inst_1_16(
		.A1(out_sel[2]),
		.A2(I2[16]),
		.B1(out_sel[3]),
		.B2(I3[16]),
		.Z(O1[16])
	);
	AO_CELL inst_2_16(
		.A1(out_sel[4]),
		.A2(I4[16]),
		.B1(out_sel[5]),
		.B2(I5[16]),
		.Z(O2[16])
	);
	AN_CELL inst_and_16(
		.A1(out_sel[6]),
		.A2(I6[16]),
		.Z(O3[16])
	);
	AO_CELL inst_0_valid(
		.A1(out_sel[0]),
		.A2(valid_in[0]),
		.B1(out_sel[1]),
		.B2(valid_in[1]),
		.Z(valid_out[0])
	);
	AO_CELL inst_1_valid(
		.A1(out_sel[2]),
		.A2(valid_in[2]),
		.B1(out_sel[3]),
		.B2(valid_in[3]),
		.Z(valid_out[1])
	);
	AO_CELL inst_2_valid(
		.A1(out_sel[4]),
		.A2(valid_in[4]),
		.B1(out_sel[5]),
		.B2(valid_in[5]),
		.Z(valid_out[2])
	);
	AN_CELL inst_and_3_valid(
		.A1(out_sel[6]),
		.A2(valid_in[6]),
		.Z(valid_out[3])
	);
endmodule
module mux_aoi_ready_valid_6_17 (
	I,
	S,
	ready_in,
	ready_out,
	valid_in,
	valid_out,
	out_sel,
	O
);
	input wire [101:0] I;
	input wire [2:0] S;
	input wire ready_in;
	output wire ready_out;
	input wire [5:0] valid_in;
	output wire valid_out;
	output wire [7:0] out_sel;
	output wire [16:0] O;
	wire [16:0] O_int0;
	wire [16:0] O_int1;
	wire [16:0] O_int2;
	wire [2:0] valid_out_temp;
	precoder_17_6 u_precoder(
		.S(S),
		.out_sel(out_sel)
	);
	mux_logic_17_6 u_mux_logic(
		.I0(I[0+:17]),
		.I1(I[17+:17]),
		.I2(I[34+:17]),
		.I3(I[51+:17]),
		.I4(I[68+:17]),
		.I5(I[85+:17]),
		.out_sel(out_sel),
		.valid_in(valid_in),
		.valid_out(valid_out_temp),
		.O0(O_int0),
		.O1(O_int1),
		.O2(O_int2)
	);
	assign O = (O_int0 | O_int1) | O_int2;
	assign ready_out = ready_in;
	assign valid_out = |valid_out_temp;
endmodule
module precoder_17_6 (
	S,
	out_sel
);
	input wire [2:0] S;
	output reg [7:0] out_sel;
	always @(*) begin : mux_sel
		case (S)
			3'd0: out_sel = 8'b00000001;
			3'd1: out_sel = 8'b00000010;
			3'd2: out_sel = 8'b00000100;
			3'd3: out_sel = 8'b00001000;
			3'd4: out_sel = 8'b00010000;
			3'd5: out_sel = 8'b00100000;
			default: out_sel = 8'b00000000;
		endcase
	end
endmodule
module mux_logic_17_6 (
	out_sel,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	valid_in,
	valid_out,
	O0,
	O1,
	O2
);
	input wire [7:0] out_sel;
	input wire [16:0] I0;
	input wire [16:0] I1;
	input wire [16:0] I2;
	input wire [16:0] I3;
	input wire [16:0] I4;
	input wire [16:0] I5;
	input wire [5:0] valid_in;
	output wire [2:0] valid_out;
	output wire [16:0] O0;
	output wire [16:0] O1;
	output wire [16:0] O2;
	AO_CELL inst_0_0(
		.A1(out_sel[0]),
		.A2(I0[0]),
		.B1(out_sel[1]),
		.B2(I1[0]),
		.Z(O0[0])
	);
	AO_CELL inst_1_0(
		.A1(out_sel[2]),
		.A2(I2[0]),
		.B1(out_sel[3]),
		.B2(I3[0]),
		.Z(O1[0])
	);
	AO_CELL inst_2_0(
		.A1(out_sel[4]),
		.A2(I4[0]),
		.B1(out_sel[5]),
		.B2(I5[0]),
		.Z(O2[0])
	);
	AO_CELL inst_0_1(
		.A1(out_sel[0]),
		.A2(I0[1]),
		.B1(out_sel[1]),
		.B2(I1[1]),
		.Z(O0[1])
	);
	AO_CELL inst_1_1(
		.A1(out_sel[2]),
		.A2(I2[1]),
		.B1(out_sel[3]),
		.B2(I3[1]),
		.Z(O1[1])
	);
	AO_CELL inst_2_1(
		.A1(out_sel[4]),
		.A2(I4[1]),
		.B1(out_sel[5]),
		.B2(I5[1]),
		.Z(O2[1])
	);
	AO_CELL inst_0_2(
		.A1(out_sel[0]),
		.A2(I0[2]),
		.B1(out_sel[1]),
		.B2(I1[2]),
		.Z(O0[2])
	);
	AO_CELL inst_1_2(
		.A1(out_sel[2]),
		.A2(I2[2]),
		.B1(out_sel[3]),
		.B2(I3[2]),
		.Z(O1[2])
	);
	AO_CELL inst_2_2(
		.A1(out_sel[4]),
		.A2(I4[2]),
		.B1(out_sel[5]),
		.B2(I5[2]),
		.Z(O2[2])
	);
	AO_CELL inst_0_3(
		.A1(out_sel[0]),
		.A2(I0[3]),
		.B1(out_sel[1]),
		.B2(I1[3]),
		.Z(O0[3])
	);
	AO_CELL inst_1_3(
		.A1(out_sel[2]),
		.A2(I2[3]),
		.B1(out_sel[3]),
		.B2(I3[3]),
		.Z(O1[3])
	);
	AO_CELL inst_2_3(
		.A1(out_sel[4]),
		.A2(I4[3]),
		.B1(out_sel[5]),
		.B2(I5[3]),
		.Z(O2[3])
	);
	AO_CELL inst_0_4(
		.A1(out_sel[0]),
		.A2(I0[4]),
		.B1(out_sel[1]),
		.B2(I1[4]),
		.Z(O0[4])
	);
	AO_CELL inst_1_4(
		.A1(out_sel[2]),
		.A2(I2[4]),
		.B1(out_sel[3]),
		.B2(I3[4]),
		.Z(O1[4])
	);
	AO_CELL inst_2_4(
		.A1(out_sel[4]),
		.A2(I4[4]),
		.B1(out_sel[5]),
		.B2(I5[4]),
		.Z(O2[4])
	);
	AO_CELL inst_0_5(
		.A1(out_sel[0]),
		.A2(I0[5]),
		.B1(out_sel[1]),
		.B2(I1[5]),
		.Z(O0[5])
	);
	AO_CELL inst_1_5(
		.A1(out_sel[2]),
		.A2(I2[5]),
		.B1(out_sel[3]),
		.B2(I3[5]),
		.Z(O1[5])
	);
	AO_CELL inst_2_5(
		.A1(out_sel[4]),
		.A2(I4[5]),
		.B1(out_sel[5]),
		.B2(I5[5]),
		.Z(O2[5])
	);
	AO_CELL inst_0_6(
		.A1(out_sel[0]),
		.A2(I0[6]),
		.B1(out_sel[1]),
		.B2(I1[6]),
		.Z(O0[6])
	);
	AO_CELL inst_1_6(
		.A1(out_sel[2]),
		.A2(I2[6]),
		.B1(out_sel[3]),
		.B2(I3[6]),
		.Z(O1[6])
	);
	AO_CELL inst_2_6(
		.A1(out_sel[4]),
		.A2(I4[6]),
		.B1(out_sel[5]),
		.B2(I5[6]),
		.Z(O2[6])
	);
	AO_CELL inst_0_7(
		.A1(out_sel[0]),
		.A2(I0[7]),
		.B1(out_sel[1]),
		.B2(I1[7]),
		.Z(O0[7])
	);
	AO_CELL inst_1_7(
		.A1(out_sel[2]),
		.A2(I2[7]),
		.B1(out_sel[3]),
		.B2(I3[7]),
		.Z(O1[7])
	);
	AO_CELL inst_2_7(
		.A1(out_sel[4]),
		.A2(I4[7]),
		.B1(out_sel[5]),
		.B2(I5[7]),
		.Z(O2[7])
	);
	AO_CELL inst_0_8(
		.A1(out_sel[0]),
		.A2(I0[8]),
		.B1(out_sel[1]),
		.B2(I1[8]),
		.Z(O0[8])
	);
	AO_CELL inst_1_8(
		.A1(out_sel[2]),
		.A2(I2[8]),
		.B1(out_sel[3]),
		.B2(I3[8]),
		.Z(O1[8])
	);
	AO_CELL inst_2_8(
		.A1(out_sel[4]),
		.A2(I4[8]),
		.B1(out_sel[5]),
		.B2(I5[8]),
		.Z(O2[8])
	);
	AO_CELL inst_0_9(
		.A1(out_sel[0]),
		.A2(I0[9]),
		.B1(out_sel[1]),
		.B2(I1[9]),
		.Z(O0[9])
	);
	AO_CELL inst_1_9(
		.A1(out_sel[2]),
		.A2(I2[9]),
		.B1(out_sel[3]),
		.B2(I3[9]),
		.Z(O1[9])
	);
	AO_CELL inst_2_9(
		.A1(out_sel[4]),
		.A2(I4[9]),
		.B1(out_sel[5]),
		.B2(I5[9]),
		.Z(O2[9])
	);
	AO_CELL inst_0_10(
		.A1(out_sel[0]),
		.A2(I0[10]),
		.B1(out_sel[1]),
		.B2(I1[10]),
		.Z(O0[10])
	);
	AO_CELL inst_1_10(
		.A1(out_sel[2]),
		.A2(I2[10]),
		.B1(out_sel[3]),
		.B2(I3[10]),
		.Z(O1[10])
	);
	AO_CELL inst_2_10(
		.A1(out_sel[4]),
		.A2(I4[10]),
		.B1(out_sel[5]),
		.B2(I5[10]),
		.Z(O2[10])
	);
	AO_CELL inst_0_11(
		.A1(out_sel[0]),
		.A2(I0[11]),
		.B1(out_sel[1]),
		.B2(I1[11]),
		.Z(O0[11])
	);
	AO_CELL inst_1_11(
		.A1(out_sel[2]),
		.A2(I2[11]),
		.B1(out_sel[3]),
		.B2(I3[11]),
		.Z(O1[11])
	);
	AO_CELL inst_2_11(
		.A1(out_sel[4]),
		.A2(I4[11]),
		.B1(out_sel[5]),
		.B2(I5[11]),
		.Z(O2[11])
	);
	AO_CELL inst_0_12(
		.A1(out_sel[0]),
		.A2(I0[12]),
		.B1(out_sel[1]),
		.B2(I1[12]),
		.Z(O0[12])
	);
	AO_CELL inst_1_12(
		.A1(out_sel[2]),
		.A2(I2[12]),
		.B1(out_sel[3]),
		.B2(I3[12]),
		.Z(O1[12])
	);
	AO_CELL inst_2_12(
		.A1(out_sel[4]),
		.A2(I4[12]),
		.B1(out_sel[5]),
		.B2(I5[12]),
		.Z(O2[12])
	);
	AO_CELL inst_0_13(
		.A1(out_sel[0]),
		.A2(I0[13]),
		.B1(out_sel[1]),
		.B2(I1[13]),
		.Z(O0[13])
	);
	AO_CELL inst_1_13(
		.A1(out_sel[2]),
		.A2(I2[13]),
		.B1(out_sel[3]),
		.B2(I3[13]),
		.Z(O1[13])
	);
	AO_CELL inst_2_13(
		.A1(out_sel[4]),
		.A2(I4[13]),
		.B1(out_sel[5]),
		.B2(I5[13]),
		.Z(O2[13])
	);
	AO_CELL inst_0_14(
		.A1(out_sel[0]),
		.A2(I0[14]),
		.B1(out_sel[1]),
		.B2(I1[14]),
		.Z(O0[14])
	);
	AO_CELL inst_1_14(
		.A1(out_sel[2]),
		.A2(I2[14]),
		.B1(out_sel[3]),
		.B2(I3[14]),
		.Z(O1[14])
	);
	AO_CELL inst_2_14(
		.A1(out_sel[4]),
		.A2(I4[14]),
		.B1(out_sel[5]),
		.B2(I5[14]),
		.Z(O2[14])
	);
	AO_CELL inst_0_15(
		.A1(out_sel[0]),
		.A2(I0[15]),
		.B1(out_sel[1]),
		.B2(I1[15]),
		.Z(O0[15])
	);
	AO_CELL inst_1_15(
		.A1(out_sel[2]),
		.A2(I2[15]),
		.B1(out_sel[3]),
		.B2(I3[15]),
		.Z(O1[15])
	);
	AO_CELL inst_2_15(
		.A1(out_sel[4]),
		.A2(I4[15]),
		.B1(out_sel[5]),
		.B2(I5[15]),
		.Z(O2[15])
	);
	AO_CELL inst_0_16(
		.A1(out_sel[0]),
		.A2(I0[16]),
		.B1(out_sel[1]),
		.B2(I1[16]),
		.Z(O0[16])
	);
	AO_CELL inst_1_16(
		.A1(out_sel[2]),
		.A2(I2[16]),
		.B1(out_sel[3]),
		.B2(I3[16]),
		.Z(O1[16])
	);
	AO_CELL inst_2_16(
		.A1(out_sel[4]),
		.A2(I4[16]),
		.B1(out_sel[5]),
		.B2(I5[16]),
		.Z(O2[16])
	);
	AO_CELL inst_0_valid(
		.A1(out_sel[0]),
		.A2(valid_in[0]),
		.B1(out_sel[1]),
		.B2(valid_in[1]),
		.Z(valid_out[0])
	);
	AO_CELL inst_1_valid(
		.A1(out_sel[2]),
		.A2(valid_in[2]),
		.B1(out_sel[3]),
		.B2(valid_in[3]),
		.Z(valid_out[1])
	);
	AO_CELL inst_2_valid(
		.A1(out_sel[4]),
		.A2(valid_in[4]),
		.B1(out_sel[5]),
		.B2(valid_in[5]),
		.Z(valid_out[2])
	);
endmodule
module mux_aoi_ready_valid_6_1 (
	I,
	S,
	ready_in,
	ready_out,
	valid_in,
	valid_out,
	out_sel,
	O
);
	input wire [5:0] I;
	input wire [2:0] S;
	input wire ready_in;
	output wire ready_out;
	input wire [5:0] valid_in;
	output wire valid_out;
	output wire [7:0] out_sel;
	output wire [0:0] O;
	wire [0:0] O_int0;
	wire [0:0] O_int1;
	wire [0:0] O_int2;
	wire [2:0] valid_out_temp;
	precoder_1_6 u_precoder(
		.S(S),
		.out_sel(out_sel)
	);
	mux_logic_1_6 u_mux_logic(
		.I0(I[0+:1]),
		.I1(I[1+:1]),
		.I2(I[2+:1]),
		.I3(I[3+:1]),
		.I4(I[4+:1]),
		.I5(I[5+:1]),
		.out_sel(out_sel),
		.valid_in(valid_in),
		.valid_out(valid_out_temp),
		.O0(O_int0),
		.O1(O_int1),
		.O2(O_int2)
	);
	assign O = (O_int0 | O_int1) | O_int2;
	assign ready_out = ready_in;
	assign valid_out = |valid_out_temp;
endmodule
module precoder_1_6 (
	S,
	out_sel
);
	input wire [2:0] S;
	output reg [7:0] out_sel;
	always @(*) begin : mux_sel
		case (S)
			3'd0: out_sel = 8'b00000001;
			3'd1: out_sel = 8'b00000010;
			3'd2: out_sel = 8'b00000100;
			3'd3: out_sel = 8'b00001000;
			3'd4: out_sel = 8'b00010000;
			3'd5: out_sel = 8'b00100000;
			default: out_sel = 8'b00000000;
		endcase
	end
endmodule
module mux_logic_1_6 (
	out_sel,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	valid_in,
	valid_out,
	O0,
	O1,
	O2
);
	input wire [7:0] out_sel;
	input wire [0:0] I0;
	input wire [0:0] I1;
	input wire [0:0] I2;
	input wire [0:0] I3;
	input wire [0:0] I4;
	input wire [0:0] I5;
	input wire [5:0] valid_in;
	output wire [2:0] valid_out;
	output wire [0:0] O0;
	output wire [0:0] O1;
	output wire [0:0] O2;
	AO_CELL inst_0_0(
		.A1(out_sel[0]),
		.A2(I0[0]),
		.B1(out_sel[1]),
		.B2(I1[0]),
		.Z(O0[0])
	);
	AO_CELL inst_1_0(
		.A1(out_sel[2]),
		.A2(I2[0]),
		.B1(out_sel[3]),
		.B2(I3[0]),
		.Z(O1[0])
	);
	AO_CELL inst_2_0(
		.A1(out_sel[4]),
		.A2(I4[0]),
		.B1(out_sel[5]),
		.B2(I5[0]),
		.Z(O2[0])
	);
	AO_CELL inst_0_valid(
		.A1(out_sel[0]),
		.A2(valid_in[0]),
		.B1(out_sel[1]),
		.B2(valid_in[1]),
		.Z(valid_out[0])
	);
	AO_CELL inst_1_valid(
		.A1(out_sel[2]),
		.A2(valid_in[2]),
		.B1(out_sel[3]),
		.B2(valid_in[3]),
		.Z(valid_out[1])
	);
	AO_CELL inst_2_valid(
		.A1(out_sel[4]),
		.A2(valid_in[4]),
		.B1(out_sel[5]),
		.B2(valid_in[5]),
		.Z(valid_out[2])
	);
endmodule
module mux_aoi_ready_valid_2_17 (
	I,
	S,
	ready_in,
	ready_out,
	valid_in,
	valid_out,
	out_sel,
	O
);
	input wire [33:0] I;
	input wire S;
	input wire ready_in;
	output wire ready_out;
	input wire [1:0] valid_in;
	output wire valid_out;
	output wire [1:0] out_sel;
	output wire [16:0] O;
	wire [16:0] O_int0;
	wire [0:0] valid_out_temp;
	precoder_17_2 u_precoder(
		.S(S),
		.out_sel(out_sel)
	);
	mux_logic_17_2 u_mux_logic(
		.I0(I[0+:17]),
		.I1(I[17+:17]),
		.out_sel(out_sel),
		.valid_in(valid_in),
		.valid_out(valid_out_temp),
		.O0(O_int0)
	);
	assign O = O_int0;
	assign ready_out = ready_in;
	assign valid_out = |valid_out_temp;
endmodule
module precoder_17_2 (
	S,
	out_sel
);
	input wire [0:0] S;
	output reg [1:0] out_sel;
	always @(*) begin : mux_sel
		case (S)
			1'd0: out_sel = 2'b01;
			1'd1: out_sel = 2'b10;
			default: out_sel = 2'b00;
		endcase
	end
endmodule
module mux_logic_17_2 (
	out_sel,
	I0,
	I1,
	valid_in,
	valid_out,
	O0
);
	input wire [1:0] out_sel;
	input wire [16:0] I0;
	input wire [16:0] I1;
	input wire [1:0] valid_in;
	output wire [0:0] valid_out;
	output wire [16:0] O0;
	AO_CELL inst_0_0(
		.A1(out_sel[0]),
		.A2(I0[0]),
		.B1(out_sel[1]),
		.B2(I1[0]),
		.Z(O0[0])
	);
	AO_CELL inst_0_1(
		.A1(out_sel[0]),
		.A2(I0[1]),
		.B1(out_sel[1]),
		.B2(I1[1]),
		.Z(O0[1])
	);
	AO_CELL inst_0_2(
		.A1(out_sel[0]),
		.A2(I0[2]),
		.B1(out_sel[1]),
		.B2(I1[2]),
		.Z(O0[2])
	);
	AO_CELL inst_0_3(
		.A1(out_sel[0]),
		.A2(I0[3]),
		.B1(out_sel[1]),
		.B2(I1[3]),
		.Z(O0[3])
	);
	AO_CELL inst_0_4(
		.A1(out_sel[0]),
		.A2(I0[4]),
		.B1(out_sel[1]),
		.B2(I1[4]),
		.Z(O0[4])
	);
	AO_CELL inst_0_5(
		.A1(out_sel[0]),
		.A2(I0[5]),
		.B1(out_sel[1]),
		.B2(I1[5]),
		.Z(O0[5])
	);
	AO_CELL inst_0_6(
		.A1(out_sel[0]),
		.A2(I0[6]),
		.B1(out_sel[1]),
		.B2(I1[6]),
		.Z(O0[6])
	);
	AO_CELL inst_0_7(
		.A1(out_sel[0]),
		.A2(I0[7]),
		.B1(out_sel[1]),
		.B2(I1[7]),
		.Z(O0[7])
	);
	AO_CELL inst_0_8(
		.A1(out_sel[0]),
		.A2(I0[8]),
		.B1(out_sel[1]),
		.B2(I1[8]),
		.Z(O0[8])
	);
	AO_CELL inst_0_9(
		.A1(out_sel[0]),
		.A2(I0[9]),
		.B1(out_sel[1]),
		.B2(I1[9]),
		.Z(O0[9])
	);
	AO_CELL inst_0_10(
		.A1(out_sel[0]),
		.A2(I0[10]),
		.B1(out_sel[1]),
		.B2(I1[10]),
		.Z(O0[10])
	);
	AO_CELL inst_0_11(
		.A1(out_sel[0]),
		.A2(I0[11]),
		.B1(out_sel[1]),
		.B2(I1[11]),
		.Z(O0[11])
	);
	AO_CELL inst_0_12(
		.A1(out_sel[0]),
		.A2(I0[12]),
		.B1(out_sel[1]),
		.B2(I1[12]),
		.Z(O0[12])
	);
	AO_CELL inst_0_13(
		.A1(out_sel[0]),
		.A2(I0[13]),
		.B1(out_sel[1]),
		.B2(I1[13]),
		.Z(O0[13])
	);
	AO_CELL inst_0_14(
		.A1(out_sel[0]),
		.A2(I0[14]),
		.B1(out_sel[1]),
		.B2(I1[14]),
		.Z(O0[14])
	);
	AO_CELL inst_0_15(
		.A1(out_sel[0]),
		.A2(I0[15]),
		.B1(out_sel[1]),
		.B2(I1[15]),
		.Z(O0[15])
	);
	AO_CELL inst_0_16(
		.A1(out_sel[0]),
		.A2(I0[16]),
		.B1(out_sel[1]),
		.B2(I1[16]),
		.Z(O0[16])
	);
	AO_CELL inst_0_valid(
		.A1(out_sel[0]),
		.A2(valid_in[0]),
		.B1(out_sel[1]),
		.B2(valid_in[1]),
		.Z(valid_out[0])
	);
endmodule
module mux_aoi_ready_valid_2_1 (
	I,
	S,
	ready_in,
	ready_out,
	valid_in,
	valid_out,
	out_sel,
	O
);
	input wire [1:0] I;
	input wire S;
	input wire ready_in;
	output wire ready_out;
	input wire [1:0] valid_in;
	output wire valid_out;
	output wire [1:0] out_sel;
	output wire [0:0] O;
	wire [0:0] O_int0;
	wire [0:0] valid_out_temp;
	precoder_1_2 u_precoder(
		.S(S),
		.out_sel(out_sel)
	);
	mux_logic_1_2 u_mux_logic(
		.I0(I[0+:1]),
		.I1(I[1+:1]),
		.out_sel(out_sel),
		.valid_in(valid_in),
		.valid_out(valid_out_temp),
		.O0(O_int0)
	);
	assign O = O_int0;
	assign ready_out = ready_in;
	assign valid_out = |valid_out_temp;
endmodule
module precoder_1_2 (
	S,
	out_sel
);
	input wire [0:0] S;
	output reg [1:0] out_sel;
	always @(*) begin : mux_sel
		case (S)
			1'd0: out_sel = 2'b01;
			1'd1: out_sel = 2'b10;
			default: out_sel = 2'b00;
		endcase
	end
endmodule
module mux_logic_1_2 (
	out_sel,
	I0,
	I1,
	valid_in,
	valid_out,
	O0
);
	input wire [1:0] out_sel;
	input wire [0:0] I0;
	input wire [0:0] I1;
	input wire [1:0] valid_in;
	output wire [0:0] valid_out;
	output wire [0:0] O0;
	AO_CELL inst_0_0(
		.A1(out_sel[0]),
		.A2(I0[0]),
		.B1(out_sel[1]),
		.B2(I1[0]),
		.Z(O0[0])
	);
	AO_CELL inst_0_valid(
		.A1(out_sel[0]),
		.A2(valid_in[0]),
		.B1(out_sel[1]),
		.B2(valid_in[1]),
		.Z(valid_out[0])
	);
endmodule
module mux_aoi_7_32 (
	I,
	S,
	out_sel,
	O
);
	input wire [223:0] I;
	input wire [2:0] S;
	output wire [7:0] out_sel;
	output wire [31:0] O;
	wire [31:0] O_int0;
	wire [31:0] O_int1;
	wire [31:0] O_int2;
	wire [31:0] O_int3;
	precoder_32_7 u_precoder(
		.S(S),
		.out_sel(out_sel)
	);
	mux_logic_32_7 u_mux_logic(
		.I0(I[0+:32]),
		.I1(I[32+:32]),
		.I2(I[64+:32]),
		.I3(I[96+:32]),
		.I4(I[128+:32]),
		.I5(I[160+:32]),
		.I6(I[192+:32]),
		.out_sel(out_sel),
		.O0(O_int0),
		.O1(O_int1),
		.O2(O_int2),
		.O3(O_int3)
	);
	assign O = ((O_int0 | O_int1) | O_int2) | O_int3;
endmodule
module precoder_32_7 (
	S,
	out_sel
);
	input wire [2:0] S;
	output reg [7:0] out_sel;
	always @(*) begin : mux_sel
		case (S)
			3'd0: out_sel = 8'b00000001;
			3'd1: out_sel = 8'b00000010;
			3'd2: out_sel = 8'b00000100;
			3'd3: out_sel = 8'b00001000;
			3'd4: out_sel = 8'b00010000;
			3'd5: out_sel = 8'b00100000;
			3'd6: out_sel = 8'b01000000;
			default: out_sel = 8'b00000000;
		endcase
	end
endmodule
module mux_logic_32_7 (
	out_sel,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	O0,
	O1,
	O2,
	O3
);
	input wire [7:0] out_sel;
	input wire [31:0] I0;
	input wire [31:0] I1;
	input wire [31:0] I2;
	input wire [31:0] I3;
	input wire [31:0] I4;
	input wire [31:0] I5;
	input wire [31:0] I6;
	output wire [31:0] O0;
	output wire [31:0] O1;
	output wire [31:0] O2;
	output wire [31:0] O3;
	AO_CELL inst_0_0(
		.A1(out_sel[0]),
		.A2(I0[0]),
		.B1(out_sel[1]),
		.B2(I1[0]),
		.Z(O0[0])
	);
	AO_CELL inst_1_0(
		.A1(out_sel[2]),
		.A2(I2[0]),
		.B1(out_sel[3]),
		.B2(I3[0]),
		.Z(O1[0])
	);
	AO_CELL inst_2_0(
		.A1(out_sel[4]),
		.A2(I4[0]),
		.B1(out_sel[5]),
		.B2(I5[0]),
		.Z(O2[0])
	);
	AN_CELL inst_and_0(
		.A1(out_sel[6]),
		.A2(I6[0]),
		.Z(O3[0])
	);
	AO_CELL inst_0_1(
		.A1(out_sel[0]),
		.A2(I0[1]),
		.B1(out_sel[1]),
		.B2(I1[1]),
		.Z(O0[1])
	);
	AO_CELL inst_1_1(
		.A1(out_sel[2]),
		.A2(I2[1]),
		.B1(out_sel[3]),
		.B2(I3[1]),
		.Z(O1[1])
	);
	AO_CELL inst_2_1(
		.A1(out_sel[4]),
		.A2(I4[1]),
		.B1(out_sel[5]),
		.B2(I5[1]),
		.Z(O2[1])
	);
	AN_CELL inst_and_1(
		.A1(out_sel[6]),
		.A2(I6[1]),
		.Z(O3[1])
	);
	AO_CELL inst_0_2(
		.A1(out_sel[0]),
		.A2(I0[2]),
		.B1(out_sel[1]),
		.B2(I1[2]),
		.Z(O0[2])
	);
	AO_CELL inst_1_2(
		.A1(out_sel[2]),
		.A2(I2[2]),
		.B1(out_sel[3]),
		.B2(I3[2]),
		.Z(O1[2])
	);
	AO_CELL inst_2_2(
		.A1(out_sel[4]),
		.A2(I4[2]),
		.B1(out_sel[5]),
		.B2(I5[2]),
		.Z(O2[2])
	);
	AN_CELL inst_and_2(
		.A1(out_sel[6]),
		.A2(I6[2]),
		.Z(O3[2])
	);
	AO_CELL inst_0_3(
		.A1(out_sel[0]),
		.A2(I0[3]),
		.B1(out_sel[1]),
		.B2(I1[3]),
		.Z(O0[3])
	);
	AO_CELL inst_1_3(
		.A1(out_sel[2]),
		.A2(I2[3]),
		.B1(out_sel[3]),
		.B2(I3[3]),
		.Z(O1[3])
	);
	AO_CELL inst_2_3(
		.A1(out_sel[4]),
		.A2(I4[3]),
		.B1(out_sel[5]),
		.B2(I5[3]),
		.Z(O2[3])
	);
	AN_CELL inst_and_3(
		.A1(out_sel[6]),
		.A2(I6[3]),
		.Z(O3[3])
	);
	AO_CELL inst_0_4(
		.A1(out_sel[0]),
		.A2(I0[4]),
		.B1(out_sel[1]),
		.B2(I1[4]),
		.Z(O0[4])
	);
	AO_CELL inst_1_4(
		.A1(out_sel[2]),
		.A2(I2[4]),
		.B1(out_sel[3]),
		.B2(I3[4]),
		.Z(O1[4])
	);
	AO_CELL inst_2_4(
		.A1(out_sel[4]),
		.A2(I4[4]),
		.B1(out_sel[5]),
		.B2(I5[4]),
		.Z(O2[4])
	);
	AN_CELL inst_and_4(
		.A1(out_sel[6]),
		.A2(I6[4]),
		.Z(O3[4])
	);
	AO_CELL inst_0_5(
		.A1(out_sel[0]),
		.A2(I0[5]),
		.B1(out_sel[1]),
		.B2(I1[5]),
		.Z(O0[5])
	);
	AO_CELL inst_1_5(
		.A1(out_sel[2]),
		.A2(I2[5]),
		.B1(out_sel[3]),
		.B2(I3[5]),
		.Z(O1[5])
	);
	AO_CELL inst_2_5(
		.A1(out_sel[4]),
		.A2(I4[5]),
		.B1(out_sel[5]),
		.B2(I5[5]),
		.Z(O2[5])
	);
	AN_CELL inst_and_5(
		.A1(out_sel[6]),
		.A2(I6[5]),
		.Z(O3[5])
	);
	AO_CELL inst_0_6(
		.A1(out_sel[0]),
		.A2(I0[6]),
		.B1(out_sel[1]),
		.B2(I1[6]),
		.Z(O0[6])
	);
	AO_CELL inst_1_6(
		.A1(out_sel[2]),
		.A2(I2[6]),
		.B1(out_sel[3]),
		.B2(I3[6]),
		.Z(O1[6])
	);
	AO_CELL inst_2_6(
		.A1(out_sel[4]),
		.A2(I4[6]),
		.B1(out_sel[5]),
		.B2(I5[6]),
		.Z(O2[6])
	);
	AN_CELL inst_and_6(
		.A1(out_sel[6]),
		.A2(I6[6]),
		.Z(O3[6])
	);
	AO_CELL inst_0_7(
		.A1(out_sel[0]),
		.A2(I0[7]),
		.B1(out_sel[1]),
		.B2(I1[7]),
		.Z(O0[7])
	);
	AO_CELL inst_1_7(
		.A1(out_sel[2]),
		.A2(I2[7]),
		.B1(out_sel[3]),
		.B2(I3[7]),
		.Z(O1[7])
	);
	AO_CELL inst_2_7(
		.A1(out_sel[4]),
		.A2(I4[7]),
		.B1(out_sel[5]),
		.B2(I5[7]),
		.Z(O2[7])
	);
	AN_CELL inst_and_7(
		.A1(out_sel[6]),
		.A2(I6[7]),
		.Z(O3[7])
	);
	AO_CELL inst_0_8(
		.A1(out_sel[0]),
		.A2(I0[8]),
		.B1(out_sel[1]),
		.B2(I1[8]),
		.Z(O0[8])
	);
	AO_CELL inst_1_8(
		.A1(out_sel[2]),
		.A2(I2[8]),
		.B1(out_sel[3]),
		.B2(I3[8]),
		.Z(O1[8])
	);
	AO_CELL inst_2_8(
		.A1(out_sel[4]),
		.A2(I4[8]),
		.B1(out_sel[5]),
		.B2(I5[8]),
		.Z(O2[8])
	);
	AN_CELL inst_and_8(
		.A1(out_sel[6]),
		.A2(I6[8]),
		.Z(O3[8])
	);
	AO_CELL inst_0_9(
		.A1(out_sel[0]),
		.A2(I0[9]),
		.B1(out_sel[1]),
		.B2(I1[9]),
		.Z(O0[9])
	);
	AO_CELL inst_1_9(
		.A1(out_sel[2]),
		.A2(I2[9]),
		.B1(out_sel[3]),
		.B2(I3[9]),
		.Z(O1[9])
	);
	AO_CELL inst_2_9(
		.A1(out_sel[4]),
		.A2(I4[9]),
		.B1(out_sel[5]),
		.B2(I5[9]),
		.Z(O2[9])
	);
	AN_CELL inst_and_9(
		.A1(out_sel[6]),
		.A2(I6[9]),
		.Z(O3[9])
	);
	AO_CELL inst_0_10(
		.A1(out_sel[0]),
		.A2(I0[10]),
		.B1(out_sel[1]),
		.B2(I1[10]),
		.Z(O0[10])
	);
	AO_CELL inst_1_10(
		.A1(out_sel[2]),
		.A2(I2[10]),
		.B1(out_sel[3]),
		.B2(I3[10]),
		.Z(O1[10])
	);
	AO_CELL inst_2_10(
		.A1(out_sel[4]),
		.A2(I4[10]),
		.B1(out_sel[5]),
		.B2(I5[10]),
		.Z(O2[10])
	);
	AN_CELL inst_and_10(
		.A1(out_sel[6]),
		.A2(I6[10]),
		.Z(O3[10])
	);
	AO_CELL inst_0_11(
		.A1(out_sel[0]),
		.A2(I0[11]),
		.B1(out_sel[1]),
		.B2(I1[11]),
		.Z(O0[11])
	);
	AO_CELL inst_1_11(
		.A1(out_sel[2]),
		.A2(I2[11]),
		.B1(out_sel[3]),
		.B2(I3[11]),
		.Z(O1[11])
	);
	AO_CELL inst_2_11(
		.A1(out_sel[4]),
		.A2(I4[11]),
		.B1(out_sel[5]),
		.B2(I5[11]),
		.Z(O2[11])
	);
	AN_CELL inst_and_11(
		.A1(out_sel[6]),
		.A2(I6[11]),
		.Z(O3[11])
	);
	AO_CELL inst_0_12(
		.A1(out_sel[0]),
		.A2(I0[12]),
		.B1(out_sel[1]),
		.B2(I1[12]),
		.Z(O0[12])
	);
	AO_CELL inst_1_12(
		.A1(out_sel[2]),
		.A2(I2[12]),
		.B1(out_sel[3]),
		.B2(I3[12]),
		.Z(O1[12])
	);
	AO_CELL inst_2_12(
		.A1(out_sel[4]),
		.A2(I4[12]),
		.B1(out_sel[5]),
		.B2(I5[12]),
		.Z(O2[12])
	);
	AN_CELL inst_and_12(
		.A1(out_sel[6]),
		.A2(I6[12]),
		.Z(O3[12])
	);
	AO_CELL inst_0_13(
		.A1(out_sel[0]),
		.A2(I0[13]),
		.B1(out_sel[1]),
		.B2(I1[13]),
		.Z(O0[13])
	);
	AO_CELL inst_1_13(
		.A1(out_sel[2]),
		.A2(I2[13]),
		.B1(out_sel[3]),
		.B2(I3[13]),
		.Z(O1[13])
	);
	AO_CELL inst_2_13(
		.A1(out_sel[4]),
		.A2(I4[13]),
		.B1(out_sel[5]),
		.B2(I5[13]),
		.Z(O2[13])
	);
	AN_CELL inst_and_13(
		.A1(out_sel[6]),
		.A2(I6[13]),
		.Z(O3[13])
	);
	AO_CELL inst_0_14(
		.A1(out_sel[0]),
		.A2(I0[14]),
		.B1(out_sel[1]),
		.B2(I1[14]),
		.Z(O0[14])
	);
	AO_CELL inst_1_14(
		.A1(out_sel[2]),
		.A2(I2[14]),
		.B1(out_sel[3]),
		.B2(I3[14]),
		.Z(O1[14])
	);
	AO_CELL inst_2_14(
		.A1(out_sel[4]),
		.A2(I4[14]),
		.B1(out_sel[5]),
		.B2(I5[14]),
		.Z(O2[14])
	);
	AN_CELL inst_and_14(
		.A1(out_sel[6]),
		.A2(I6[14]),
		.Z(O3[14])
	);
	AO_CELL inst_0_15(
		.A1(out_sel[0]),
		.A2(I0[15]),
		.B1(out_sel[1]),
		.B2(I1[15]),
		.Z(O0[15])
	);
	AO_CELL inst_1_15(
		.A1(out_sel[2]),
		.A2(I2[15]),
		.B1(out_sel[3]),
		.B2(I3[15]),
		.Z(O1[15])
	);
	AO_CELL inst_2_15(
		.A1(out_sel[4]),
		.A2(I4[15]),
		.B1(out_sel[5]),
		.B2(I5[15]),
		.Z(O2[15])
	);
	AN_CELL inst_and_15(
		.A1(out_sel[6]),
		.A2(I6[15]),
		.Z(O3[15])
	);
	AO_CELL inst_0_16(
		.A1(out_sel[0]),
		.A2(I0[16]),
		.B1(out_sel[1]),
		.B2(I1[16]),
		.Z(O0[16])
	);
	AO_CELL inst_1_16(
		.A1(out_sel[2]),
		.A2(I2[16]),
		.B1(out_sel[3]),
		.B2(I3[16]),
		.Z(O1[16])
	);
	AO_CELL inst_2_16(
		.A1(out_sel[4]),
		.A2(I4[16]),
		.B1(out_sel[5]),
		.B2(I5[16]),
		.Z(O2[16])
	);
	AN_CELL inst_and_16(
		.A1(out_sel[6]),
		.A2(I6[16]),
		.Z(O3[16])
	);
	AO_CELL inst_0_17(
		.A1(out_sel[0]),
		.A2(I0[17]),
		.B1(out_sel[1]),
		.B2(I1[17]),
		.Z(O0[17])
	);
	AO_CELL inst_1_17(
		.A1(out_sel[2]),
		.A2(I2[17]),
		.B1(out_sel[3]),
		.B2(I3[17]),
		.Z(O1[17])
	);
	AO_CELL inst_2_17(
		.A1(out_sel[4]),
		.A2(I4[17]),
		.B1(out_sel[5]),
		.B2(I5[17]),
		.Z(O2[17])
	);
	AN_CELL inst_and_17(
		.A1(out_sel[6]),
		.A2(I6[17]),
		.Z(O3[17])
	);
	AO_CELL inst_0_18(
		.A1(out_sel[0]),
		.A2(I0[18]),
		.B1(out_sel[1]),
		.B2(I1[18]),
		.Z(O0[18])
	);
	AO_CELL inst_1_18(
		.A1(out_sel[2]),
		.A2(I2[18]),
		.B1(out_sel[3]),
		.B2(I3[18]),
		.Z(O1[18])
	);
	AO_CELL inst_2_18(
		.A1(out_sel[4]),
		.A2(I4[18]),
		.B1(out_sel[5]),
		.B2(I5[18]),
		.Z(O2[18])
	);
	AN_CELL inst_and_18(
		.A1(out_sel[6]),
		.A2(I6[18]),
		.Z(O3[18])
	);
	AO_CELL inst_0_19(
		.A1(out_sel[0]),
		.A2(I0[19]),
		.B1(out_sel[1]),
		.B2(I1[19]),
		.Z(O0[19])
	);
	AO_CELL inst_1_19(
		.A1(out_sel[2]),
		.A2(I2[19]),
		.B1(out_sel[3]),
		.B2(I3[19]),
		.Z(O1[19])
	);
	AO_CELL inst_2_19(
		.A1(out_sel[4]),
		.A2(I4[19]),
		.B1(out_sel[5]),
		.B2(I5[19]),
		.Z(O2[19])
	);
	AN_CELL inst_and_19(
		.A1(out_sel[6]),
		.A2(I6[19]),
		.Z(O3[19])
	);
	AO_CELL inst_0_20(
		.A1(out_sel[0]),
		.A2(I0[20]),
		.B1(out_sel[1]),
		.B2(I1[20]),
		.Z(O0[20])
	);
	AO_CELL inst_1_20(
		.A1(out_sel[2]),
		.A2(I2[20]),
		.B1(out_sel[3]),
		.B2(I3[20]),
		.Z(O1[20])
	);
	AO_CELL inst_2_20(
		.A1(out_sel[4]),
		.A2(I4[20]),
		.B1(out_sel[5]),
		.B2(I5[20]),
		.Z(O2[20])
	);
	AN_CELL inst_and_20(
		.A1(out_sel[6]),
		.A2(I6[20]),
		.Z(O3[20])
	);
	AO_CELL inst_0_21(
		.A1(out_sel[0]),
		.A2(I0[21]),
		.B1(out_sel[1]),
		.B2(I1[21]),
		.Z(O0[21])
	);
	AO_CELL inst_1_21(
		.A1(out_sel[2]),
		.A2(I2[21]),
		.B1(out_sel[3]),
		.B2(I3[21]),
		.Z(O1[21])
	);
	AO_CELL inst_2_21(
		.A1(out_sel[4]),
		.A2(I4[21]),
		.B1(out_sel[5]),
		.B2(I5[21]),
		.Z(O2[21])
	);
	AN_CELL inst_and_21(
		.A1(out_sel[6]),
		.A2(I6[21]),
		.Z(O3[21])
	);
	AO_CELL inst_0_22(
		.A1(out_sel[0]),
		.A2(I0[22]),
		.B1(out_sel[1]),
		.B2(I1[22]),
		.Z(O0[22])
	);
	AO_CELL inst_1_22(
		.A1(out_sel[2]),
		.A2(I2[22]),
		.B1(out_sel[3]),
		.B2(I3[22]),
		.Z(O1[22])
	);
	AO_CELL inst_2_22(
		.A1(out_sel[4]),
		.A2(I4[22]),
		.B1(out_sel[5]),
		.B2(I5[22]),
		.Z(O2[22])
	);
	AN_CELL inst_and_22(
		.A1(out_sel[6]),
		.A2(I6[22]),
		.Z(O3[22])
	);
	AO_CELL inst_0_23(
		.A1(out_sel[0]),
		.A2(I0[23]),
		.B1(out_sel[1]),
		.B2(I1[23]),
		.Z(O0[23])
	);
	AO_CELL inst_1_23(
		.A1(out_sel[2]),
		.A2(I2[23]),
		.B1(out_sel[3]),
		.B2(I3[23]),
		.Z(O1[23])
	);
	AO_CELL inst_2_23(
		.A1(out_sel[4]),
		.A2(I4[23]),
		.B1(out_sel[5]),
		.B2(I5[23]),
		.Z(O2[23])
	);
	AN_CELL inst_and_23(
		.A1(out_sel[6]),
		.A2(I6[23]),
		.Z(O3[23])
	);
	AO_CELL inst_0_24(
		.A1(out_sel[0]),
		.A2(I0[24]),
		.B1(out_sel[1]),
		.B2(I1[24]),
		.Z(O0[24])
	);
	AO_CELL inst_1_24(
		.A1(out_sel[2]),
		.A2(I2[24]),
		.B1(out_sel[3]),
		.B2(I3[24]),
		.Z(O1[24])
	);
	AO_CELL inst_2_24(
		.A1(out_sel[4]),
		.A2(I4[24]),
		.B1(out_sel[5]),
		.B2(I5[24]),
		.Z(O2[24])
	);
	AN_CELL inst_and_24(
		.A1(out_sel[6]),
		.A2(I6[24]),
		.Z(O3[24])
	);
	AO_CELL inst_0_25(
		.A1(out_sel[0]),
		.A2(I0[25]),
		.B1(out_sel[1]),
		.B2(I1[25]),
		.Z(O0[25])
	);
	AO_CELL inst_1_25(
		.A1(out_sel[2]),
		.A2(I2[25]),
		.B1(out_sel[3]),
		.B2(I3[25]),
		.Z(O1[25])
	);
	AO_CELL inst_2_25(
		.A1(out_sel[4]),
		.A2(I4[25]),
		.B1(out_sel[5]),
		.B2(I5[25]),
		.Z(O2[25])
	);
	AN_CELL inst_and_25(
		.A1(out_sel[6]),
		.A2(I6[25]),
		.Z(O3[25])
	);
	AO_CELL inst_0_26(
		.A1(out_sel[0]),
		.A2(I0[26]),
		.B1(out_sel[1]),
		.B2(I1[26]),
		.Z(O0[26])
	);
	AO_CELL inst_1_26(
		.A1(out_sel[2]),
		.A2(I2[26]),
		.B1(out_sel[3]),
		.B2(I3[26]),
		.Z(O1[26])
	);
	AO_CELL inst_2_26(
		.A1(out_sel[4]),
		.A2(I4[26]),
		.B1(out_sel[5]),
		.B2(I5[26]),
		.Z(O2[26])
	);
	AN_CELL inst_and_26(
		.A1(out_sel[6]),
		.A2(I6[26]),
		.Z(O3[26])
	);
	AO_CELL inst_0_27(
		.A1(out_sel[0]),
		.A2(I0[27]),
		.B1(out_sel[1]),
		.B2(I1[27]),
		.Z(O0[27])
	);
	AO_CELL inst_1_27(
		.A1(out_sel[2]),
		.A2(I2[27]),
		.B1(out_sel[3]),
		.B2(I3[27]),
		.Z(O1[27])
	);
	AO_CELL inst_2_27(
		.A1(out_sel[4]),
		.A2(I4[27]),
		.B1(out_sel[5]),
		.B2(I5[27]),
		.Z(O2[27])
	);
	AN_CELL inst_and_27(
		.A1(out_sel[6]),
		.A2(I6[27]),
		.Z(O3[27])
	);
	AO_CELL inst_0_28(
		.A1(out_sel[0]),
		.A2(I0[28]),
		.B1(out_sel[1]),
		.B2(I1[28]),
		.Z(O0[28])
	);
	AO_CELL inst_1_28(
		.A1(out_sel[2]),
		.A2(I2[28]),
		.B1(out_sel[3]),
		.B2(I3[28]),
		.Z(O1[28])
	);
	AO_CELL inst_2_28(
		.A1(out_sel[4]),
		.A2(I4[28]),
		.B1(out_sel[5]),
		.B2(I5[28]),
		.Z(O2[28])
	);
	AN_CELL inst_and_28(
		.A1(out_sel[6]),
		.A2(I6[28]),
		.Z(O3[28])
	);
	AO_CELL inst_0_29(
		.A1(out_sel[0]),
		.A2(I0[29]),
		.B1(out_sel[1]),
		.B2(I1[29]),
		.Z(O0[29])
	);
	AO_CELL inst_1_29(
		.A1(out_sel[2]),
		.A2(I2[29]),
		.B1(out_sel[3]),
		.B2(I3[29]),
		.Z(O1[29])
	);
	AO_CELL inst_2_29(
		.A1(out_sel[4]),
		.A2(I4[29]),
		.B1(out_sel[5]),
		.B2(I5[29]),
		.Z(O2[29])
	);
	AN_CELL inst_and_29(
		.A1(out_sel[6]),
		.A2(I6[29]),
		.Z(O3[29])
	);
	AO_CELL inst_0_30(
		.A1(out_sel[0]),
		.A2(I0[30]),
		.B1(out_sel[1]),
		.B2(I1[30]),
		.Z(O0[30])
	);
	AO_CELL inst_1_30(
		.A1(out_sel[2]),
		.A2(I2[30]),
		.B1(out_sel[3]),
		.B2(I3[30]),
		.Z(O1[30])
	);
	AO_CELL inst_2_30(
		.A1(out_sel[4]),
		.A2(I4[30]),
		.B1(out_sel[5]),
		.B2(I5[30]),
		.Z(O2[30])
	);
	AN_CELL inst_and_30(
		.A1(out_sel[6]),
		.A2(I6[30]),
		.Z(O3[30])
	);
	AO_CELL inst_0_31(
		.A1(out_sel[0]),
		.A2(I0[31]),
		.B1(out_sel[1]),
		.B2(I1[31]),
		.Z(O0[31])
	);
	AO_CELL inst_1_31(
		.A1(out_sel[2]),
		.A2(I2[31]),
		.B1(out_sel[3]),
		.B2(I3[31]),
		.Z(O1[31])
	);
	AO_CELL inst_2_31(
		.A1(out_sel[4]),
		.A2(I4[31]),
		.B1(out_sel[5]),
		.B2(I5[31]),
		.Z(O2[31])
	);
	AN_CELL inst_and_31(
		.A1(out_sel[6]),
		.A2(I6[31]),
		.Z(O3[31])
	);
endmodule
module mux_aoi_6_32 (
	I,
	S,
	out_sel,
	O
);
	input wire [191:0] I;
	input wire [2:0] S;
	output wire [7:0] out_sel;
	output wire [31:0] O;
	wire [31:0] O_int0;
	wire [31:0] O_int1;
	wire [31:0] O_int2;
	precoder_32_6 u_precoder(
		.S(S),
		.out_sel(out_sel)
	);
	mux_logic_32_6 u_mux_logic(
		.I0(I[0+:32]),
		.I1(I[32+:32]),
		.I2(I[64+:32]),
		.I3(I[96+:32]),
		.I4(I[128+:32]),
		.I5(I[160+:32]),
		.out_sel(out_sel),
		.O0(O_int0),
		.O1(O_int1),
		.O2(O_int2)
	);
	assign O = (O_int0 | O_int1) | O_int2;
endmodule
module precoder_32_6 (
	S,
	out_sel
);
	input wire [2:0] S;
	output reg [7:0] out_sel;
	always @(*) begin : mux_sel
		case (S)
			3'd0: out_sel = 8'b00000001;
			3'd1: out_sel = 8'b00000010;
			3'd2: out_sel = 8'b00000100;
			3'd3: out_sel = 8'b00001000;
			3'd4: out_sel = 8'b00010000;
			3'd5: out_sel = 8'b00100000;
			default: out_sel = 8'b00000000;
		endcase
	end
endmodule
module mux_logic_32_6 (
	out_sel,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	O0,
	O1,
	O2
);
	input wire [7:0] out_sel;
	input wire [31:0] I0;
	input wire [31:0] I1;
	input wire [31:0] I2;
	input wire [31:0] I3;
	input wire [31:0] I4;
	input wire [31:0] I5;
	output wire [31:0] O0;
	output wire [31:0] O1;
	output wire [31:0] O2;
	AO_CELL inst_0_0(
		.A1(out_sel[0]),
		.A2(I0[0]),
		.B1(out_sel[1]),
		.B2(I1[0]),
		.Z(O0[0])
	);
	AO_CELL inst_1_0(
		.A1(out_sel[2]),
		.A2(I2[0]),
		.B1(out_sel[3]),
		.B2(I3[0]),
		.Z(O1[0])
	);
	AO_CELL inst_2_0(
		.A1(out_sel[4]),
		.A2(I4[0]),
		.B1(out_sel[5]),
		.B2(I5[0]),
		.Z(O2[0])
	);
	AO_CELL inst_0_1(
		.A1(out_sel[0]),
		.A2(I0[1]),
		.B1(out_sel[1]),
		.B2(I1[1]),
		.Z(O0[1])
	);
	AO_CELL inst_1_1(
		.A1(out_sel[2]),
		.A2(I2[1]),
		.B1(out_sel[3]),
		.B2(I3[1]),
		.Z(O1[1])
	);
	AO_CELL inst_2_1(
		.A1(out_sel[4]),
		.A2(I4[1]),
		.B1(out_sel[5]),
		.B2(I5[1]),
		.Z(O2[1])
	);
	AO_CELL inst_0_2(
		.A1(out_sel[0]),
		.A2(I0[2]),
		.B1(out_sel[1]),
		.B2(I1[2]),
		.Z(O0[2])
	);
	AO_CELL inst_1_2(
		.A1(out_sel[2]),
		.A2(I2[2]),
		.B1(out_sel[3]),
		.B2(I3[2]),
		.Z(O1[2])
	);
	AO_CELL inst_2_2(
		.A1(out_sel[4]),
		.A2(I4[2]),
		.B1(out_sel[5]),
		.B2(I5[2]),
		.Z(O2[2])
	);
	AO_CELL inst_0_3(
		.A1(out_sel[0]),
		.A2(I0[3]),
		.B1(out_sel[1]),
		.B2(I1[3]),
		.Z(O0[3])
	);
	AO_CELL inst_1_3(
		.A1(out_sel[2]),
		.A2(I2[3]),
		.B1(out_sel[3]),
		.B2(I3[3]),
		.Z(O1[3])
	);
	AO_CELL inst_2_3(
		.A1(out_sel[4]),
		.A2(I4[3]),
		.B1(out_sel[5]),
		.B2(I5[3]),
		.Z(O2[3])
	);
	AO_CELL inst_0_4(
		.A1(out_sel[0]),
		.A2(I0[4]),
		.B1(out_sel[1]),
		.B2(I1[4]),
		.Z(O0[4])
	);
	AO_CELL inst_1_4(
		.A1(out_sel[2]),
		.A2(I2[4]),
		.B1(out_sel[3]),
		.B2(I3[4]),
		.Z(O1[4])
	);
	AO_CELL inst_2_4(
		.A1(out_sel[4]),
		.A2(I4[4]),
		.B1(out_sel[5]),
		.B2(I5[4]),
		.Z(O2[4])
	);
	AO_CELL inst_0_5(
		.A1(out_sel[0]),
		.A2(I0[5]),
		.B1(out_sel[1]),
		.B2(I1[5]),
		.Z(O0[5])
	);
	AO_CELL inst_1_5(
		.A1(out_sel[2]),
		.A2(I2[5]),
		.B1(out_sel[3]),
		.B2(I3[5]),
		.Z(O1[5])
	);
	AO_CELL inst_2_5(
		.A1(out_sel[4]),
		.A2(I4[5]),
		.B1(out_sel[5]),
		.B2(I5[5]),
		.Z(O2[5])
	);
	AO_CELL inst_0_6(
		.A1(out_sel[0]),
		.A2(I0[6]),
		.B1(out_sel[1]),
		.B2(I1[6]),
		.Z(O0[6])
	);
	AO_CELL inst_1_6(
		.A1(out_sel[2]),
		.A2(I2[6]),
		.B1(out_sel[3]),
		.B2(I3[6]),
		.Z(O1[6])
	);
	AO_CELL inst_2_6(
		.A1(out_sel[4]),
		.A2(I4[6]),
		.B1(out_sel[5]),
		.B2(I5[6]),
		.Z(O2[6])
	);
	AO_CELL inst_0_7(
		.A1(out_sel[0]),
		.A2(I0[7]),
		.B1(out_sel[1]),
		.B2(I1[7]),
		.Z(O0[7])
	);
	AO_CELL inst_1_7(
		.A1(out_sel[2]),
		.A2(I2[7]),
		.B1(out_sel[3]),
		.B2(I3[7]),
		.Z(O1[7])
	);
	AO_CELL inst_2_7(
		.A1(out_sel[4]),
		.A2(I4[7]),
		.B1(out_sel[5]),
		.B2(I5[7]),
		.Z(O2[7])
	);
	AO_CELL inst_0_8(
		.A1(out_sel[0]),
		.A2(I0[8]),
		.B1(out_sel[1]),
		.B2(I1[8]),
		.Z(O0[8])
	);
	AO_CELL inst_1_8(
		.A1(out_sel[2]),
		.A2(I2[8]),
		.B1(out_sel[3]),
		.B2(I3[8]),
		.Z(O1[8])
	);
	AO_CELL inst_2_8(
		.A1(out_sel[4]),
		.A2(I4[8]),
		.B1(out_sel[5]),
		.B2(I5[8]),
		.Z(O2[8])
	);
	AO_CELL inst_0_9(
		.A1(out_sel[0]),
		.A2(I0[9]),
		.B1(out_sel[1]),
		.B2(I1[9]),
		.Z(O0[9])
	);
	AO_CELL inst_1_9(
		.A1(out_sel[2]),
		.A2(I2[9]),
		.B1(out_sel[3]),
		.B2(I3[9]),
		.Z(O1[9])
	);
	AO_CELL inst_2_9(
		.A1(out_sel[4]),
		.A2(I4[9]),
		.B1(out_sel[5]),
		.B2(I5[9]),
		.Z(O2[9])
	);
	AO_CELL inst_0_10(
		.A1(out_sel[0]),
		.A2(I0[10]),
		.B1(out_sel[1]),
		.B2(I1[10]),
		.Z(O0[10])
	);
	AO_CELL inst_1_10(
		.A1(out_sel[2]),
		.A2(I2[10]),
		.B1(out_sel[3]),
		.B2(I3[10]),
		.Z(O1[10])
	);
	AO_CELL inst_2_10(
		.A1(out_sel[4]),
		.A2(I4[10]),
		.B1(out_sel[5]),
		.B2(I5[10]),
		.Z(O2[10])
	);
	AO_CELL inst_0_11(
		.A1(out_sel[0]),
		.A2(I0[11]),
		.B1(out_sel[1]),
		.B2(I1[11]),
		.Z(O0[11])
	);
	AO_CELL inst_1_11(
		.A1(out_sel[2]),
		.A2(I2[11]),
		.B1(out_sel[3]),
		.B2(I3[11]),
		.Z(O1[11])
	);
	AO_CELL inst_2_11(
		.A1(out_sel[4]),
		.A2(I4[11]),
		.B1(out_sel[5]),
		.B2(I5[11]),
		.Z(O2[11])
	);
	AO_CELL inst_0_12(
		.A1(out_sel[0]),
		.A2(I0[12]),
		.B1(out_sel[1]),
		.B2(I1[12]),
		.Z(O0[12])
	);
	AO_CELL inst_1_12(
		.A1(out_sel[2]),
		.A2(I2[12]),
		.B1(out_sel[3]),
		.B2(I3[12]),
		.Z(O1[12])
	);
	AO_CELL inst_2_12(
		.A1(out_sel[4]),
		.A2(I4[12]),
		.B1(out_sel[5]),
		.B2(I5[12]),
		.Z(O2[12])
	);
	AO_CELL inst_0_13(
		.A1(out_sel[0]),
		.A2(I0[13]),
		.B1(out_sel[1]),
		.B2(I1[13]),
		.Z(O0[13])
	);
	AO_CELL inst_1_13(
		.A1(out_sel[2]),
		.A2(I2[13]),
		.B1(out_sel[3]),
		.B2(I3[13]),
		.Z(O1[13])
	);
	AO_CELL inst_2_13(
		.A1(out_sel[4]),
		.A2(I4[13]),
		.B1(out_sel[5]),
		.B2(I5[13]),
		.Z(O2[13])
	);
	AO_CELL inst_0_14(
		.A1(out_sel[0]),
		.A2(I0[14]),
		.B1(out_sel[1]),
		.B2(I1[14]),
		.Z(O0[14])
	);
	AO_CELL inst_1_14(
		.A1(out_sel[2]),
		.A2(I2[14]),
		.B1(out_sel[3]),
		.B2(I3[14]),
		.Z(O1[14])
	);
	AO_CELL inst_2_14(
		.A1(out_sel[4]),
		.A2(I4[14]),
		.B1(out_sel[5]),
		.B2(I5[14]),
		.Z(O2[14])
	);
	AO_CELL inst_0_15(
		.A1(out_sel[0]),
		.A2(I0[15]),
		.B1(out_sel[1]),
		.B2(I1[15]),
		.Z(O0[15])
	);
	AO_CELL inst_1_15(
		.A1(out_sel[2]),
		.A2(I2[15]),
		.B1(out_sel[3]),
		.B2(I3[15]),
		.Z(O1[15])
	);
	AO_CELL inst_2_15(
		.A1(out_sel[4]),
		.A2(I4[15]),
		.B1(out_sel[5]),
		.B2(I5[15]),
		.Z(O2[15])
	);
	AO_CELL inst_0_16(
		.A1(out_sel[0]),
		.A2(I0[16]),
		.B1(out_sel[1]),
		.B2(I1[16]),
		.Z(O0[16])
	);
	AO_CELL inst_1_16(
		.A1(out_sel[2]),
		.A2(I2[16]),
		.B1(out_sel[3]),
		.B2(I3[16]),
		.Z(O1[16])
	);
	AO_CELL inst_2_16(
		.A1(out_sel[4]),
		.A2(I4[16]),
		.B1(out_sel[5]),
		.B2(I5[16]),
		.Z(O2[16])
	);
	AO_CELL inst_0_17(
		.A1(out_sel[0]),
		.A2(I0[17]),
		.B1(out_sel[1]),
		.B2(I1[17]),
		.Z(O0[17])
	);
	AO_CELL inst_1_17(
		.A1(out_sel[2]),
		.A2(I2[17]),
		.B1(out_sel[3]),
		.B2(I3[17]),
		.Z(O1[17])
	);
	AO_CELL inst_2_17(
		.A1(out_sel[4]),
		.A2(I4[17]),
		.B1(out_sel[5]),
		.B2(I5[17]),
		.Z(O2[17])
	);
	AO_CELL inst_0_18(
		.A1(out_sel[0]),
		.A2(I0[18]),
		.B1(out_sel[1]),
		.B2(I1[18]),
		.Z(O0[18])
	);
	AO_CELL inst_1_18(
		.A1(out_sel[2]),
		.A2(I2[18]),
		.B1(out_sel[3]),
		.B2(I3[18]),
		.Z(O1[18])
	);
	AO_CELL inst_2_18(
		.A1(out_sel[4]),
		.A2(I4[18]),
		.B1(out_sel[5]),
		.B2(I5[18]),
		.Z(O2[18])
	);
	AO_CELL inst_0_19(
		.A1(out_sel[0]),
		.A2(I0[19]),
		.B1(out_sel[1]),
		.B2(I1[19]),
		.Z(O0[19])
	);
	AO_CELL inst_1_19(
		.A1(out_sel[2]),
		.A2(I2[19]),
		.B1(out_sel[3]),
		.B2(I3[19]),
		.Z(O1[19])
	);
	AO_CELL inst_2_19(
		.A1(out_sel[4]),
		.A2(I4[19]),
		.B1(out_sel[5]),
		.B2(I5[19]),
		.Z(O2[19])
	);
	AO_CELL inst_0_20(
		.A1(out_sel[0]),
		.A2(I0[20]),
		.B1(out_sel[1]),
		.B2(I1[20]),
		.Z(O0[20])
	);
	AO_CELL inst_1_20(
		.A1(out_sel[2]),
		.A2(I2[20]),
		.B1(out_sel[3]),
		.B2(I3[20]),
		.Z(O1[20])
	);
	AO_CELL inst_2_20(
		.A1(out_sel[4]),
		.A2(I4[20]),
		.B1(out_sel[5]),
		.B2(I5[20]),
		.Z(O2[20])
	);
	AO_CELL inst_0_21(
		.A1(out_sel[0]),
		.A2(I0[21]),
		.B1(out_sel[1]),
		.B2(I1[21]),
		.Z(O0[21])
	);
	AO_CELL inst_1_21(
		.A1(out_sel[2]),
		.A2(I2[21]),
		.B1(out_sel[3]),
		.B2(I3[21]),
		.Z(O1[21])
	);
	AO_CELL inst_2_21(
		.A1(out_sel[4]),
		.A2(I4[21]),
		.B1(out_sel[5]),
		.B2(I5[21]),
		.Z(O2[21])
	);
	AO_CELL inst_0_22(
		.A1(out_sel[0]),
		.A2(I0[22]),
		.B1(out_sel[1]),
		.B2(I1[22]),
		.Z(O0[22])
	);
	AO_CELL inst_1_22(
		.A1(out_sel[2]),
		.A2(I2[22]),
		.B1(out_sel[3]),
		.B2(I3[22]),
		.Z(O1[22])
	);
	AO_CELL inst_2_22(
		.A1(out_sel[4]),
		.A2(I4[22]),
		.B1(out_sel[5]),
		.B2(I5[22]),
		.Z(O2[22])
	);
	AO_CELL inst_0_23(
		.A1(out_sel[0]),
		.A2(I0[23]),
		.B1(out_sel[1]),
		.B2(I1[23]),
		.Z(O0[23])
	);
	AO_CELL inst_1_23(
		.A1(out_sel[2]),
		.A2(I2[23]),
		.B1(out_sel[3]),
		.B2(I3[23]),
		.Z(O1[23])
	);
	AO_CELL inst_2_23(
		.A1(out_sel[4]),
		.A2(I4[23]),
		.B1(out_sel[5]),
		.B2(I5[23]),
		.Z(O2[23])
	);
	AO_CELL inst_0_24(
		.A1(out_sel[0]),
		.A2(I0[24]),
		.B1(out_sel[1]),
		.B2(I1[24]),
		.Z(O0[24])
	);
	AO_CELL inst_1_24(
		.A1(out_sel[2]),
		.A2(I2[24]),
		.B1(out_sel[3]),
		.B2(I3[24]),
		.Z(O1[24])
	);
	AO_CELL inst_2_24(
		.A1(out_sel[4]),
		.A2(I4[24]),
		.B1(out_sel[5]),
		.B2(I5[24]),
		.Z(O2[24])
	);
	AO_CELL inst_0_25(
		.A1(out_sel[0]),
		.A2(I0[25]),
		.B1(out_sel[1]),
		.B2(I1[25]),
		.Z(O0[25])
	);
	AO_CELL inst_1_25(
		.A1(out_sel[2]),
		.A2(I2[25]),
		.B1(out_sel[3]),
		.B2(I3[25]),
		.Z(O1[25])
	);
	AO_CELL inst_2_25(
		.A1(out_sel[4]),
		.A2(I4[25]),
		.B1(out_sel[5]),
		.B2(I5[25]),
		.Z(O2[25])
	);
	AO_CELL inst_0_26(
		.A1(out_sel[0]),
		.A2(I0[26]),
		.B1(out_sel[1]),
		.B2(I1[26]),
		.Z(O0[26])
	);
	AO_CELL inst_1_26(
		.A1(out_sel[2]),
		.A2(I2[26]),
		.B1(out_sel[3]),
		.B2(I3[26]),
		.Z(O1[26])
	);
	AO_CELL inst_2_26(
		.A1(out_sel[4]),
		.A2(I4[26]),
		.B1(out_sel[5]),
		.B2(I5[26]),
		.Z(O2[26])
	);
	AO_CELL inst_0_27(
		.A1(out_sel[0]),
		.A2(I0[27]),
		.B1(out_sel[1]),
		.B2(I1[27]),
		.Z(O0[27])
	);
	AO_CELL inst_1_27(
		.A1(out_sel[2]),
		.A2(I2[27]),
		.B1(out_sel[3]),
		.B2(I3[27]),
		.Z(O1[27])
	);
	AO_CELL inst_2_27(
		.A1(out_sel[4]),
		.A2(I4[27]),
		.B1(out_sel[5]),
		.B2(I5[27]),
		.Z(O2[27])
	);
	AO_CELL inst_0_28(
		.A1(out_sel[0]),
		.A2(I0[28]),
		.B1(out_sel[1]),
		.B2(I1[28]),
		.Z(O0[28])
	);
	AO_CELL inst_1_28(
		.A1(out_sel[2]),
		.A2(I2[28]),
		.B1(out_sel[3]),
		.B2(I3[28]),
		.Z(O1[28])
	);
	AO_CELL inst_2_28(
		.A1(out_sel[4]),
		.A2(I4[28]),
		.B1(out_sel[5]),
		.B2(I5[28]),
		.Z(O2[28])
	);
	AO_CELL inst_0_29(
		.A1(out_sel[0]),
		.A2(I0[29]),
		.B1(out_sel[1]),
		.B2(I1[29]),
		.Z(O0[29])
	);
	AO_CELL inst_1_29(
		.A1(out_sel[2]),
		.A2(I2[29]),
		.B1(out_sel[3]),
		.B2(I3[29]),
		.Z(O1[29])
	);
	AO_CELL inst_2_29(
		.A1(out_sel[4]),
		.A2(I4[29]),
		.B1(out_sel[5]),
		.B2(I5[29]),
		.Z(O2[29])
	);
	AO_CELL inst_0_30(
		.A1(out_sel[0]),
		.A2(I0[30]),
		.B1(out_sel[1]),
		.B2(I1[30]),
		.Z(O0[30])
	);
	AO_CELL inst_1_30(
		.A1(out_sel[2]),
		.A2(I2[30]),
		.B1(out_sel[3]),
		.B2(I3[30]),
		.Z(O1[30])
	);
	AO_CELL inst_2_30(
		.A1(out_sel[4]),
		.A2(I4[30]),
		.B1(out_sel[5]),
		.B2(I5[30]),
		.Z(O2[30])
	);
	AO_CELL inst_0_31(
		.A1(out_sel[0]),
		.A2(I0[31]),
		.B1(out_sel[1]),
		.B2(I1[31]),
		.Z(O0[31])
	);
	AO_CELL inst_1_31(
		.A1(out_sel[2]),
		.A2(I2[31]),
		.B1(out_sel[3]),
		.B2(I3[31]),
		.Z(O1[31])
	);
	AO_CELL inst_2_31(
		.A1(out_sel[4]),
		.A2(I4[31]),
		.B1(out_sel[5]),
		.B2(I5[31]),
		.Z(O2[31])
	);
endmodule
module mux_aoi_47_32 (
	I,
	S,
	out_sel,
	O
);
	input wire [1503:0] I;
	input wire [5:0] S;
	output wire [63:0] out_sel;
	output wire [31:0] O;
	wire [31:0] O_int0;
	wire [31:0] O_int1;
	wire [31:0] O_int2;
	wire [31:0] O_int3;
	wire [31:0] O_int4;
	wire [31:0] O_int5;
	wire [31:0] O_int6;
	wire [31:0] O_int7;
	wire [31:0] O_int8;
	wire [31:0] O_int9;
	wire [31:0] O_int10;
	wire [31:0] O_int11;
	wire [31:0] O_int12;
	wire [31:0] O_int13;
	wire [31:0] O_int14;
	wire [31:0] O_int15;
	wire [31:0] O_int16;
	wire [31:0] O_int17;
	wire [31:0] O_int18;
	wire [31:0] O_int19;
	wire [31:0] O_int20;
	wire [31:0] O_int21;
	wire [31:0] O_int22;
	wire [31:0] O_int23;
	precoder_32_47 u_precoder(
		.S(S),
		.out_sel(out_sel)
	);
	mux_logic_32_47 u_mux_logic(
		.I0(I[0+:32]),
		.I1(I[32+:32]),
		.I2(I[64+:32]),
		.I3(I[96+:32]),
		.I4(I[128+:32]),
		.I5(I[160+:32]),
		.I6(I[192+:32]),
		.I7(I[224+:32]),
		.I8(I[256+:32]),
		.I9(I[288+:32]),
		.I10(I[320+:32]),
		.I11(I[352+:32]),
		.I12(I[384+:32]),
		.I13(I[416+:32]),
		.I14(I[448+:32]),
		.I15(I[480+:32]),
		.I16(I[512+:32]),
		.I17(I[544+:32]),
		.I18(I[576+:32]),
		.I19(I[608+:32]),
		.I20(I[640+:32]),
		.I21(I[672+:32]),
		.I22(I[704+:32]),
		.I23(I[736+:32]),
		.I24(I[768+:32]),
		.I25(I[800+:32]),
		.I26(I[832+:32]),
		.I27(I[864+:32]),
		.I28(I[896+:32]),
		.I29(I[928+:32]),
		.I30(I[960+:32]),
		.I31(I[992+:32]),
		.I32(I[1024+:32]),
		.I33(I[1056+:32]),
		.I34(I[1088+:32]),
		.I35(I[1120+:32]),
		.I36(I[1152+:32]),
		.I37(I[1184+:32]),
		.I38(I[1216+:32]),
		.I39(I[1248+:32]),
		.I40(I[1280+:32]),
		.I41(I[1312+:32]),
		.I42(I[1344+:32]),
		.I43(I[1376+:32]),
		.I44(I[1408+:32]),
		.I45(I[1440+:32]),
		.I46(I[1472+:32]),
		.out_sel(out_sel),
		.O0(O_int0),
		.O1(O_int1),
		.O2(O_int2),
		.O3(O_int3),
		.O4(O_int4),
		.O5(O_int5),
		.O6(O_int6),
		.O7(O_int7),
		.O8(O_int8),
		.O9(O_int9),
		.O10(O_int10),
		.O11(O_int11),
		.O12(O_int12),
		.O13(O_int13),
		.O14(O_int14),
		.O15(O_int15),
		.O16(O_int16),
		.O17(O_int17),
		.O18(O_int18),
		.O19(O_int19),
		.O20(O_int20),
		.O21(O_int21),
		.O22(O_int22),
		.O23(O_int23)
	);
	assign O = ((((((((((((((((((((((O_int0 | O_int1) | O_int2) | O_int3) | O_int4) | O_int5) | O_int6) | O_int7) | O_int8) | O_int9) | O_int10) | O_int11) | O_int12) | O_int13) | O_int14) | O_int15) | O_int16) | O_int17) | O_int18) | O_int19) | O_int20) | O_int21) | O_int22) | O_int23;
endmodule
module precoder_32_47 (
	S,
	out_sel
);
	input wire [5:0] S;
	output reg [63:0] out_sel;
	always @(*) begin : mux_sel
		case (S)
			6'd0: out_sel = 64'b0000000000000000000000000000000000000000000000000000000000000001;
			6'd1: out_sel = 64'b0000000000000000000000000000000000000000000000000000000000000010;
			6'd2: out_sel = 64'b0000000000000000000000000000000000000000000000000000000000000100;
			6'd3: out_sel = 64'b0000000000000000000000000000000000000000000000000000000000001000;
			6'd4: out_sel = 64'b0000000000000000000000000000000000000000000000000000000000010000;
			6'd5: out_sel = 64'b0000000000000000000000000000000000000000000000000000000000100000;
			6'd6: out_sel = 64'b0000000000000000000000000000000000000000000000000000000001000000;
			6'd7: out_sel = 64'b0000000000000000000000000000000000000000000000000000000010000000;
			6'd8: out_sel = 64'b0000000000000000000000000000000000000000000000000000000100000000;
			6'd9: out_sel = 64'b0000000000000000000000000000000000000000000000000000001000000000;
			6'd10: out_sel = 64'b0000000000000000000000000000000000000000000000000000010000000000;
			6'd11: out_sel = 64'b0000000000000000000000000000000000000000000000000000100000000000;
			6'd12: out_sel = 64'b0000000000000000000000000000000000000000000000000001000000000000;
			6'd13: out_sel = 64'b0000000000000000000000000000000000000000000000000010000000000000;
			6'd14: out_sel = 64'b0000000000000000000000000000000000000000000000000100000000000000;
			6'd15: out_sel = 64'b0000000000000000000000000000000000000000000000001000000000000000;
			6'd16: out_sel = 64'b0000000000000000000000000000000000000000000000010000000000000000;
			6'd17: out_sel = 64'b0000000000000000000000000000000000000000000000100000000000000000;
			6'd18: out_sel = 64'b0000000000000000000000000000000000000000000001000000000000000000;
			6'd19: out_sel = 64'b0000000000000000000000000000000000000000000010000000000000000000;
			6'd20: out_sel = 64'b0000000000000000000000000000000000000000000100000000000000000000;
			6'd21: out_sel = 64'b0000000000000000000000000000000000000000001000000000000000000000;
			6'd22: out_sel = 64'b0000000000000000000000000000000000000000010000000000000000000000;
			6'd23: out_sel = 64'b0000000000000000000000000000000000000000100000000000000000000000;
			6'd24: out_sel = 64'b0000000000000000000000000000000000000001000000000000000000000000;
			6'd25: out_sel = 64'b0000000000000000000000000000000000000010000000000000000000000000;
			6'd26: out_sel = 64'b0000000000000000000000000000000000000100000000000000000000000000;
			6'd27: out_sel = 64'b0000000000000000000000000000000000001000000000000000000000000000;
			6'd28: out_sel = 64'b0000000000000000000000000000000000010000000000000000000000000000;
			6'd29: out_sel = 64'b0000000000000000000000000000000000100000000000000000000000000000;
			6'd30: out_sel = 64'b0000000000000000000000000000000001000000000000000000000000000000;
			6'd31: out_sel = 64'b0000000000000000000000000000000010000000000000000000000000000000;
			6'd32: out_sel = 64'b0000000000000000000000000000000100000000000000000000000000000000;
			6'd33: out_sel = 64'b0000000000000000000000000000001000000000000000000000000000000000;
			6'd34: out_sel = 64'b0000000000000000000000000000010000000000000000000000000000000000;
			6'd35: out_sel = 64'b0000000000000000000000000000100000000000000000000000000000000000;
			6'd36: out_sel = 64'b0000000000000000000000000001000000000000000000000000000000000000;
			6'd37: out_sel = 64'b0000000000000000000000000010000000000000000000000000000000000000;
			6'd38: out_sel = 64'b0000000000000000000000000100000000000000000000000000000000000000;
			6'd39: out_sel = 64'b0000000000000000000000001000000000000000000000000000000000000000;
			6'd40: out_sel = 64'b0000000000000000000000010000000000000000000000000000000000000000;
			6'd41: out_sel = 64'b0000000000000000000000100000000000000000000000000000000000000000;
			6'd42: out_sel = 64'b0000000000000000000001000000000000000000000000000000000000000000;
			6'd43: out_sel = 64'b0000000000000000000010000000000000000000000000000000000000000000;
			6'd44: out_sel = 64'b0000000000000000000100000000000000000000000000000000000000000000;
			6'd45: out_sel = 64'b0000000000000000001000000000000000000000000000000000000000000000;
			6'd46: out_sel = 64'b0000000000000000010000000000000000000000000000000000000000000000;
			default: out_sel = 64'b0000000000000000000000000000000000000000000000000000000000000000;
		endcase
	end
endmodule
module mux_logic_32_47 (
	out_sel,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	I9,
	I10,
	I11,
	I12,
	I13,
	I14,
	I15,
	I16,
	I17,
	I18,
	I19,
	I20,
	I21,
	I22,
	I23,
	I24,
	I25,
	I26,
	I27,
	I28,
	I29,
	I30,
	I31,
	I32,
	I33,
	I34,
	I35,
	I36,
	I37,
	I38,
	I39,
	I40,
	I41,
	I42,
	I43,
	I44,
	I45,
	I46,
	O0,
	O1,
	O2,
	O3,
	O4,
	O5,
	O6,
	O7,
	O8,
	O9,
	O10,
	O11,
	O12,
	O13,
	O14,
	O15,
	O16,
	O17,
	O18,
	O19,
	O20,
	O21,
	O22,
	O23
);
	input wire [63:0] out_sel;
	input wire [31:0] I0;
	input wire [31:0] I1;
	input wire [31:0] I2;
	input wire [31:0] I3;
	input wire [31:0] I4;
	input wire [31:0] I5;
	input wire [31:0] I6;
	input wire [31:0] I7;
	input wire [31:0] I8;
	input wire [31:0] I9;
	input wire [31:0] I10;
	input wire [31:0] I11;
	input wire [31:0] I12;
	input wire [31:0] I13;
	input wire [31:0] I14;
	input wire [31:0] I15;
	input wire [31:0] I16;
	input wire [31:0] I17;
	input wire [31:0] I18;
	input wire [31:0] I19;
	input wire [31:0] I20;
	input wire [31:0] I21;
	input wire [31:0] I22;
	input wire [31:0] I23;
	input wire [31:0] I24;
	input wire [31:0] I25;
	input wire [31:0] I26;
	input wire [31:0] I27;
	input wire [31:0] I28;
	input wire [31:0] I29;
	input wire [31:0] I30;
	input wire [31:0] I31;
	input wire [31:0] I32;
	input wire [31:0] I33;
	input wire [31:0] I34;
	input wire [31:0] I35;
	input wire [31:0] I36;
	input wire [31:0] I37;
	input wire [31:0] I38;
	input wire [31:0] I39;
	input wire [31:0] I40;
	input wire [31:0] I41;
	input wire [31:0] I42;
	input wire [31:0] I43;
	input wire [31:0] I44;
	input wire [31:0] I45;
	input wire [31:0] I46;
	output wire [31:0] O0;
	output wire [31:0] O1;
	output wire [31:0] O2;
	output wire [31:0] O3;
	output wire [31:0] O4;
	output wire [31:0] O5;
	output wire [31:0] O6;
	output wire [31:0] O7;
	output wire [31:0] O8;
	output wire [31:0] O9;
	output wire [31:0] O10;
	output wire [31:0] O11;
	output wire [31:0] O12;
	output wire [31:0] O13;
	output wire [31:0] O14;
	output wire [31:0] O15;
	output wire [31:0] O16;
	output wire [31:0] O17;
	output wire [31:0] O18;
	output wire [31:0] O19;
	output wire [31:0] O20;
	output wire [31:0] O21;
	output wire [31:0] O22;
	output wire [31:0] O23;
	AO_CELL inst_0_0(
		.A1(out_sel[0]),
		.A2(I0[0]),
		.B1(out_sel[1]),
		.B2(I1[0]),
		.Z(O0[0])
	);
	AO_CELL inst_1_0(
		.A1(out_sel[2]),
		.A2(I2[0]),
		.B1(out_sel[3]),
		.B2(I3[0]),
		.Z(O1[0])
	);
	AO_CELL inst_2_0(
		.A1(out_sel[4]),
		.A2(I4[0]),
		.B1(out_sel[5]),
		.B2(I5[0]),
		.Z(O2[0])
	);
	AO_CELL inst_3_0(
		.A1(out_sel[6]),
		.A2(I6[0]),
		.B1(out_sel[7]),
		.B2(I7[0]),
		.Z(O3[0])
	);
	AO_CELL inst_4_0(
		.A1(out_sel[8]),
		.A2(I8[0]),
		.B1(out_sel[9]),
		.B2(I9[0]),
		.Z(O4[0])
	);
	AO_CELL inst_5_0(
		.A1(out_sel[10]),
		.A2(I10[0]),
		.B1(out_sel[11]),
		.B2(I11[0]),
		.Z(O5[0])
	);
	AO_CELL inst_6_0(
		.A1(out_sel[12]),
		.A2(I12[0]),
		.B1(out_sel[13]),
		.B2(I13[0]),
		.Z(O6[0])
	);
	AO_CELL inst_7_0(
		.A1(out_sel[14]),
		.A2(I14[0]),
		.B1(out_sel[15]),
		.B2(I15[0]),
		.Z(O7[0])
	);
	AO_CELL inst_8_0(
		.A1(out_sel[16]),
		.A2(I16[0]),
		.B1(out_sel[17]),
		.B2(I17[0]),
		.Z(O8[0])
	);
	AO_CELL inst_9_0(
		.A1(out_sel[18]),
		.A2(I18[0]),
		.B1(out_sel[19]),
		.B2(I19[0]),
		.Z(O9[0])
	);
	AO_CELL inst_10_0(
		.A1(out_sel[20]),
		.A2(I20[0]),
		.B1(out_sel[21]),
		.B2(I21[0]),
		.Z(O10[0])
	);
	AO_CELL inst_11_0(
		.A1(out_sel[22]),
		.A2(I22[0]),
		.B1(out_sel[23]),
		.B2(I23[0]),
		.Z(O11[0])
	);
	AO_CELL inst_12_0(
		.A1(out_sel[24]),
		.A2(I24[0]),
		.B1(out_sel[25]),
		.B2(I25[0]),
		.Z(O12[0])
	);
	AO_CELL inst_13_0(
		.A1(out_sel[26]),
		.A2(I26[0]),
		.B1(out_sel[27]),
		.B2(I27[0]),
		.Z(O13[0])
	);
	AO_CELL inst_14_0(
		.A1(out_sel[28]),
		.A2(I28[0]),
		.B1(out_sel[29]),
		.B2(I29[0]),
		.Z(O14[0])
	);
	AO_CELL inst_15_0(
		.A1(out_sel[30]),
		.A2(I30[0]),
		.B1(out_sel[31]),
		.B2(I31[0]),
		.Z(O15[0])
	);
	AO_CELL inst_16_0(
		.A1(out_sel[32]),
		.A2(I32[0]),
		.B1(out_sel[33]),
		.B2(I33[0]),
		.Z(O16[0])
	);
	AO_CELL inst_17_0(
		.A1(out_sel[34]),
		.A2(I34[0]),
		.B1(out_sel[35]),
		.B2(I35[0]),
		.Z(O17[0])
	);
	AO_CELL inst_18_0(
		.A1(out_sel[36]),
		.A2(I36[0]),
		.B1(out_sel[37]),
		.B2(I37[0]),
		.Z(O18[0])
	);
	AO_CELL inst_19_0(
		.A1(out_sel[38]),
		.A2(I38[0]),
		.B1(out_sel[39]),
		.B2(I39[0]),
		.Z(O19[0])
	);
	AO_CELL inst_20_0(
		.A1(out_sel[40]),
		.A2(I40[0]),
		.B1(out_sel[41]),
		.B2(I41[0]),
		.Z(O20[0])
	);
	AO_CELL inst_21_0(
		.A1(out_sel[42]),
		.A2(I42[0]),
		.B1(out_sel[43]),
		.B2(I43[0]),
		.Z(O21[0])
	);
	AO_CELL inst_22_0(
		.A1(out_sel[44]),
		.A2(I44[0]),
		.B1(out_sel[45]),
		.B2(I45[0]),
		.Z(O22[0])
	);
	AN_CELL inst_and_0(
		.A1(out_sel[46]),
		.A2(I46[0]),
		.Z(O23[0])
	);
	AO_CELL inst_0_1(
		.A1(out_sel[0]),
		.A2(I0[1]),
		.B1(out_sel[1]),
		.B2(I1[1]),
		.Z(O0[1])
	);
	AO_CELL inst_1_1(
		.A1(out_sel[2]),
		.A2(I2[1]),
		.B1(out_sel[3]),
		.B2(I3[1]),
		.Z(O1[1])
	);
	AO_CELL inst_2_1(
		.A1(out_sel[4]),
		.A2(I4[1]),
		.B1(out_sel[5]),
		.B2(I5[1]),
		.Z(O2[1])
	);
	AO_CELL inst_3_1(
		.A1(out_sel[6]),
		.A2(I6[1]),
		.B1(out_sel[7]),
		.B2(I7[1]),
		.Z(O3[1])
	);
	AO_CELL inst_4_1(
		.A1(out_sel[8]),
		.A2(I8[1]),
		.B1(out_sel[9]),
		.B2(I9[1]),
		.Z(O4[1])
	);
	AO_CELL inst_5_1(
		.A1(out_sel[10]),
		.A2(I10[1]),
		.B1(out_sel[11]),
		.B2(I11[1]),
		.Z(O5[1])
	);
	AO_CELL inst_6_1(
		.A1(out_sel[12]),
		.A2(I12[1]),
		.B1(out_sel[13]),
		.B2(I13[1]),
		.Z(O6[1])
	);
	AO_CELL inst_7_1(
		.A1(out_sel[14]),
		.A2(I14[1]),
		.B1(out_sel[15]),
		.B2(I15[1]),
		.Z(O7[1])
	);
	AO_CELL inst_8_1(
		.A1(out_sel[16]),
		.A2(I16[1]),
		.B1(out_sel[17]),
		.B2(I17[1]),
		.Z(O8[1])
	);
	AO_CELL inst_9_1(
		.A1(out_sel[18]),
		.A2(I18[1]),
		.B1(out_sel[19]),
		.B2(I19[1]),
		.Z(O9[1])
	);
	AO_CELL inst_10_1(
		.A1(out_sel[20]),
		.A2(I20[1]),
		.B1(out_sel[21]),
		.B2(I21[1]),
		.Z(O10[1])
	);
	AO_CELL inst_11_1(
		.A1(out_sel[22]),
		.A2(I22[1]),
		.B1(out_sel[23]),
		.B2(I23[1]),
		.Z(O11[1])
	);
	AO_CELL inst_12_1(
		.A1(out_sel[24]),
		.A2(I24[1]),
		.B1(out_sel[25]),
		.B2(I25[1]),
		.Z(O12[1])
	);
	AO_CELL inst_13_1(
		.A1(out_sel[26]),
		.A2(I26[1]),
		.B1(out_sel[27]),
		.B2(I27[1]),
		.Z(O13[1])
	);
	AO_CELL inst_14_1(
		.A1(out_sel[28]),
		.A2(I28[1]),
		.B1(out_sel[29]),
		.B2(I29[1]),
		.Z(O14[1])
	);
	AO_CELL inst_15_1(
		.A1(out_sel[30]),
		.A2(I30[1]),
		.B1(out_sel[31]),
		.B2(I31[1]),
		.Z(O15[1])
	);
	AO_CELL inst_16_1(
		.A1(out_sel[32]),
		.A2(I32[1]),
		.B1(out_sel[33]),
		.B2(I33[1]),
		.Z(O16[1])
	);
	AO_CELL inst_17_1(
		.A1(out_sel[34]),
		.A2(I34[1]),
		.B1(out_sel[35]),
		.B2(I35[1]),
		.Z(O17[1])
	);
	AO_CELL inst_18_1(
		.A1(out_sel[36]),
		.A2(I36[1]),
		.B1(out_sel[37]),
		.B2(I37[1]),
		.Z(O18[1])
	);
	AO_CELL inst_19_1(
		.A1(out_sel[38]),
		.A2(I38[1]),
		.B1(out_sel[39]),
		.B2(I39[1]),
		.Z(O19[1])
	);
	AO_CELL inst_20_1(
		.A1(out_sel[40]),
		.A2(I40[1]),
		.B1(out_sel[41]),
		.B2(I41[1]),
		.Z(O20[1])
	);
	AO_CELL inst_21_1(
		.A1(out_sel[42]),
		.A2(I42[1]),
		.B1(out_sel[43]),
		.B2(I43[1]),
		.Z(O21[1])
	);
	AO_CELL inst_22_1(
		.A1(out_sel[44]),
		.A2(I44[1]),
		.B1(out_sel[45]),
		.B2(I45[1]),
		.Z(O22[1])
	);
	AN_CELL inst_and_1(
		.A1(out_sel[46]),
		.A2(I46[1]),
		.Z(O23[1])
	);
	AO_CELL inst_0_2(
		.A1(out_sel[0]),
		.A2(I0[2]),
		.B1(out_sel[1]),
		.B2(I1[2]),
		.Z(O0[2])
	);
	AO_CELL inst_1_2(
		.A1(out_sel[2]),
		.A2(I2[2]),
		.B1(out_sel[3]),
		.B2(I3[2]),
		.Z(O1[2])
	);
	AO_CELL inst_2_2(
		.A1(out_sel[4]),
		.A2(I4[2]),
		.B1(out_sel[5]),
		.B2(I5[2]),
		.Z(O2[2])
	);
	AO_CELL inst_3_2(
		.A1(out_sel[6]),
		.A2(I6[2]),
		.B1(out_sel[7]),
		.B2(I7[2]),
		.Z(O3[2])
	);
	AO_CELL inst_4_2(
		.A1(out_sel[8]),
		.A2(I8[2]),
		.B1(out_sel[9]),
		.B2(I9[2]),
		.Z(O4[2])
	);
	AO_CELL inst_5_2(
		.A1(out_sel[10]),
		.A2(I10[2]),
		.B1(out_sel[11]),
		.B2(I11[2]),
		.Z(O5[2])
	);
	AO_CELL inst_6_2(
		.A1(out_sel[12]),
		.A2(I12[2]),
		.B1(out_sel[13]),
		.B2(I13[2]),
		.Z(O6[2])
	);
	AO_CELL inst_7_2(
		.A1(out_sel[14]),
		.A2(I14[2]),
		.B1(out_sel[15]),
		.B2(I15[2]),
		.Z(O7[2])
	);
	AO_CELL inst_8_2(
		.A1(out_sel[16]),
		.A2(I16[2]),
		.B1(out_sel[17]),
		.B2(I17[2]),
		.Z(O8[2])
	);
	AO_CELL inst_9_2(
		.A1(out_sel[18]),
		.A2(I18[2]),
		.B1(out_sel[19]),
		.B2(I19[2]),
		.Z(O9[2])
	);
	AO_CELL inst_10_2(
		.A1(out_sel[20]),
		.A2(I20[2]),
		.B1(out_sel[21]),
		.B2(I21[2]),
		.Z(O10[2])
	);
	AO_CELL inst_11_2(
		.A1(out_sel[22]),
		.A2(I22[2]),
		.B1(out_sel[23]),
		.B2(I23[2]),
		.Z(O11[2])
	);
	AO_CELL inst_12_2(
		.A1(out_sel[24]),
		.A2(I24[2]),
		.B1(out_sel[25]),
		.B2(I25[2]),
		.Z(O12[2])
	);
	AO_CELL inst_13_2(
		.A1(out_sel[26]),
		.A2(I26[2]),
		.B1(out_sel[27]),
		.B2(I27[2]),
		.Z(O13[2])
	);
	AO_CELL inst_14_2(
		.A1(out_sel[28]),
		.A2(I28[2]),
		.B1(out_sel[29]),
		.B2(I29[2]),
		.Z(O14[2])
	);
	AO_CELL inst_15_2(
		.A1(out_sel[30]),
		.A2(I30[2]),
		.B1(out_sel[31]),
		.B2(I31[2]),
		.Z(O15[2])
	);
	AO_CELL inst_16_2(
		.A1(out_sel[32]),
		.A2(I32[2]),
		.B1(out_sel[33]),
		.B2(I33[2]),
		.Z(O16[2])
	);
	AO_CELL inst_17_2(
		.A1(out_sel[34]),
		.A2(I34[2]),
		.B1(out_sel[35]),
		.B2(I35[2]),
		.Z(O17[2])
	);
	AO_CELL inst_18_2(
		.A1(out_sel[36]),
		.A2(I36[2]),
		.B1(out_sel[37]),
		.B2(I37[2]),
		.Z(O18[2])
	);
	AO_CELL inst_19_2(
		.A1(out_sel[38]),
		.A2(I38[2]),
		.B1(out_sel[39]),
		.B2(I39[2]),
		.Z(O19[2])
	);
	AO_CELL inst_20_2(
		.A1(out_sel[40]),
		.A2(I40[2]),
		.B1(out_sel[41]),
		.B2(I41[2]),
		.Z(O20[2])
	);
	AO_CELL inst_21_2(
		.A1(out_sel[42]),
		.A2(I42[2]),
		.B1(out_sel[43]),
		.B2(I43[2]),
		.Z(O21[2])
	);
	AO_CELL inst_22_2(
		.A1(out_sel[44]),
		.A2(I44[2]),
		.B1(out_sel[45]),
		.B2(I45[2]),
		.Z(O22[2])
	);
	AN_CELL inst_and_2(
		.A1(out_sel[46]),
		.A2(I46[2]),
		.Z(O23[2])
	);
	AO_CELL inst_0_3(
		.A1(out_sel[0]),
		.A2(I0[3]),
		.B1(out_sel[1]),
		.B2(I1[3]),
		.Z(O0[3])
	);
	AO_CELL inst_1_3(
		.A1(out_sel[2]),
		.A2(I2[3]),
		.B1(out_sel[3]),
		.B2(I3[3]),
		.Z(O1[3])
	);
	AO_CELL inst_2_3(
		.A1(out_sel[4]),
		.A2(I4[3]),
		.B1(out_sel[5]),
		.B2(I5[3]),
		.Z(O2[3])
	);
	AO_CELL inst_3_3(
		.A1(out_sel[6]),
		.A2(I6[3]),
		.B1(out_sel[7]),
		.B2(I7[3]),
		.Z(O3[3])
	);
	AO_CELL inst_4_3(
		.A1(out_sel[8]),
		.A2(I8[3]),
		.B1(out_sel[9]),
		.B2(I9[3]),
		.Z(O4[3])
	);
	AO_CELL inst_5_3(
		.A1(out_sel[10]),
		.A2(I10[3]),
		.B1(out_sel[11]),
		.B2(I11[3]),
		.Z(O5[3])
	);
	AO_CELL inst_6_3(
		.A1(out_sel[12]),
		.A2(I12[3]),
		.B1(out_sel[13]),
		.B2(I13[3]),
		.Z(O6[3])
	);
	AO_CELL inst_7_3(
		.A1(out_sel[14]),
		.A2(I14[3]),
		.B1(out_sel[15]),
		.B2(I15[3]),
		.Z(O7[3])
	);
	AO_CELL inst_8_3(
		.A1(out_sel[16]),
		.A2(I16[3]),
		.B1(out_sel[17]),
		.B2(I17[3]),
		.Z(O8[3])
	);
	AO_CELL inst_9_3(
		.A1(out_sel[18]),
		.A2(I18[3]),
		.B1(out_sel[19]),
		.B2(I19[3]),
		.Z(O9[3])
	);
	AO_CELL inst_10_3(
		.A1(out_sel[20]),
		.A2(I20[3]),
		.B1(out_sel[21]),
		.B2(I21[3]),
		.Z(O10[3])
	);
	AO_CELL inst_11_3(
		.A1(out_sel[22]),
		.A2(I22[3]),
		.B1(out_sel[23]),
		.B2(I23[3]),
		.Z(O11[3])
	);
	AO_CELL inst_12_3(
		.A1(out_sel[24]),
		.A2(I24[3]),
		.B1(out_sel[25]),
		.B2(I25[3]),
		.Z(O12[3])
	);
	AO_CELL inst_13_3(
		.A1(out_sel[26]),
		.A2(I26[3]),
		.B1(out_sel[27]),
		.B2(I27[3]),
		.Z(O13[3])
	);
	AO_CELL inst_14_3(
		.A1(out_sel[28]),
		.A2(I28[3]),
		.B1(out_sel[29]),
		.B2(I29[3]),
		.Z(O14[3])
	);
	AO_CELL inst_15_3(
		.A1(out_sel[30]),
		.A2(I30[3]),
		.B1(out_sel[31]),
		.B2(I31[3]),
		.Z(O15[3])
	);
	AO_CELL inst_16_3(
		.A1(out_sel[32]),
		.A2(I32[3]),
		.B1(out_sel[33]),
		.B2(I33[3]),
		.Z(O16[3])
	);
	AO_CELL inst_17_3(
		.A1(out_sel[34]),
		.A2(I34[3]),
		.B1(out_sel[35]),
		.B2(I35[3]),
		.Z(O17[3])
	);
	AO_CELL inst_18_3(
		.A1(out_sel[36]),
		.A2(I36[3]),
		.B1(out_sel[37]),
		.B2(I37[3]),
		.Z(O18[3])
	);
	AO_CELL inst_19_3(
		.A1(out_sel[38]),
		.A2(I38[3]),
		.B1(out_sel[39]),
		.B2(I39[3]),
		.Z(O19[3])
	);
	AO_CELL inst_20_3(
		.A1(out_sel[40]),
		.A2(I40[3]),
		.B1(out_sel[41]),
		.B2(I41[3]),
		.Z(O20[3])
	);
	AO_CELL inst_21_3(
		.A1(out_sel[42]),
		.A2(I42[3]),
		.B1(out_sel[43]),
		.B2(I43[3]),
		.Z(O21[3])
	);
	AO_CELL inst_22_3(
		.A1(out_sel[44]),
		.A2(I44[3]),
		.B1(out_sel[45]),
		.B2(I45[3]),
		.Z(O22[3])
	);
	AN_CELL inst_and_3(
		.A1(out_sel[46]),
		.A2(I46[3]),
		.Z(O23[3])
	);
	AO_CELL inst_0_4(
		.A1(out_sel[0]),
		.A2(I0[4]),
		.B1(out_sel[1]),
		.B2(I1[4]),
		.Z(O0[4])
	);
	AO_CELL inst_1_4(
		.A1(out_sel[2]),
		.A2(I2[4]),
		.B1(out_sel[3]),
		.B2(I3[4]),
		.Z(O1[4])
	);
	AO_CELL inst_2_4(
		.A1(out_sel[4]),
		.A2(I4[4]),
		.B1(out_sel[5]),
		.B2(I5[4]),
		.Z(O2[4])
	);
	AO_CELL inst_3_4(
		.A1(out_sel[6]),
		.A2(I6[4]),
		.B1(out_sel[7]),
		.B2(I7[4]),
		.Z(O3[4])
	);
	AO_CELL inst_4_4(
		.A1(out_sel[8]),
		.A2(I8[4]),
		.B1(out_sel[9]),
		.B2(I9[4]),
		.Z(O4[4])
	);
	AO_CELL inst_5_4(
		.A1(out_sel[10]),
		.A2(I10[4]),
		.B1(out_sel[11]),
		.B2(I11[4]),
		.Z(O5[4])
	);
	AO_CELL inst_6_4(
		.A1(out_sel[12]),
		.A2(I12[4]),
		.B1(out_sel[13]),
		.B2(I13[4]),
		.Z(O6[4])
	);
	AO_CELL inst_7_4(
		.A1(out_sel[14]),
		.A2(I14[4]),
		.B1(out_sel[15]),
		.B2(I15[4]),
		.Z(O7[4])
	);
	AO_CELL inst_8_4(
		.A1(out_sel[16]),
		.A2(I16[4]),
		.B1(out_sel[17]),
		.B2(I17[4]),
		.Z(O8[4])
	);
	AO_CELL inst_9_4(
		.A1(out_sel[18]),
		.A2(I18[4]),
		.B1(out_sel[19]),
		.B2(I19[4]),
		.Z(O9[4])
	);
	AO_CELL inst_10_4(
		.A1(out_sel[20]),
		.A2(I20[4]),
		.B1(out_sel[21]),
		.B2(I21[4]),
		.Z(O10[4])
	);
	AO_CELL inst_11_4(
		.A1(out_sel[22]),
		.A2(I22[4]),
		.B1(out_sel[23]),
		.B2(I23[4]),
		.Z(O11[4])
	);
	AO_CELL inst_12_4(
		.A1(out_sel[24]),
		.A2(I24[4]),
		.B1(out_sel[25]),
		.B2(I25[4]),
		.Z(O12[4])
	);
	AO_CELL inst_13_4(
		.A1(out_sel[26]),
		.A2(I26[4]),
		.B1(out_sel[27]),
		.B2(I27[4]),
		.Z(O13[4])
	);
	AO_CELL inst_14_4(
		.A1(out_sel[28]),
		.A2(I28[4]),
		.B1(out_sel[29]),
		.B2(I29[4]),
		.Z(O14[4])
	);
	AO_CELL inst_15_4(
		.A1(out_sel[30]),
		.A2(I30[4]),
		.B1(out_sel[31]),
		.B2(I31[4]),
		.Z(O15[4])
	);
	AO_CELL inst_16_4(
		.A1(out_sel[32]),
		.A2(I32[4]),
		.B1(out_sel[33]),
		.B2(I33[4]),
		.Z(O16[4])
	);
	AO_CELL inst_17_4(
		.A1(out_sel[34]),
		.A2(I34[4]),
		.B1(out_sel[35]),
		.B2(I35[4]),
		.Z(O17[4])
	);
	AO_CELL inst_18_4(
		.A1(out_sel[36]),
		.A2(I36[4]),
		.B1(out_sel[37]),
		.B2(I37[4]),
		.Z(O18[4])
	);
	AO_CELL inst_19_4(
		.A1(out_sel[38]),
		.A2(I38[4]),
		.B1(out_sel[39]),
		.B2(I39[4]),
		.Z(O19[4])
	);
	AO_CELL inst_20_4(
		.A1(out_sel[40]),
		.A2(I40[4]),
		.B1(out_sel[41]),
		.B2(I41[4]),
		.Z(O20[4])
	);
	AO_CELL inst_21_4(
		.A1(out_sel[42]),
		.A2(I42[4]),
		.B1(out_sel[43]),
		.B2(I43[4]),
		.Z(O21[4])
	);
	AO_CELL inst_22_4(
		.A1(out_sel[44]),
		.A2(I44[4]),
		.B1(out_sel[45]),
		.B2(I45[4]),
		.Z(O22[4])
	);
	AN_CELL inst_and_4(
		.A1(out_sel[46]),
		.A2(I46[4]),
		.Z(O23[4])
	);
	AO_CELL inst_0_5(
		.A1(out_sel[0]),
		.A2(I0[5]),
		.B1(out_sel[1]),
		.B2(I1[5]),
		.Z(O0[5])
	);
	AO_CELL inst_1_5(
		.A1(out_sel[2]),
		.A2(I2[5]),
		.B1(out_sel[3]),
		.B2(I3[5]),
		.Z(O1[5])
	);
	AO_CELL inst_2_5(
		.A1(out_sel[4]),
		.A2(I4[5]),
		.B1(out_sel[5]),
		.B2(I5[5]),
		.Z(O2[5])
	);
	AO_CELL inst_3_5(
		.A1(out_sel[6]),
		.A2(I6[5]),
		.B1(out_sel[7]),
		.B2(I7[5]),
		.Z(O3[5])
	);
	AO_CELL inst_4_5(
		.A1(out_sel[8]),
		.A2(I8[5]),
		.B1(out_sel[9]),
		.B2(I9[5]),
		.Z(O4[5])
	);
	AO_CELL inst_5_5(
		.A1(out_sel[10]),
		.A2(I10[5]),
		.B1(out_sel[11]),
		.B2(I11[5]),
		.Z(O5[5])
	);
	AO_CELL inst_6_5(
		.A1(out_sel[12]),
		.A2(I12[5]),
		.B1(out_sel[13]),
		.B2(I13[5]),
		.Z(O6[5])
	);
	AO_CELL inst_7_5(
		.A1(out_sel[14]),
		.A2(I14[5]),
		.B1(out_sel[15]),
		.B2(I15[5]),
		.Z(O7[5])
	);
	AO_CELL inst_8_5(
		.A1(out_sel[16]),
		.A2(I16[5]),
		.B1(out_sel[17]),
		.B2(I17[5]),
		.Z(O8[5])
	);
	AO_CELL inst_9_5(
		.A1(out_sel[18]),
		.A2(I18[5]),
		.B1(out_sel[19]),
		.B2(I19[5]),
		.Z(O9[5])
	);
	AO_CELL inst_10_5(
		.A1(out_sel[20]),
		.A2(I20[5]),
		.B1(out_sel[21]),
		.B2(I21[5]),
		.Z(O10[5])
	);
	AO_CELL inst_11_5(
		.A1(out_sel[22]),
		.A2(I22[5]),
		.B1(out_sel[23]),
		.B2(I23[5]),
		.Z(O11[5])
	);
	AO_CELL inst_12_5(
		.A1(out_sel[24]),
		.A2(I24[5]),
		.B1(out_sel[25]),
		.B2(I25[5]),
		.Z(O12[5])
	);
	AO_CELL inst_13_5(
		.A1(out_sel[26]),
		.A2(I26[5]),
		.B1(out_sel[27]),
		.B2(I27[5]),
		.Z(O13[5])
	);
	AO_CELL inst_14_5(
		.A1(out_sel[28]),
		.A2(I28[5]),
		.B1(out_sel[29]),
		.B2(I29[5]),
		.Z(O14[5])
	);
	AO_CELL inst_15_5(
		.A1(out_sel[30]),
		.A2(I30[5]),
		.B1(out_sel[31]),
		.B2(I31[5]),
		.Z(O15[5])
	);
	AO_CELL inst_16_5(
		.A1(out_sel[32]),
		.A2(I32[5]),
		.B1(out_sel[33]),
		.B2(I33[5]),
		.Z(O16[5])
	);
	AO_CELL inst_17_5(
		.A1(out_sel[34]),
		.A2(I34[5]),
		.B1(out_sel[35]),
		.B2(I35[5]),
		.Z(O17[5])
	);
	AO_CELL inst_18_5(
		.A1(out_sel[36]),
		.A2(I36[5]),
		.B1(out_sel[37]),
		.B2(I37[5]),
		.Z(O18[5])
	);
	AO_CELL inst_19_5(
		.A1(out_sel[38]),
		.A2(I38[5]),
		.B1(out_sel[39]),
		.B2(I39[5]),
		.Z(O19[5])
	);
	AO_CELL inst_20_5(
		.A1(out_sel[40]),
		.A2(I40[5]),
		.B1(out_sel[41]),
		.B2(I41[5]),
		.Z(O20[5])
	);
	AO_CELL inst_21_5(
		.A1(out_sel[42]),
		.A2(I42[5]),
		.B1(out_sel[43]),
		.B2(I43[5]),
		.Z(O21[5])
	);
	AO_CELL inst_22_5(
		.A1(out_sel[44]),
		.A2(I44[5]),
		.B1(out_sel[45]),
		.B2(I45[5]),
		.Z(O22[5])
	);
	AN_CELL inst_and_5(
		.A1(out_sel[46]),
		.A2(I46[5]),
		.Z(O23[5])
	);
	AO_CELL inst_0_6(
		.A1(out_sel[0]),
		.A2(I0[6]),
		.B1(out_sel[1]),
		.B2(I1[6]),
		.Z(O0[6])
	);
	AO_CELL inst_1_6(
		.A1(out_sel[2]),
		.A2(I2[6]),
		.B1(out_sel[3]),
		.B2(I3[6]),
		.Z(O1[6])
	);
	AO_CELL inst_2_6(
		.A1(out_sel[4]),
		.A2(I4[6]),
		.B1(out_sel[5]),
		.B2(I5[6]),
		.Z(O2[6])
	);
	AO_CELL inst_3_6(
		.A1(out_sel[6]),
		.A2(I6[6]),
		.B1(out_sel[7]),
		.B2(I7[6]),
		.Z(O3[6])
	);
	AO_CELL inst_4_6(
		.A1(out_sel[8]),
		.A2(I8[6]),
		.B1(out_sel[9]),
		.B2(I9[6]),
		.Z(O4[6])
	);
	AO_CELL inst_5_6(
		.A1(out_sel[10]),
		.A2(I10[6]),
		.B1(out_sel[11]),
		.B2(I11[6]),
		.Z(O5[6])
	);
	AO_CELL inst_6_6(
		.A1(out_sel[12]),
		.A2(I12[6]),
		.B1(out_sel[13]),
		.B2(I13[6]),
		.Z(O6[6])
	);
	AO_CELL inst_7_6(
		.A1(out_sel[14]),
		.A2(I14[6]),
		.B1(out_sel[15]),
		.B2(I15[6]),
		.Z(O7[6])
	);
	AO_CELL inst_8_6(
		.A1(out_sel[16]),
		.A2(I16[6]),
		.B1(out_sel[17]),
		.B2(I17[6]),
		.Z(O8[6])
	);
	AO_CELL inst_9_6(
		.A1(out_sel[18]),
		.A2(I18[6]),
		.B1(out_sel[19]),
		.B2(I19[6]),
		.Z(O9[6])
	);
	AO_CELL inst_10_6(
		.A1(out_sel[20]),
		.A2(I20[6]),
		.B1(out_sel[21]),
		.B2(I21[6]),
		.Z(O10[6])
	);
	AO_CELL inst_11_6(
		.A1(out_sel[22]),
		.A2(I22[6]),
		.B1(out_sel[23]),
		.B2(I23[6]),
		.Z(O11[6])
	);
	AO_CELL inst_12_6(
		.A1(out_sel[24]),
		.A2(I24[6]),
		.B1(out_sel[25]),
		.B2(I25[6]),
		.Z(O12[6])
	);
	AO_CELL inst_13_6(
		.A1(out_sel[26]),
		.A2(I26[6]),
		.B1(out_sel[27]),
		.B2(I27[6]),
		.Z(O13[6])
	);
	AO_CELL inst_14_6(
		.A1(out_sel[28]),
		.A2(I28[6]),
		.B1(out_sel[29]),
		.B2(I29[6]),
		.Z(O14[6])
	);
	AO_CELL inst_15_6(
		.A1(out_sel[30]),
		.A2(I30[6]),
		.B1(out_sel[31]),
		.B2(I31[6]),
		.Z(O15[6])
	);
	AO_CELL inst_16_6(
		.A1(out_sel[32]),
		.A2(I32[6]),
		.B1(out_sel[33]),
		.B2(I33[6]),
		.Z(O16[6])
	);
	AO_CELL inst_17_6(
		.A1(out_sel[34]),
		.A2(I34[6]),
		.B1(out_sel[35]),
		.B2(I35[6]),
		.Z(O17[6])
	);
	AO_CELL inst_18_6(
		.A1(out_sel[36]),
		.A2(I36[6]),
		.B1(out_sel[37]),
		.B2(I37[6]),
		.Z(O18[6])
	);
	AO_CELL inst_19_6(
		.A1(out_sel[38]),
		.A2(I38[6]),
		.B1(out_sel[39]),
		.B2(I39[6]),
		.Z(O19[6])
	);
	AO_CELL inst_20_6(
		.A1(out_sel[40]),
		.A2(I40[6]),
		.B1(out_sel[41]),
		.B2(I41[6]),
		.Z(O20[6])
	);
	AO_CELL inst_21_6(
		.A1(out_sel[42]),
		.A2(I42[6]),
		.B1(out_sel[43]),
		.B2(I43[6]),
		.Z(O21[6])
	);
	AO_CELL inst_22_6(
		.A1(out_sel[44]),
		.A2(I44[6]),
		.B1(out_sel[45]),
		.B2(I45[6]),
		.Z(O22[6])
	);
	AN_CELL inst_and_6(
		.A1(out_sel[46]),
		.A2(I46[6]),
		.Z(O23[6])
	);
	AO_CELL inst_0_7(
		.A1(out_sel[0]),
		.A2(I0[7]),
		.B1(out_sel[1]),
		.B2(I1[7]),
		.Z(O0[7])
	);
	AO_CELL inst_1_7(
		.A1(out_sel[2]),
		.A2(I2[7]),
		.B1(out_sel[3]),
		.B2(I3[7]),
		.Z(O1[7])
	);
	AO_CELL inst_2_7(
		.A1(out_sel[4]),
		.A2(I4[7]),
		.B1(out_sel[5]),
		.B2(I5[7]),
		.Z(O2[7])
	);
	AO_CELL inst_3_7(
		.A1(out_sel[6]),
		.A2(I6[7]),
		.B1(out_sel[7]),
		.B2(I7[7]),
		.Z(O3[7])
	);
	AO_CELL inst_4_7(
		.A1(out_sel[8]),
		.A2(I8[7]),
		.B1(out_sel[9]),
		.B2(I9[7]),
		.Z(O4[7])
	);
	AO_CELL inst_5_7(
		.A1(out_sel[10]),
		.A2(I10[7]),
		.B1(out_sel[11]),
		.B2(I11[7]),
		.Z(O5[7])
	);
	AO_CELL inst_6_7(
		.A1(out_sel[12]),
		.A2(I12[7]),
		.B1(out_sel[13]),
		.B2(I13[7]),
		.Z(O6[7])
	);
	AO_CELL inst_7_7(
		.A1(out_sel[14]),
		.A2(I14[7]),
		.B1(out_sel[15]),
		.B2(I15[7]),
		.Z(O7[7])
	);
	AO_CELL inst_8_7(
		.A1(out_sel[16]),
		.A2(I16[7]),
		.B1(out_sel[17]),
		.B2(I17[7]),
		.Z(O8[7])
	);
	AO_CELL inst_9_7(
		.A1(out_sel[18]),
		.A2(I18[7]),
		.B1(out_sel[19]),
		.B2(I19[7]),
		.Z(O9[7])
	);
	AO_CELL inst_10_7(
		.A1(out_sel[20]),
		.A2(I20[7]),
		.B1(out_sel[21]),
		.B2(I21[7]),
		.Z(O10[7])
	);
	AO_CELL inst_11_7(
		.A1(out_sel[22]),
		.A2(I22[7]),
		.B1(out_sel[23]),
		.B2(I23[7]),
		.Z(O11[7])
	);
	AO_CELL inst_12_7(
		.A1(out_sel[24]),
		.A2(I24[7]),
		.B1(out_sel[25]),
		.B2(I25[7]),
		.Z(O12[7])
	);
	AO_CELL inst_13_7(
		.A1(out_sel[26]),
		.A2(I26[7]),
		.B1(out_sel[27]),
		.B2(I27[7]),
		.Z(O13[7])
	);
	AO_CELL inst_14_7(
		.A1(out_sel[28]),
		.A2(I28[7]),
		.B1(out_sel[29]),
		.B2(I29[7]),
		.Z(O14[7])
	);
	AO_CELL inst_15_7(
		.A1(out_sel[30]),
		.A2(I30[7]),
		.B1(out_sel[31]),
		.B2(I31[7]),
		.Z(O15[7])
	);
	AO_CELL inst_16_7(
		.A1(out_sel[32]),
		.A2(I32[7]),
		.B1(out_sel[33]),
		.B2(I33[7]),
		.Z(O16[7])
	);
	AO_CELL inst_17_7(
		.A1(out_sel[34]),
		.A2(I34[7]),
		.B1(out_sel[35]),
		.B2(I35[7]),
		.Z(O17[7])
	);
	AO_CELL inst_18_7(
		.A1(out_sel[36]),
		.A2(I36[7]),
		.B1(out_sel[37]),
		.B2(I37[7]),
		.Z(O18[7])
	);
	AO_CELL inst_19_7(
		.A1(out_sel[38]),
		.A2(I38[7]),
		.B1(out_sel[39]),
		.B2(I39[7]),
		.Z(O19[7])
	);
	AO_CELL inst_20_7(
		.A1(out_sel[40]),
		.A2(I40[7]),
		.B1(out_sel[41]),
		.B2(I41[7]),
		.Z(O20[7])
	);
	AO_CELL inst_21_7(
		.A1(out_sel[42]),
		.A2(I42[7]),
		.B1(out_sel[43]),
		.B2(I43[7]),
		.Z(O21[7])
	);
	AO_CELL inst_22_7(
		.A1(out_sel[44]),
		.A2(I44[7]),
		.B1(out_sel[45]),
		.B2(I45[7]),
		.Z(O22[7])
	);
	AN_CELL inst_and_7(
		.A1(out_sel[46]),
		.A2(I46[7]),
		.Z(O23[7])
	);
	AO_CELL inst_0_8(
		.A1(out_sel[0]),
		.A2(I0[8]),
		.B1(out_sel[1]),
		.B2(I1[8]),
		.Z(O0[8])
	);
	AO_CELL inst_1_8(
		.A1(out_sel[2]),
		.A2(I2[8]),
		.B1(out_sel[3]),
		.B2(I3[8]),
		.Z(O1[8])
	);
	AO_CELL inst_2_8(
		.A1(out_sel[4]),
		.A2(I4[8]),
		.B1(out_sel[5]),
		.B2(I5[8]),
		.Z(O2[8])
	);
	AO_CELL inst_3_8(
		.A1(out_sel[6]),
		.A2(I6[8]),
		.B1(out_sel[7]),
		.B2(I7[8]),
		.Z(O3[8])
	);
	AO_CELL inst_4_8(
		.A1(out_sel[8]),
		.A2(I8[8]),
		.B1(out_sel[9]),
		.B2(I9[8]),
		.Z(O4[8])
	);
	AO_CELL inst_5_8(
		.A1(out_sel[10]),
		.A2(I10[8]),
		.B1(out_sel[11]),
		.B2(I11[8]),
		.Z(O5[8])
	);
	AO_CELL inst_6_8(
		.A1(out_sel[12]),
		.A2(I12[8]),
		.B1(out_sel[13]),
		.B2(I13[8]),
		.Z(O6[8])
	);
	AO_CELL inst_7_8(
		.A1(out_sel[14]),
		.A2(I14[8]),
		.B1(out_sel[15]),
		.B2(I15[8]),
		.Z(O7[8])
	);
	AO_CELL inst_8_8(
		.A1(out_sel[16]),
		.A2(I16[8]),
		.B1(out_sel[17]),
		.B2(I17[8]),
		.Z(O8[8])
	);
	AO_CELL inst_9_8(
		.A1(out_sel[18]),
		.A2(I18[8]),
		.B1(out_sel[19]),
		.B2(I19[8]),
		.Z(O9[8])
	);
	AO_CELL inst_10_8(
		.A1(out_sel[20]),
		.A2(I20[8]),
		.B1(out_sel[21]),
		.B2(I21[8]),
		.Z(O10[8])
	);
	AO_CELL inst_11_8(
		.A1(out_sel[22]),
		.A2(I22[8]),
		.B1(out_sel[23]),
		.B2(I23[8]),
		.Z(O11[8])
	);
	AO_CELL inst_12_8(
		.A1(out_sel[24]),
		.A2(I24[8]),
		.B1(out_sel[25]),
		.B2(I25[8]),
		.Z(O12[8])
	);
	AO_CELL inst_13_8(
		.A1(out_sel[26]),
		.A2(I26[8]),
		.B1(out_sel[27]),
		.B2(I27[8]),
		.Z(O13[8])
	);
	AO_CELL inst_14_8(
		.A1(out_sel[28]),
		.A2(I28[8]),
		.B1(out_sel[29]),
		.B2(I29[8]),
		.Z(O14[8])
	);
	AO_CELL inst_15_8(
		.A1(out_sel[30]),
		.A2(I30[8]),
		.B1(out_sel[31]),
		.B2(I31[8]),
		.Z(O15[8])
	);
	AO_CELL inst_16_8(
		.A1(out_sel[32]),
		.A2(I32[8]),
		.B1(out_sel[33]),
		.B2(I33[8]),
		.Z(O16[8])
	);
	AO_CELL inst_17_8(
		.A1(out_sel[34]),
		.A2(I34[8]),
		.B1(out_sel[35]),
		.B2(I35[8]),
		.Z(O17[8])
	);
	AO_CELL inst_18_8(
		.A1(out_sel[36]),
		.A2(I36[8]),
		.B1(out_sel[37]),
		.B2(I37[8]),
		.Z(O18[8])
	);
	AO_CELL inst_19_8(
		.A1(out_sel[38]),
		.A2(I38[8]),
		.B1(out_sel[39]),
		.B2(I39[8]),
		.Z(O19[8])
	);
	AO_CELL inst_20_8(
		.A1(out_sel[40]),
		.A2(I40[8]),
		.B1(out_sel[41]),
		.B2(I41[8]),
		.Z(O20[8])
	);
	AO_CELL inst_21_8(
		.A1(out_sel[42]),
		.A2(I42[8]),
		.B1(out_sel[43]),
		.B2(I43[8]),
		.Z(O21[8])
	);
	AO_CELL inst_22_8(
		.A1(out_sel[44]),
		.A2(I44[8]),
		.B1(out_sel[45]),
		.B2(I45[8]),
		.Z(O22[8])
	);
	AN_CELL inst_and_8(
		.A1(out_sel[46]),
		.A2(I46[8]),
		.Z(O23[8])
	);
	AO_CELL inst_0_9(
		.A1(out_sel[0]),
		.A2(I0[9]),
		.B1(out_sel[1]),
		.B2(I1[9]),
		.Z(O0[9])
	);
	AO_CELL inst_1_9(
		.A1(out_sel[2]),
		.A2(I2[9]),
		.B1(out_sel[3]),
		.B2(I3[9]),
		.Z(O1[9])
	);
	AO_CELL inst_2_9(
		.A1(out_sel[4]),
		.A2(I4[9]),
		.B1(out_sel[5]),
		.B2(I5[9]),
		.Z(O2[9])
	);
	AO_CELL inst_3_9(
		.A1(out_sel[6]),
		.A2(I6[9]),
		.B1(out_sel[7]),
		.B2(I7[9]),
		.Z(O3[9])
	);
	AO_CELL inst_4_9(
		.A1(out_sel[8]),
		.A2(I8[9]),
		.B1(out_sel[9]),
		.B2(I9[9]),
		.Z(O4[9])
	);
	AO_CELL inst_5_9(
		.A1(out_sel[10]),
		.A2(I10[9]),
		.B1(out_sel[11]),
		.B2(I11[9]),
		.Z(O5[9])
	);
	AO_CELL inst_6_9(
		.A1(out_sel[12]),
		.A2(I12[9]),
		.B1(out_sel[13]),
		.B2(I13[9]),
		.Z(O6[9])
	);
	AO_CELL inst_7_9(
		.A1(out_sel[14]),
		.A2(I14[9]),
		.B1(out_sel[15]),
		.B2(I15[9]),
		.Z(O7[9])
	);
	AO_CELL inst_8_9(
		.A1(out_sel[16]),
		.A2(I16[9]),
		.B1(out_sel[17]),
		.B2(I17[9]),
		.Z(O8[9])
	);
	AO_CELL inst_9_9(
		.A1(out_sel[18]),
		.A2(I18[9]),
		.B1(out_sel[19]),
		.B2(I19[9]),
		.Z(O9[9])
	);
	AO_CELL inst_10_9(
		.A1(out_sel[20]),
		.A2(I20[9]),
		.B1(out_sel[21]),
		.B2(I21[9]),
		.Z(O10[9])
	);
	AO_CELL inst_11_9(
		.A1(out_sel[22]),
		.A2(I22[9]),
		.B1(out_sel[23]),
		.B2(I23[9]),
		.Z(O11[9])
	);
	AO_CELL inst_12_9(
		.A1(out_sel[24]),
		.A2(I24[9]),
		.B1(out_sel[25]),
		.B2(I25[9]),
		.Z(O12[9])
	);
	AO_CELL inst_13_9(
		.A1(out_sel[26]),
		.A2(I26[9]),
		.B1(out_sel[27]),
		.B2(I27[9]),
		.Z(O13[9])
	);
	AO_CELL inst_14_9(
		.A1(out_sel[28]),
		.A2(I28[9]),
		.B1(out_sel[29]),
		.B2(I29[9]),
		.Z(O14[9])
	);
	AO_CELL inst_15_9(
		.A1(out_sel[30]),
		.A2(I30[9]),
		.B1(out_sel[31]),
		.B2(I31[9]),
		.Z(O15[9])
	);
	AO_CELL inst_16_9(
		.A1(out_sel[32]),
		.A2(I32[9]),
		.B1(out_sel[33]),
		.B2(I33[9]),
		.Z(O16[9])
	);
	AO_CELL inst_17_9(
		.A1(out_sel[34]),
		.A2(I34[9]),
		.B1(out_sel[35]),
		.B2(I35[9]),
		.Z(O17[9])
	);
	AO_CELL inst_18_9(
		.A1(out_sel[36]),
		.A2(I36[9]),
		.B1(out_sel[37]),
		.B2(I37[9]),
		.Z(O18[9])
	);
	AO_CELL inst_19_9(
		.A1(out_sel[38]),
		.A2(I38[9]),
		.B1(out_sel[39]),
		.B2(I39[9]),
		.Z(O19[9])
	);
	AO_CELL inst_20_9(
		.A1(out_sel[40]),
		.A2(I40[9]),
		.B1(out_sel[41]),
		.B2(I41[9]),
		.Z(O20[9])
	);
	AO_CELL inst_21_9(
		.A1(out_sel[42]),
		.A2(I42[9]),
		.B1(out_sel[43]),
		.B2(I43[9]),
		.Z(O21[9])
	);
	AO_CELL inst_22_9(
		.A1(out_sel[44]),
		.A2(I44[9]),
		.B1(out_sel[45]),
		.B2(I45[9]),
		.Z(O22[9])
	);
	AN_CELL inst_and_9(
		.A1(out_sel[46]),
		.A2(I46[9]),
		.Z(O23[9])
	);
	AO_CELL inst_0_10(
		.A1(out_sel[0]),
		.A2(I0[10]),
		.B1(out_sel[1]),
		.B2(I1[10]),
		.Z(O0[10])
	);
	AO_CELL inst_1_10(
		.A1(out_sel[2]),
		.A2(I2[10]),
		.B1(out_sel[3]),
		.B2(I3[10]),
		.Z(O1[10])
	);
	AO_CELL inst_2_10(
		.A1(out_sel[4]),
		.A2(I4[10]),
		.B1(out_sel[5]),
		.B2(I5[10]),
		.Z(O2[10])
	);
	AO_CELL inst_3_10(
		.A1(out_sel[6]),
		.A2(I6[10]),
		.B1(out_sel[7]),
		.B2(I7[10]),
		.Z(O3[10])
	);
	AO_CELL inst_4_10(
		.A1(out_sel[8]),
		.A2(I8[10]),
		.B1(out_sel[9]),
		.B2(I9[10]),
		.Z(O4[10])
	);
	AO_CELL inst_5_10(
		.A1(out_sel[10]),
		.A2(I10[10]),
		.B1(out_sel[11]),
		.B2(I11[10]),
		.Z(O5[10])
	);
	AO_CELL inst_6_10(
		.A1(out_sel[12]),
		.A2(I12[10]),
		.B1(out_sel[13]),
		.B2(I13[10]),
		.Z(O6[10])
	);
	AO_CELL inst_7_10(
		.A1(out_sel[14]),
		.A2(I14[10]),
		.B1(out_sel[15]),
		.B2(I15[10]),
		.Z(O7[10])
	);
	AO_CELL inst_8_10(
		.A1(out_sel[16]),
		.A2(I16[10]),
		.B1(out_sel[17]),
		.B2(I17[10]),
		.Z(O8[10])
	);
	AO_CELL inst_9_10(
		.A1(out_sel[18]),
		.A2(I18[10]),
		.B1(out_sel[19]),
		.B2(I19[10]),
		.Z(O9[10])
	);
	AO_CELL inst_10_10(
		.A1(out_sel[20]),
		.A2(I20[10]),
		.B1(out_sel[21]),
		.B2(I21[10]),
		.Z(O10[10])
	);
	AO_CELL inst_11_10(
		.A1(out_sel[22]),
		.A2(I22[10]),
		.B1(out_sel[23]),
		.B2(I23[10]),
		.Z(O11[10])
	);
	AO_CELL inst_12_10(
		.A1(out_sel[24]),
		.A2(I24[10]),
		.B1(out_sel[25]),
		.B2(I25[10]),
		.Z(O12[10])
	);
	AO_CELL inst_13_10(
		.A1(out_sel[26]),
		.A2(I26[10]),
		.B1(out_sel[27]),
		.B2(I27[10]),
		.Z(O13[10])
	);
	AO_CELL inst_14_10(
		.A1(out_sel[28]),
		.A2(I28[10]),
		.B1(out_sel[29]),
		.B2(I29[10]),
		.Z(O14[10])
	);
	AO_CELL inst_15_10(
		.A1(out_sel[30]),
		.A2(I30[10]),
		.B1(out_sel[31]),
		.B2(I31[10]),
		.Z(O15[10])
	);
	AO_CELL inst_16_10(
		.A1(out_sel[32]),
		.A2(I32[10]),
		.B1(out_sel[33]),
		.B2(I33[10]),
		.Z(O16[10])
	);
	AO_CELL inst_17_10(
		.A1(out_sel[34]),
		.A2(I34[10]),
		.B1(out_sel[35]),
		.B2(I35[10]),
		.Z(O17[10])
	);
	AO_CELL inst_18_10(
		.A1(out_sel[36]),
		.A2(I36[10]),
		.B1(out_sel[37]),
		.B2(I37[10]),
		.Z(O18[10])
	);
	AO_CELL inst_19_10(
		.A1(out_sel[38]),
		.A2(I38[10]),
		.B1(out_sel[39]),
		.B2(I39[10]),
		.Z(O19[10])
	);
	AO_CELL inst_20_10(
		.A1(out_sel[40]),
		.A2(I40[10]),
		.B1(out_sel[41]),
		.B2(I41[10]),
		.Z(O20[10])
	);
	AO_CELL inst_21_10(
		.A1(out_sel[42]),
		.A2(I42[10]),
		.B1(out_sel[43]),
		.B2(I43[10]),
		.Z(O21[10])
	);
	AO_CELL inst_22_10(
		.A1(out_sel[44]),
		.A2(I44[10]),
		.B1(out_sel[45]),
		.B2(I45[10]),
		.Z(O22[10])
	);
	AN_CELL inst_and_10(
		.A1(out_sel[46]),
		.A2(I46[10]),
		.Z(O23[10])
	);
	AO_CELL inst_0_11(
		.A1(out_sel[0]),
		.A2(I0[11]),
		.B1(out_sel[1]),
		.B2(I1[11]),
		.Z(O0[11])
	);
	AO_CELL inst_1_11(
		.A1(out_sel[2]),
		.A2(I2[11]),
		.B1(out_sel[3]),
		.B2(I3[11]),
		.Z(O1[11])
	);
	AO_CELL inst_2_11(
		.A1(out_sel[4]),
		.A2(I4[11]),
		.B1(out_sel[5]),
		.B2(I5[11]),
		.Z(O2[11])
	);
	AO_CELL inst_3_11(
		.A1(out_sel[6]),
		.A2(I6[11]),
		.B1(out_sel[7]),
		.B2(I7[11]),
		.Z(O3[11])
	);
	AO_CELL inst_4_11(
		.A1(out_sel[8]),
		.A2(I8[11]),
		.B1(out_sel[9]),
		.B2(I9[11]),
		.Z(O4[11])
	);
	AO_CELL inst_5_11(
		.A1(out_sel[10]),
		.A2(I10[11]),
		.B1(out_sel[11]),
		.B2(I11[11]),
		.Z(O5[11])
	);
	AO_CELL inst_6_11(
		.A1(out_sel[12]),
		.A2(I12[11]),
		.B1(out_sel[13]),
		.B2(I13[11]),
		.Z(O6[11])
	);
	AO_CELL inst_7_11(
		.A1(out_sel[14]),
		.A2(I14[11]),
		.B1(out_sel[15]),
		.B2(I15[11]),
		.Z(O7[11])
	);
	AO_CELL inst_8_11(
		.A1(out_sel[16]),
		.A2(I16[11]),
		.B1(out_sel[17]),
		.B2(I17[11]),
		.Z(O8[11])
	);
	AO_CELL inst_9_11(
		.A1(out_sel[18]),
		.A2(I18[11]),
		.B1(out_sel[19]),
		.B2(I19[11]),
		.Z(O9[11])
	);
	AO_CELL inst_10_11(
		.A1(out_sel[20]),
		.A2(I20[11]),
		.B1(out_sel[21]),
		.B2(I21[11]),
		.Z(O10[11])
	);
	AO_CELL inst_11_11(
		.A1(out_sel[22]),
		.A2(I22[11]),
		.B1(out_sel[23]),
		.B2(I23[11]),
		.Z(O11[11])
	);
	AO_CELL inst_12_11(
		.A1(out_sel[24]),
		.A2(I24[11]),
		.B1(out_sel[25]),
		.B2(I25[11]),
		.Z(O12[11])
	);
	AO_CELL inst_13_11(
		.A1(out_sel[26]),
		.A2(I26[11]),
		.B1(out_sel[27]),
		.B2(I27[11]),
		.Z(O13[11])
	);
	AO_CELL inst_14_11(
		.A1(out_sel[28]),
		.A2(I28[11]),
		.B1(out_sel[29]),
		.B2(I29[11]),
		.Z(O14[11])
	);
	AO_CELL inst_15_11(
		.A1(out_sel[30]),
		.A2(I30[11]),
		.B1(out_sel[31]),
		.B2(I31[11]),
		.Z(O15[11])
	);
	AO_CELL inst_16_11(
		.A1(out_sel[32]),
		.A2(I32[11]),
		.B1(out_sel[33]),
		.B2(I33[11]),
		.Z(O16[11])
	);
	AO_CELL inst_17_11(
		.A1(out_sel[34]),
		.A2(I34[11]),
		.B1(out_sel[35]),
		.B2(I35[11]),
		.Z(O17[11])
	);
	AO_CELL inst_18_11(
		.A1(out_sel[36]),
		.A2(I36[11]),
		.B1(out_sel[37]),
		.B2(I37[11]),
		.Z(O18[11])
	);
	AO_CELL inst_19_11(
		.A1(out_sel[38]),
		.A2(I38[11]),
		.B1(out_sel[39]),
		.B2(I39[11]),
		.Z(O19[11])
	);
	AO_CELL inst_20_11(
		.A1(out_sel[40]),
		.A2(I40[11]),
		.B1(out_sel[41]),
		.B2(I41[11]),
		.Z(O20[11])
	);
	AO_CELL inst_21_11(
		.A1(out_sel[42]),
		.A2(I42[11]),
		.B1(out_sel[43]),
		.B2(I43[11]),
		.Z(O21[11])
	);
	AO_CELL inst_22_11(
		.A1(out_sel[44]),
		.A2(I44[11]),
		.B1(out_sel[45]),
		.B2(I45[11]),
		.Z(O22[11])
	);
	AN_CELL inst_and_11(
		.A1(out_sel[46]),
		.A2(I46[11]),
		.Z(O23[11])
	);
	AO_CELL inst_0_12(
		.A1(out_sel[0]),
		.A2(I0[12]),
		.B1(out_sel[1]),
		.B2(I1[12]),
		.Z(O0[12])
	);
	AO_CELL inst_1_12(
		.A1(out_sel[2]),
		.A2(I2[12]),
		.B1(out_sel[3]),
		.B2(I3[12]),
		.Z(O1[12])
	);
	AO_CELL inst_2_12(
		.A1(out_sel[4]),
		.A2(I4[12]),
		.B1(out_sel[5]),
		.B2(I5[12]),
		.Z(O2[12])
	);
	AO_CELL inst_3_12(
		.A1(out_sel[6]),
		.A2(I6[12]),
		.B1(out_sel[7]),
		.B2(I7[12]),
		.Z(O3[12])
	);
	AO_CELL inst_4_12(
		.A1(out_sel[8]),
		.A2(I8[12]),
		.B1(out_sel[9]),
		.B2(I9[12]),
		.Z(O4[12])
	);
	AO_CELL inst_5_12(
		.A1(out_sel[10]),
		.A2(I10[12]),
		.B1(out_sel[11]),
		.B2(I11[12]),
		.Z(O5[12])
	);
	AO_CELL inst_6_12(
		.A1(out_sel[12]),
		.A2(I12[12]),
		.B1(out_sel[13]),
		.B2(I13[12]),
		.Z(O6[12])
	);
	AO_CELL inst_7_12(
		.A1(out_sel[14]),
		.A2(I14[12]),
		.B1(out_sel[15]),
		.B2(I15[12]),
		.Z(O7[12])
	);
	AO_CELL inst_8_12(
		.A1(out_sel[16]),
		.A2(I16[12]),
		.B1(out_sel[17]),
		.B2(I17[12]),
		.Z(O8[12])
	);
	AO_CELL inst_9_12(
		.A1(out_sel[18]),
		.A2(I18[12]),
		.B1(out_sel[19]),
		.B2(I19[12]),
		.Z(O9[12])
	);
	AO_CELL inst_10_12(
		.A1(out_sel[20]),
		.A2(I20[12]),
		.B1(out_sel[21]),
		.B2(I21[12]),
		.Z(O10[12])
	);
	AO_CELL inst_11_12(
		.A1(out_sel[22]),
		.A2(I22[12]),
		.B1(out_sel[23]),
		.B2(I23[12]),
		.Z(O11[12])
	);
	AO_CELL inst_12_12(
		.A1(out_sel[24]),
		.A2(I24[12]),
		.B1(out_sel[25]),
		.B2(I25[12]),
		.Z(O12[12])
	);
	AO_CELL inst_13_12(
		.A1(out_sel[26]),
		.A2(I26[12]),
		.B1(out_sel[27]),
		.B2(I27[12]),
		.Z(O13[12])
	);
	AO_CELL inst_14_12(
		.A1(out_sel[28]),
		.A2(I28[12]),
		.B1(out_sel[29]),
		.B2(I29[12]),
		.Z(O14[12])
	);
	AO_CELL inst_15_12(
		.A1(out_sel[30]),
		.A2(I30[12]),
		.B1(out_sel[31]),
		.B2(I31[12]),
		.Z(O15[12])
	);
	AO_CELL inst_16_12(
		.A1(out_sel[32]),
		.A2(I32[12]),
		.B1(out_sel[33]),
		.B2(I33[12]),
		.Z(O16[12])
	);
	AO_CELL inst_17_12(
		.A1(out_sel[34]),
		.A2(I34[12]),
		.B1(out_sel[35]),
		.B2(I35[12]),
		.Z(O17[12])
	);
	AO_CELL inst_18_12(
		.A1(out_sel[36]),
		.A2(I36[12]),
		.B1(out_sel[37]),
		.B2(I37[12]),
		.Z(O18[12])
	);
	AO_CELL inst_19_12(
		.A1(out_sel[38]),
		.A2(I38[12]),
		.B1(out_sel[39]),
		.B2(I39[12]),
		.Z(O19[12])
	);
	AO_CELL inst_20_12(
		.A1(out_sel[40]),
		.A2(I40[12]),
		.B1(out_sel[41]),
		.B2(I41[12]),
		.Z(O20[12])
	);
	AO_CELL inst_21_12(
		.A1(out_sel[42]),
		.A2(I42[12]),
		.B1(out_sel[43]),
		.B2(I43[12]),
		.Z(O21[12])
	);
	AO_CELL inst_22_12(
		.A1(out_sel[44]),
		.A2(I44[12]),
		.B1(out_sel[45]),
		.B2(I45[12]),
		.Z(O22[12])
	);
	AN_CELL inst_and_12(
		.A1(out_sel[46]),
		.A2(I46[12]),
		.Z(O23[12])
	);
	AO_CELL inst_0_13(
		.A1(out_sel[0]),
		.A2(I0[13]),
		.B1(out_sel[1]),
		.B2(I1[13]),
		.Z(O0[13])
	);
	AO_CELL inst_1_13(
		.A1(out_sel[2]),
		.A2(I2[13]),
		.B1(out_sel[3]),
		.B2(I3[13]),
		.Z(O1[13])
	);
	AO_CELL inst_2_13(
		.A1(out_sel[4]),
		.A2(I4[13]),
		.B1(out_sel[5]),
		.B2(I5[13]),
		.Z(O2[13])
	);
	AO_CELL inst_3_13(
		.A1(out_sel[6]),
		.A2(I6[13]),
		.B1(out_sel[7]),
		.B2(I7[13]),
		.Z(O3[13])
	);
	AO_CELL inst_4_13(
		.A1(out_sel[8]),
		.A2(I8[13]),
		.B1(out_sel[9]),
		.B2(I9[13]),
		.Z(O4[13])
	);
	AO_CELL inst_5_13(
		.A1(out_sel[10]),
		.A2(I10[13]),
		.B1(out_sel[11]),
		.B2(I11[13]),
		.Z(O5[13])
	);
	AO_CELL inst_6_13(
		.A1(out_sel[12]),
		.A2(I12[13]),
		.B1(out_sel[13]),
		.B2(I13[13]),
		.Z(O6[13])
	);
	AO_CELL inst_7_13(
		.A1(out_sel[14]),
		.A2(I14[13]),
		.B1(out_sel[15]),
		.B2(I15[13]),
		.Z(O7[13])
	);
	AO_CELL inst_8_13(
		.A1(out_sel[16]),
		.A2(I16[13]),
		.B1(out_sel[17]),
		.B2(I17[13]),
		.Z(O8[13])
	);
	AO_CELL inst_9_13(
		.A1(out_sel[18]),
		.A2(I18[13]),
		.B1(out_sel[19]),
		.B2(I19[13]),
		.Z(O9[13])
	);
	AO_CELL inst_10_13(
		.A1(out_sel[20]),
		.A2(I20[13]),
		.B1(out_sel[21]),
		.B2(I21[13]),
		.Z(O10[13])
	);
	AO_CELL inst_11_13(
		.A1(out_sel[22]),
		.A2(I22[13]),
		.B1(out_sel[23]),
		.B2(I23[13]),
		.Z(O11[13])
	);
	AO_CELL inst_12_13(
		.A1(out_sel[24]),
		.A2(I24[13]),
		.B1(out_sel[25]),
		.B2(I25[13]),
		.Z(O12[13])
	);
	AO_CELL inst_13_13(
		.A1(out_sel[26]),
		.A2(I26[13]),
		.B1(out_sel[27]),
		.B2(I27[13]),
		.Z(O13[13])
	);
	AO_CELL inst_14_13(
		.A1(out_sel[28]),
		.A2(I28[13]),
		.B1(out_sel[29]),
		.B2(I29[13]),
		.Z(O14[13])
	);
	AO_CELL inst_15_13(
		.A1(out_sel[30]),
		.A2(I30[13]),
		.B1(out_sel[31]),
		.B2(I31[13]),
		.Z(O15[13])
	);
	AO_CELL inst_16_13(
		.A1(out_sel[32]),
		.A2(I32[13]),
		.B1(out_sel[33]),
		.B2(I33[13]),
		.Z(O16[13])
	);
	AO_CELL inst_17_13(
		.A1(out_sel[34]),
		.A2(I34[13]),
		.B1(out_sel[35]),
		.B2(I35[13]),
		.Z(O17[13])
	);
	AO_CELL inst_18_13(
		.A1(out_sel[36]),
		.A2(I36[13]),
		.B1(out_sel[37]),
		.B2(I37[13]),
		.Z(O18[13])
	);
	AO_CELL inst_19_13(
		.A1(out_sel[38]),
		.A2(I38[13]),
		.B1(out_sel[39]),
		.B2(I39[13]),
		.Z(O19[13])
	);
	AO_CELL inst_20_13(
		.A1(out_sel[40]),
		.A2(I40[13]),
		.B1(out_sel[41]),
		.B2(I41[13]),
		.Z(O20[13])
	);
	AO_CELL inst_21_13(
		.A1(out_sel[42]),
		.A2(I42[13]),
		.B1(out_sel[43]),
		.B2(I43[13]),
		.Z(O21[13])
	);
	AO_CELL inst_22_13(
		.A1(out_sel[44]),
		.A2(I44[13]),
		.B1(out_sel[45]),
		.B2(I45[13]),
		.Z(O22[13])
	);
	AN_CELL inst_and_13(
		.A1(out_sel[46]),
		.A2(I46[13]),
		.Z(O23[13])
	);
	AO_CELL inst_0_14(
		.A1(out_sel[0]),
		.A2(I0[14]),
		.B1(out_sel[1]),
		.B2(I1[14]),
		.Z(O0[14])
	);
	AO_CELL inst_1_14(
		.A1(out_sel[2]),
		.A2(I2[14]),
		.B1(out_sel[3]),
		.B2(I3[14]),
		.Z(O1[14])
	);
	AO_CELL inst_2_14(
		.A1(out_sel[4]),
		.A2(I4[14]),
		.B1(out_sel[5]),
		.B2(I5[14]),
		.Z(O2[14])
	);
	AO_CELL inst_3_14(
		.A1(out_sel[6]),
		.A2(I6[14]),
		.B1(out_sel[7]),
		.B2(I7[14]),
		.Z(O3[14])
	);
	AO_CELL inst_4_14(
		.A1(out_sel[8]),
		.A2(I8[14]),
		.B1(out_sel[9]),
		.B2(I9[14]),
		.Z(O4[14])
	);
	AO_CELL inst_5_14(
		.A1(out_sel[10]),
		.A2(I10[14]),
		.B1(out_sel[11]),
		.B2(I11[14]),
		.Z(O5[14])
	);
	AO_CELL inst_6_14(
		.A1(out_sel[12]),
		.A2(I12[14]),
		.B1(out_sel[13]),
		.B2(I13[14]),
		.Z(O6[14])
	);
	AO_CELL inst_7_14(
		.A1(out_sel[14]),
		.A2(I14[14]),
		.B1(out_sel[15]),
		.B2(I15[14]),
		.Z(O7[14])
	);
	AO_CELL inst_8_14(
		.A1(out_sel[16]),
		.A2(I16[14]),
		.B1(out_sel[17]),
		.B2(I17[14]),
		.Z(O8[14])
	);
	AO_CELL inst_9_14(
		.A1(out_sel[18]),
		.A2(I18[14]),
		.B1(out_sel[19]),
		.B2(I19[14]),
		.Z(O9[14])
	);
	AO_CELL inst_10_14(
		.A1(out_sel[20]),
		.A2(I20[14]),
		.B1(out_sel[21]),
		.B2(I21[14]),
		.Z(O10[14])
	);
	AO_CELL inst_11_14(
		.A1(out_sel[22]),
		.A2(I22[14]),
		.B1(out_sel[23]),
		.B2(I23[14]),
		.Z(O11[14])
	);
	AO_CELL inst_12_14(
		.A1(out_sel[24]),
		.A2(I24[14]),
		.B1(out_sel[25]),
		.B2(I25[14]),
		.Z(O12[14])
	);
	AO_CELL inst_13_14(
		.A1(out_sel[26]),
		.A2(I26[14]),
		.B1(out_sel[27]),
		.B2(I27[14]),
		.Z(O13[14])
	);
	AO_CELL inst_14_14(
		.A1(out_sel[28]),
		.A2(I28[14]),
		.B1(out_sel[29]),
		.B2(I29[14]),
		.Z(O14[14])
	);
	AO_CELL inst_15_14(
		.A1(out_sel[30]),
		.A2(I30[14]),
		.B1(out_sel[31]),
		.B2(I31[14]),
		.Z(O15[14])
	);
	AO_CELL inst_16_14(
		.A1(out_sel[32]),
		.A2(I32[14]),
		.B1(out_sel[33]),
		.B2(I33[14]),
		.Z(O16[14])
	);
	AO_CELL inst_17_14(
		.A1(out_sel[34]),
		.A2(I34[14]),
		.B1(out_sel[35]),
		.B2(I35[14]),
		.Z(O17[14])
	);
	AO_CELL inst_18_14(
		.A1(out_sel[36]),
		.A2(I36[14]),
		.B1(out_sel[37]),
		.B2(I37[14]),
		.Z(O18[14])
	);
	AO_CELL inst_19_14(
		.A1(out_sel[38]),
		.A2(I38[14]),
		.B1(out_sel[39]),
		.B2(I39[14]),
		.Z(O19[14])
	);
	AO_CELL inst_20_14(
		.A1(out_sel[40]),
		.A2(I40[14]),
		.B1(out_sel[41]),
		.B2(I41[14]),
		.Z(O20[14])
	);
	AO_CELL inst_21_14(
		.A1(out_sel[42]),
		.A2(I42[14]),
		.B1(out_sel[43]),
		.B2(I43[14]),
		.Z(O21[14])
	);
	AO_CELL inst_22_14(
		.A1(out_sel[44]),
		.A2(I44[14]),
		.B1(out_sel[45]),
		.B2(I45[14]),
		.Z(O22[14])
	);
	AN_CELL inst_and_14(
		.A1(out_sel[46]),
		.A2(I46[14]),
		.Z(O23[14])
	);
	AO_CELL inst_0_15(
		.A1(out_sel[0]),
		.A2(I0[15]),
		.B1(out_sel[1]),
		.B2(I1[15]),
		.Z(O0[15])
	);
	AO_CELL inst_1_15(
		.A1(out_sel[2]),
		.A2(I2[15]),
		.B1(out_sel[3]),
		.B2(I3[15]),
		.Z(O1[15])
	);
	AO_CELL inst_2_15(
		.A1(out_sel[4]),
		.A2(I4[15]),
		.B1(out_sel[5]),
		.B2(I5[15]),
		.Z(O2[15])
	);
	AO_CELL inst_3_15(
		.A1(out_sel[6]),
		.A2(I6[15]),
		.B1(out_sel[7]),
		.B2(I7[15]),
		.Z(O3[15])
	);
	AO_CELL inst_4_15(
		.A1(out_sel[8]),
		.A2(I8[15]),
		.B1(out_sel[9]),
		.B2(I9[15]),
		.Z(O4[15])
	);
	AO_CELL inst_5_15(
		.A1(out_sel[10]),
		.A2(I10[15]),
		.B1(out_sel[11]),
		.B2(I11[15]),
		.Z(O5[15])
	);
	AO_CELL inst_6_15(
		.A1(out_sel[12]),
		.A2(I12[15]),
		.B1(out_sel[13]),
		.B2(I13[15]),
		.Z(O6[15])
	);
	AO_CELL inst_7_15(
		.A1(out_sel[14]),
		.A2(I14[15]),
		.B1(out_sel[15]),
		.B2(I15[15]),
		.Z(O7[15])
	);
	AO_CELL inst_8_15(
		.A1(out_sel[16]),
		.A2(I16[15]),
		.B1(out_sel[17]),
		.B2(I17[15]),
		.Z(O8[15])
	);
	AO_CELL inst_9_15(
		.A1(out_sel[18]),
		.A2(I18[15]),
		.B1(out_sel[19]),
		.B2(I19[15]),
		.Z(O9[15])
	);
	AO_CELL inst_10_15(
		.A1(out_sel[20]),
		.A2(I20[15]),
		.B1(out_sel[21]),
		.B2(I21[15]),
		.Z(O10[15])
	);
	AO_CELL inst_11_15(
		.A1(out_sel[22]),
		.A2(I22[15]),
		.B1(out_sel[23]),
		.B2(I23[15]),
		.Z(O11[15])
	);
	AO_CELL inst_12_15(
		.A1(out_sel[24]),
		.A2(I24[15]),
		.B1(out_sel[25]),
		.B2(I25[15]),
		.Z(O12[15])
	);
	AO_CELL inst_13_15(
		.A1(out_sel[26]),
		.A2(I26[15]),
		.B1(out_sel[27]),
		.B2(I27[15]),
		.Z(O13[15])
	);
	AO_CELL inst_14_15(
		.A1(out_sel[28]),
		.A2(I28[15]),
		.B1(out_sel[29]),
		.B2(I29[15]),
		.Z(O14[15])
	);
	AO_CELL inst_15_15(
		.A1(out_sel[30]),
		.A2(I30[15]),
		.B1(out_sel[31]),
		.B2(I31[15]),
		.Z(O15[15])
	);
	AO_CELL inst_16_15(
		.A1(out_sel[32]),
		.A2(I32[15]),
		.B1(out_sel[33]),
		.B2(I33[15]),
		.Z(O16[15])
	);
	AO_CELL inst_17_15(
		.A1(out_sel[34]),
		.A2(I34[15]),
		.B1(out_sel[35]),
		.B2(I35[15]),
		.Z(O17[15])
	);
	AO_CELL inst_18_15(
		.A1(out_sel[36]),
		.A2(I36[15]),
		.B1(out_sel[37]),
		.B2(I37[15]),
		.Z(O18[15])
	);
	AO_CELL inst_19_15(
		.A1(out_sel[38]),
		.A2(I38[15]),
		.B1(out_sel[39]),
		.B2(I39[15]),
		.Z(O19[15])
	);
	AO_CELL inst_20_15(
		.A1(out_sel[40]),
		.A2(I40[15]),
		.B1(out_sel[41]),
		.B2(I41[15]),
		.Z(O20[15])
	);
	AO_CELL inst_21_15(
		.A1(out_sel[42]),
		.A2(I42[15]),
		.B1(out_sel[43]),
		.B2(I43[15]),
		.Z(O21[15])
	);
	AO_CELL inst_22_15(
		.A1(out_sel[44]),
		.A2(I44[15]),
		.B1(out_sel[45]),
		.B2(I45[15]),
		.Z(O22[15])
	);
	AN_CELL inst_and_15(
		.A1(out_sel[46]),
		.A2(I46[15]),
		.Z(O23[15])
	);
	AO_CELL inst_0_16(
		.A1(out_sel[0]),
		.A2(I0[16]),
		.B1(out_sel[1]),
		.B2(I1[16]),
		.Z(O0[16])
	);
	AO_CELL inst_1_16(
		.A1(out_sel[2]),
		.A2(I2[16]),
		.B1(out_sel[3]),
		.B2(I3[16]),
		.Z(O1[16])
	);
	AO_CELL inst_2_16(
		.A1(out_sel[4]),
		.A2(I4[16]),
		.B1(out_sel[5]),
		.B2(I5[16]),
		.Z(O2[16])
	);
	AO_CELL inst_3_16(
		.A1(out_sel[6]),
		.A2(I6[16]),
		.B1(out_sel[7]),
		.B2(I7[16]),
		.Z(O3[16])
	);
	AO_CELL inst_4_16(
		.A1(out_sel[8]),
		.A2(I8[16]),
		.B1(out_sel[9]),
		.B2(I9[16]),
		.Z(O4[16])
	);
	AO_CELL inst_5_16(
		.A1(out_sel[10]),
		.A2(I10[16]),
		.B1(out_sel[11]),
		.B2(I11[16]),
		.Z(O5[16])
	);
	AO_CELL inst_6_16(
		.A1(out_sel[12]),
		.A2(I12[16]),
		.B1(out_sel[13]),
		.B2(I13[16]),
		.Z(O6[16])
	);
	AO_CELL inst_7_16(
		.A1(out_sel[14]),
		.A2(I14[16]),
		.B1(out_sel[15]),
		.B2(I15[16]),
		.Z(O7[16])
	);
	AO_CELL inst_8_16(
		.A1(out_sel[16]),
		.A2(I16[16]),
		.B1(out_sel[17]),
		.B2(I17[16]),
		.Z(O8[16])
	);
	AO_CELL inst_9_16(
		.A1(out_sel[18]),
		.A2(I18[16]),
		.B1(out_sel[19]),
		.B2(I19[16]),
		.Z(O9[16])
	);
	AO_CELL inst_10_16(
		.A1(out_sel[20]),
		.A2(I20[16]),
		.B1(out_sel[21]),
		.B2(I21[16]),
		.Z(O10[16])
	);
	AO_CELL inst_11_16(
		.A1(out_sel[22]),
		.A2(I22[16]),
		.B1(out_sel[23]),
		.B2(I23[16]),
		.Z(O11[16])
	);
	AO_CELL inst_12_16(
		.A1(out_sel[24]),
		.A2(I24[16]),
		.B1(out_sel[25]),
		.B2(I25[16]),
		.Z(O12[16])
	);
	AO_CELL inst_13_16(
		.A1(out_sel[26]),
		.A2(I26[16]),
		.B1(out_sel[27]),
		.B2(I27[16]),
		.Z(O13[16])
	);
	AO_CELL inst_14_16(
		.A1(out_sel[28]),
		.A2(I28[16]),
		.B1(out_sel[29]),
		.B2(I29[16]),
		.Z(O14[16])
	);
	AO_CELL inst_15_16(
		.A1(out_sel[30]),
		.A2(I30[16]),
		.B1(out_sel[31]),
		.B2(I31[16]),
		.Z(O15[16])
	);
	AO_CELL inst_16_16(
		.A1(out_sel[32]),
		.A2(I32[16]),
		.B1(out_sel[33]),
		.B2(I33[16]),
		.Z(O16[16])
	);
	AO_CELL inst_17_16(
		.A1(out_sel[34]),
		.A2(I34[16]),
		.B1(out_sel[35]),
		.B2(I35[16]),
		.Z(O17[16])
	);
	AO_CELL inst_18_16(
		.A1(out_sel[36]),
		.A2(I36[16]),
		.B1(out_sel[37]),
		.B2(I37[16]),
		.Z(O18[16])
	);
	AO_CELL inst_19_16(
		.A1(out_sel[38]),
		.A2(I38[16]),
		.B1(out_sel[39]),
		.B2(I39[16]),
		.Z(O19[16])
	);
	AO_CELL inst_20_16(
		.A1(out_sel[40]),
		.A2(I40[16]),
		.B1(out_sel[41]),
		.B2(I41[16]),
		.Z(O20[16])
	);
	AO_CELL inst_21_16(
		.A1(out_sel[42]),
		.A2(I42[16]),
		.B1(out_sel[43]),
		.B2(I43[16]),
		.Z(O21[16])
	);
	AO_CELL inst_22_16(
		.A1(out_sel[44]),
		.A2(I44[16]),
		.B1(out_sel[45]),
		.B2(I45[16]),
		.Z(O22[16])
	);
	AN_CELL inst_and_16(
		.A1(out_sel[46]),
		.A2(I46[16]),
		.Z(O23[16])
	);
	AO_CELL inst_0_17(
		.A1(out_sel[0]),
		.A2(I0[17]),
		.B1(out_sel[1]),
		.B2(I1[17]),
		.Z(O0[17])
	);
	AO_CELL inst_1_17(
		.A1(out_sel[2]),
		.A2(I2[17]),
		.B1(out_sel[3]),
		.B2(I3[17]),
		.Z(O1[17])
	);
	AO_CELL inst_2_17(
		.A1(out_sel[4]),
		.A2(I4[17]),
		.B1(out_sel[5]),
		.B2(I5[17]),
		.Z(O2[17])
	);
	AO_CELL inst_3_17(
		.A1(out_sel[6]),
		.A2(I6[17]),
		.B1(out_sel[7]),
		.B2(I7[17]),
		.Z(O3[17])
	);
	AO_CELL inst_4_17(
		.A1(out_sel[8]),
		.A2(I8[17]),
		.B1(out_sel[9]),
		.B2(I9[17]),
		.Z(O4[17])
	);
	AO_CELL inst_5_17(
		.A1(out_sel[10]),
		.A2(I10[17]),
		.B1(out_sel[11]),
		.B2(I11[17]),
		.Z(O5[17])
	);
	AO_CELL inst_6_17(
		.A1(out_sel[12]),
		.A2(I12[17]),
		.B1(out_sel[13]),
		.B2(I13[17]),
		.Z(O6[17])
	);
	AO_CELL inst_7_17(
		.A1(out_sel[14]),
		.A2(I14[17]),
		.B1(out_sel[15]),
		.B2(I15[17]),
		.Z(O7[17])
	);
	AO_CELL inst_8_17(
		.A1(out_sel[16]),
		.A2(I16[17]),
		.B1(out_sel[17]),
		.B2(I17[17]),
		.Z(O8[17])
	);
	AO_CELL inst_9_17(
		.A1(out_sel[18]),
		.A2(I18[17]),
		.B1(out_sel[19]),
		.B2(I19[17]),
		.Z(O9[17])
	);
	AO_CELL inst_10_17(
		.A1(out_sel[20]),
		.A2(I20[17]),
		.B1(out_sel[21]),
		.B2(I21[17]),
		.Z(O10[17])
	);
	AO_CELL inst_11_17(
		.A1(out_sel[22]),
		.A2(I22[17]),
		.B1(out_sel[23]),
		.B2(I23[17]),
		.Z(O11[17])
	);
	AO_CELL inst_12_17(
		.A1(out_sel[24]),
		.A2(I24[17]),
		.B1(out_sel[25]),
		.B2(I25[17]),
		.Z(O12[17])
	);
	AO_CELL inst_13_17(
		.A1(out_sel[26]),
		.A2(I26[17]),
		.B1(out_sel[27]),
		.B2(I27[17]),
		.Z(O13[17])
	);
	AO_CELL inst_14_17(
		.A1(out_sel[28]),
		.A2(I28[17]),
		.B1(out_sel[29]),
		.B2(I29[17]),
		.Z(O14[17])
	);
	AO_CELL inst_15_17(
		.A1(out_sel[30]),
		.A2(I30[17]),
		.B1(out_sel[31]),
		.B2(I31[17]),
		.Z(O15[17])
	);
	AO_CELL inst_16_17(
		.A1(out_sel[32]),
		.A2(I32[17]),
		.B1(out_sel[33]),
		.B2(I33[17]),
		.Z(O16[17])
	);
	AO_CELL inst_17_17(
		.A1(out_sel[34]),
		.A2(I34[17]),
		.B1(out_sel[35]),
		.B2(I35[17]),
		.Z(O17[17])
	);
	AO_CELL inst_18_17(
		.A1(out_sel[36]),
		.A2(I36[17]),
		.B1(out_sel[37]),
		.B2(I37[17]),
		.Z(O18[17])
	);
	AO_CELL inst_19_17(
		.A1(out_sel[38]),
		.A2(I38[17]),
		.B1(out_sel[39]),
		.B2(I39[17]),
		.Z(O19[17])
	);
	AO_CELL inst_20_17(
		.A1(out_sel[40]),
		.A2(I40[17]),
		.B1(out_sel[41]),
		.B2(I41[17]),
		.Z(O20[17])
	);
	AO_CELL inst_21_17(
		.A1(out_sel[42]),
		.A2(I42[17]),
		.B1(out_sel[43]),
		.B2(I43[17]),
		.Z(O21[17])
	);
	AO_CELL inst_22_17(
		.A1(out_sel[44]),
		.A2(I44[17]),
		.B1(out_sel[45]),
		.B2(I45[17]),
		.Z(O22[17])
	);
	AN_CELL inst_and_17(
		.A1(out_sel[46]),
		.A2(I46[17]),
		.Z(O23[17])
	);
	AO_CELL inst_0_18(
		.A1(out_sel[0]),
		.A2(I0[18]),
		.B1(out_sel[1]),
		.B2(I1[18]),
		.Z(O0[18])
	);
	AO_CELL inst_1_18(
		.A1(out_sel[2]),
		.A2(I2[18]),
		.B1(out_sel[3]),
		.B2(I3[18]),
		.Z(O1[18])
	);
	AO_CELL inst_2_18(
		.A1(out_sel[4]),
		.A2(I4[18]),
		.B1(out_sel[5]),
		.B2(I5[18]),
		.Z(O2[18])
	);
	AO_CELL inst_3_18(
		.A1(out_sel[6]),
		.A2(I6[18]),
		.B1(out_sel[7]),
		.B2(I7[18]),
		.Z(O3[18])
	);
	AO_CELL inst_4_18(
		.A1(out_sel[8]),
		.A2(I8[18]),
		.B1(out_sel[9]),
		.B2(I9[18]),
		.Z(O4[18])
	);
	AO_CELL inst_5_18(
		.A1(out_sel[10]),
		.A2(I10[18]),
		.B1(out_sel[11]),
		.B2(I11[18]),
		.Z(O5[18])
	);
	AO_CELL inst_6_18(
		.A1(out_sel[12]),
		.A2(I12[18]),
		.B1(out_sel[13]),
		.B2(I13[18]),
		.Z(O6[18])
	);
	AO_CELL inst_7_18(
		.A1(out_sel[14]),
		.A2(I14[18]),
		.B1(out_sel[15]),
		.B2(I15[18]),
		.Z(O7[18])
	);
	AO_CELL inst_8_18(
		.A1(out_sel[16]),
		.A2(I16[18]),
		.B1(out_sel[17]),
		.B2(I17[18]),
		.Z(O8[18])
	);
	AO_CELL inst_9_18(
		.A1(out_sel[18]),
		.A2(I18[18]),
		.B1(out_sel[19]),
		.B2(I19[18]),
		.Z(O9[18])
	);
	AO_CELL inst_10_18(
		.A1(out_sel[20]),
		.A2(I20[18]),
		.B1(out_sel[21]),
		.B2(I21[18]),
		.Z(O10[18])
	);
	AO_CELL inst_11_18(
		.A1(out_sel[22]),
		.A2(I22[18]),
		.B1(out_sel[23]),
		.B2(I23[18]),
		.Z(O11[18])
	);
	AO_CELL inst_12_18(
		.A1(out_sel[24]),
		.A2(I24[18]),
		.B1(out_sel[25]),
		.B2(I25[18]),
		.Z(O12[18])
	);
	AO_CELL inst_13_18(
		.A1(out_sel[26]),
		.A2(I26[18]),
		.B1(out_sel[27]),
		.B2(I27[18]),
		.Z(O13[18])
	);
	AO_CELL inst_14_18(
		.A1(out_sel[28]),
		.A2(I28[18]),
		.B1(out_sel[29]),
		.B2(I29[18]),
		.Z(O14[18])
	);
	AO_CELL inst_15_18(
		.A1(out_sel[30]),
		.A2(I30[18]),
		.B1(out_sel[31]),
		.B2(I31[18]),
		.Z(O15[18])
	);
	AO_CELL inst_16_18(
		.A1(out_sel[32]),
		.A2(I32[18]),
		.B1(out_sel[33]),
		.B2(I33[18]),
		.Z(O16[18])
	);
	AO_CELL inst_17_18(
		.A1(out_sel[34]),
		.A2(I34[18]),
		.B1(out_sel[35]),
		.B2(I35[18]),
		.Z(O17[18])
	);
	AO_CELL inst_18_18(
		.A1(out_sel[36]),
		.A2(I36[18]),
		.B1(out_sel[37]),
		.B2(I37[18]),
		.Z(O18[18])
	);
	AO_CELL inst_19_18(
		.A1(out_sel[38]),
		.A2(I38[18]),
		.B1(out_sel[39]),
		.B2(I39[18]),
		.Z(O19[18])
	);
	AO_CELL inst_20_18(
		.A1(out_sel[40]),
		.A2(I40[18]),
		.B1(out_sel[41]),
		.B2(I41[18]),
		.Z(O20[18])
	);
	AO_CELL inst_21_18(
		.A1(out_sel[42]),
		.A2(I42[18]),
		.B1(out_sel[43]),
		.B2(I43[18]),
		.Z(O21[18])
	);
	AO_CELL inst_22_18(
		.A1(out_sel[44]),
		.A2(I44[18]),
		.B1(out_sel[45]),
		.B2(I45[18]),
		.Z(O22[18])
	);
	AN_CELL inst_and_18(
		.A1(out_sel[46]),
		.A2(I46[18]),
		.Z(O23[18])
	);
	AO_CELL inst_0_19(
		.A1(out_sel[0]),
		.A2(I0[19]),
		.B1(out_sel[1]),
		.B2(I1[19]),
		.Z(O0[19])
	);
	AO_CELL inst_1_19(
		.A1(out_sel[2]),
		.A2(I2[19]),
		.B1(out_sel[3]),
		.B2(I3[19]),
		.Z(O1[19])
	);
	AO_CELL inst_2_19(
		.A1(out_sel[4]),
		.A2(I4[19]),
		.B1(out_sel[5]),
		.B2(I5[19]),
		.Z(O2[19])
	);
	AO_CELL inst_3_19(
		.A1(out_sel[6]),
		.A2(I6[19]),
		.B1(out_sel[7]),
		.B2(I7[19]),
		.Z(O3[19])
	);
	AO_CELL inst_4_19(
		.A1(out_sel[8]),
		.A2(I8[19]),
		.B1(out_sel[9]),
		.B2(I9[19]),
		.Z(O4[19])
	);
	AO_CELL inst_5_19(
		.A1(out_sel[10]),
		.A2(I10[19]),
		.B1(out_sel[11]),
		.B2(I11[19]),
		.Z(O5[19])
	);
	AO_CELL inst_6_19(
		.A1(out_sel[12]),
		.A2(I12[19]),
		.B1(out_sel[13]),
		.B2(I13[19]),
		.Z(O6[19])
	);
	AO_CELL inst_7_19(
		.A1(out_sel[14]),
		.A2(I14[19]),
		.B1(out_sel[15]),
		.B2(I15[19]),
		.Z(O7[19])
	);
	AO_CELL inst_8_19(
		.A1(out_sel[16]),
		.A2(I16[19]),
		.B1(out_sel[17]),
		.B2(I17[19]),
		.Z(O8[19])
	);
	AO_CELL inst_9_19(
		.A1(out_sel[18]),
		.A2(I18[19]),
		.B1(out_sel[19]),
		.B2(I19[19]),
		.Z(O9[19])
	);
	AO_CELL inst_10_19(
		.A1(out_sel[20]),
		.A2(I20[19]),
		.B1(out_sel[21]),
		.B2(I21[19]),
		.Z(O10[19])
	);
	AO_CELL inst_11_19(
		.A1(out_sel[22]),
		.A2(I22[19]),
		.B1(out_sel[23]),
		.B2(I23[19]),
		.Z(O11[19])
	);
	AO_CELL inst_12_19(
		.A1(out_sel[24]),
		.A2(I24[19]),
		.B1(out_sel[25]),
		.B2(I25[19]),
		.Z(O12[19])
	);
	AO_CELL inst_13_19(
		.A1(out_sel[26]),
		.A2(I26[19]),
		.B1(out_sel[27]),
		.B2(I27[19]),
		.Z(O13[19])
	);
	AO_CELL inst_14_19(
		.A1(out_sel[28]),
		.A2(I28[19]),
		.B1(out_sel[29]),
		.B2(I29[19]),
		.Z(O14[19])
	);
	AO_CELL inst_15_19(
		.A1(out_sel[30]),
		.A2(I30[19]),
		.B1(out_sel[31]),
		.B2(I31[19]),
		.Z(O15[19])
	);
	AO_CELL inst_16_19(
		.A1(out_sel[32]),
		.A2(I32[19]),
		.B1(out_sel[33]),
		.B2(I33[19]),
		.Z(O16[19])
	);
	AO_CELL inst_17_19(
		.A1(out_sel[34]),
		.A2(I34[19]),
		.B1(out_sel[35]),
		.B2(I35[19]),
		.Z(O17[19])
	);
	AO_CELL inst_18_19(
		.A1(out_sel[36]),
		.A2(I36[19]),
		.B1(out_sel[37]),
		.B2(I37[19]),
		.Z(O18[19])
	);
	AO_CELL inst_19_19(
		.A1(out_sel[38]),
		.A2(I38[19]),
		.B1(out_sel[39]),
		.B2(I39[19]),
		.Z(O19[19])
	);
	AO_CELL inst_20_19(
		.A1(out_sel[40]),
		.A2(I40[19]),
		.B1(out_sel[41]),
		.B2(I41[19]),
		.Z(O20[19])
	);
	AO_CELL inst_21_19(
		.A1(out_sel[42]),
		.A2(I42[19]),
		.B1(out_sel[43]),
		.B2(I43[19]),
		.Z(O21[19])
	);
	AO_CELL inst_22_19(
		.A1(out_sel[44]),
		.A2(I44[19]),
		.B1(out_sel[45]),
		.B2(I45[19]),
		.Z(O22[19])
	);
	AN_CELL inst_and_19(
		.A1(out_sel[46]),
		.A2(I46[19]),
		.Z(O23[19])
	);
	AO_CELL inst_0_20(
		.A1(out_sel[0]),
		.A2(I0[20]),
		.B1(out_sel[1]),
		.B2(I1[20]),
		.Z(O0[20])
	);
	AO_CELL inst_1_20(
		.A1(out_sel[2]),
		.A2(I2[20]),
		.B1(out_sel[3]),
		.B2(I3[20]),
		.Z(O1[20])
	);
	AO_CELL inst_2_20(
		.A1(out_sel[4]),
		.A2(I4[20]),
		.B1(out_sel[5]),
		.B2(I5[20]),
		.Z(O2[20])
	);
	AO_CELL inst_3_20(
		.A1(out_sel[6]),
		.A2(I6[20]),
		.B1(out_sel[7]),
		.B2(I7[20]),
		.Z(O3[20])
	);
	AO_CELL inst_4_20(
		.A1(out_sel[8]),
		.A2(I8[20]),
		.B1(out_sel[9]),
		.B2(I9[20]),
		.Z(O4[20])
	);
	AO_CELL inst_5_20(
		.A1(out_sel[10]),
		.A2(I10[20]),
		.B1(out_sel[11]),
		.B2(I11[20]),
		.Z(O5[20])
	);
	AO_CELL inst_6_20(
		.A1(out_sel[12]),
		.A2(I12[20]),
		.B1(out_sel[13]),
		.B2(I13[20]),
		.Z(O6[20])
	);
	AO_CELL inst_7_20(
		.A1(out_sel[14]),
		.A2(I14[20]),
		.B1(out_sel[15]),
		.B2(I15[20]),
		.Z(O7[20])
	);
	AO_CELL inst_8_20(
		.A1(out_sel[16]),
		.A2(I16[20]),
		.B1(out_sel[17]),
		.B2(I17[20]),
		.Z(O8[20])
	);
	AO_CELL inst_9_20(
		.A1(out_sel[18]),
		.A2(I18[20]),
		.B1(out_sel[19]),
		.B2(I19[20]),
		.Z(O9[20])
	);
	AO_CELL inst_10_20(
		.A1(out_sel[20]),
		.A2(I20[20]),
		.B1(out_sel[21]),
		.B2(I21[20]),
		.Z(O10[20])
	);
	AO_CELL inst_11_20(
		.A1(out_sel[22]),
		.A2(I22[20]),
		.B1(out_sel[23]),
		.B2(I23[20]),
		.Z(O11[20])
	);
	AO_CELL inst_12_20(
		.A1(out_sel[24]),
		.A2(I24[20]),
		.B1(out_sel[25]),
		.B2(I25[20]),
		.Z(O12[20])
	);
	AO_CELL inst_13_20(
		.A1(out_sel[26]),
		.A2(I26[20]),
		.B1(out_sel[27]),
		.B2(I27[20]),
		.Z(O13[20])
	);
	AO_CELL inst_14_20(
		.A1(out_sel[28]),
		.A2(I28[20]),
		.B1(out_sel[29]),
		.B2(I29[20]),
		.Z(O14[20])
	);
	AO_CELL inst_15_20(
		.A1(out_sel[30]),
		.A2(I30[20]),
		.B1(out_sel[31]),
		.B2(I31[20]),
		.Z(O15[20])
	);
	AO_CELL inst_16_20(
		.A1(out_sel[32]),
		.A2(I32[20]),
		.B1(out_sel[33]),
		.B2(I33[20]),
		.Z(O16[20])
	);
	AO_CELL inst_17_20(
		.A1(out_sel[34]),
		.A2(I34[20]),
		.B1(out_sel[35]),
		.B2(I35[20]),
		.Z(O17[20])
	);
	AO_CELL inst_18_20(
		.A1(out_sel[36]),
		.A2(I36[20]),
		.B1(out_sel[37]),
		.B2(I37[20]),
		.Z(O18[20])
	);
	AO_CELL inst_19_20(
		.A1(out_sel[38]),
		.A2(I38[20]),
		.B1(out_sel[39]),
		.B2(I39[20]),
		.Z(O19[20])
	);
	AO_CELL inst_20_20(
		.A1(out_sel[40]),
		.A2(I40[20]),
		.B1(out_sel[41]),
		.B2(I41[20]),
		.Z(O20[20])
	);
	AO_CELL inst_21_20(
		.A1(out_sel[42]),
		.A2(I42[20]),
		.B1(out_sel[43]),
		.B2(I43[20]),
		.Z(O21[20])
	);
	AO_CELL inst_22_20(
		.A1(out_sel[44]),
		.A2(I44[20]),
		.B1(out_sel[45]),
		.B2(I45[20]),
		.Z(O22[20])
	);
	AN_CELL inst_and_20(
		.A1(out_sel[46]),
		.A2(I46[20]),
		.Z(O23[20])
	);
	AO_CELL inst_0_21(
		.A1(out_sel[0]),
		.A2(I0[21]),
		.B1(out_sel[1]),
		.B2(I1[21]),
		.Z(O0[21])
	);
	AO_CELL inst_1_21(
		.A1(out_sel[2]),
		.A2(I2[21]),
		.B1(out_sel[3]),
		.B2(I3[21]),
		.Z(O1[21])
	);
	AO_CELL inst_2_21(
		.A1(out_sel[4]),
		.A2(I4[21]),
		.B1(out_sel[5]),
		.B2(I5[21]),
		.Z(O2[21])
	);
	AO_CELL inst_3_21(
		.A1(out_sel[6]),
		.A2(I6[21]),
		.B1(out_sel[7]),
		.B2(I7[21]),
		.Z(O3[21])
	);
	AO_CELL inst_4_21(
		.A1(out_sel[8]),
		.A2(I8[21]),
		.B1(out_sel[9]),
		.B2(I9[21]),
		.Z(O4[21])
	);
	AO_CELL inst_5_21(
		.A1(out_sel[10]),
		.A2(I10[21]),
		.B1(out_sel[11]),
		.B2(I11[21]),
		.Z(O5[21])
	);
	AO_CELL inst_6_21(
		.A1(out_sel[12]),
		.A2(I12[21]),
		.B1(out_sel[13]),
		.B2(I13[21]),
		.Z(O6[21])
	);
	AO_CELL inst_7_21(
		.A1(out_sel[14]),
		.A2(I14[21]),
		.B1(out_sel[15]),
		.B2(I15[21]),
		.Z(O7[21])
	);
	AO_CELL inst_8_21(
		.A1(out_sel[16]),
		.A2(I16[21]),
		.B1(out_sel[17]),
		.B2(I17[21]),
		.Z(O8[21])
	);
	AO_CELL inst_9_21(
		.A1(out_sel[18]),
		.A2(I18[21]),
		.B1(out_sel[19]),
		.B2(I19[21]),
		.Z(O9[21])
	);
	AO_CELL inst_10_21(
		.A1(out_sel[20]),
		.A2(I20[21]),
		.B1(out_sel[21]),
		.B2(I21[21]),
		.Z(O10[21])
	);
	AO_CELL inst_11_21(
		.A1(out_sel[22]),
		.A2(I22[21]),
		.B1(out_sel[23]),
		.B2(I23[21]),
		.Z(O11[21])
	);
	AO_CELL inst_12_21(
		.A1(out_sel[24]),
		.A2(I24[21]),
		.B1(out_sel[25]),
		.B2(I25[21]),
		.Z(O12[21])
	);
	AO_CELL inst_13_21(
		.A1(out_sel[26]),
		.A2(I26[21]),
		.B1(out_sel[27]),
		.B2(I27[21]),
		.Z(O13[21])
	);
	AO_CELL inst_14_21(
		.A1(out_sel[28]),
		.A2(I28[21]),
		.B1(out_sel[29]),
		.B2(I29[21]),
		.Z(O14[21])
	);
	AO_CELL inst_15_21(
		.A1(out_sel[30]),
		.A2(I30[21]),
		.B1(out_sel[31]),
		.B2(I31[21]),
		.Z(O15[21])
	);
	AO_CELL inst_16_21(
		.A1(out_sel[32]),
		.A2(I32[21]),
		.B1(out_sel[33]),
		.B2(I33[21]),
		.Z(O16[21])
	);
	AO_CELL inst_17_21(
		.A1(out_sel[34]),
		.A2(I34[21]),
		.B1(out_sel[35]),
		.B2(I35[21]),
		.Z(O17[21])
	);
	AO_CELL inst_18_21(
		.A1(out_sel[36]),
		.A2(I36[21]),
		.B1(out_sel[37]),
		.B2(I37[21]),
		.Z(O18[21])
	);
	AO_CELL inst_19_21(
		.A1(out_sel[38]),
		.A2(I38[21]),
		.B1(out_sel[39]),
		.B2(I39[21]),
		.Z(O19[21])
	);
	AO_CELL inst_20_21(
		.A1(out_sel[40]),
		.A2(I40[21]),
		.B1(out_sel[41]),
		.B2(I41[21]),
		.Z(O20[21])
	);
	AO_CELL inst_21_21(
		.A1(out_sel[42]),
		.A2(I42[21]),
		.B1(out_sel[43]),
		.B2(I43[21]),
		.Z(O21[21])
	);
	AO_CELL inst_22_21(
		.A1(out_sel[44]),
		.A2(I44[21]),
		.B1(out_sel[45]),
		.B2(I45[21]),
		.Z(O22[21])
	);
	AN_CELL inst_and_21(
		.A1(out_sel[46]),
		.A2(I46[21]),
		.Z(O23[21])
	);
	AO_CELL inst_0_22(
		.A1(out_sel[0]),
		.A2(I0[22]),
		.B1(out_sel[1]),
		.B2(I1[22]),
		.Z(O0[22])
	);
	AO_CELL inst_1_22(
		.A1(out_sel[2]),
		.A2(I2[22]),
		.B1(out_sel[3]),
		.B2(I3[22]),
		.Z(O1[22])
	);
	AO_CELL inst_2_22(
		.A1(out_sel[4]),
		.A2(I4[22]),
		.B1(out_sel[5]),
		.B2(I5[22]),
		.Z(O2[22])
	);
	AO_CELL inst_3_22(
		.A1(out_sel[6]),
		.A2(I6[22]),
		.B1(out_sel[7]),
		.B2(I7[22]),
		.Z(O3[22])
	);
	AO_CELL inst_4_22(
		.A1(out_sel[8]),
		.A2(I8[22]),
		.B1(out_sel[9]),
		.B2(I9[22]),
		.Z(O4[22])
	);
	AO_CELL inst_5_22(
		.A1(out_sel[10]),
		.A2(I10[22]),
		.B1(out_sel[11]),
		.B2(I11[22]),
		.Z(O5[22])
	);
	AO_CELL inst_6_22(
		.A1(out_sel[12]),
		.A2(I12[22]),
		.B1(out_sel[13]),
		.B2(I13[22]),
		.Z(O6[22])
	);
	AO_CELL inst_7_22(
		.A1(out_sel[14]),
		.A2(I14[22]),
		.B1(out_sel[15]),
		.B2(I15[22]),
		.Z(O7[22])
	);
	AO_CELL inst_8_22(
		.A1(out_sel[16]),
		.A2(I16[22]),
		.B1(out_sel[17]),
		.B2(I17[22]),
		.Z(O8[22])
	);
	AO_CELL inst_9_22(
		.A1(out_sel[18]),
		.A2(I18[22]),
		.B1(out_sel[19]),
		.B2(I19[22]),
		.Z(O9[22])
	);
	AO_CELL inst_10_22(
		.A1(out_sel[20]),
		.A2(I20[22]),
		.B1(out_sel[21]),
		.B2(I21[22]),
		.Z(O10[22])
	);
	AO_CELL inst_11_22(
		.A1(out_sel[22]),
		.A2(I22[22]),
		.B1(out_sel[23]),
		.B2(I23[22]),
		.Z(O11[22])
	);
	AO_CELL inst_12_22(
		.A1(out_sel[24]),
		.A2(I24[22]),
		.B1(out_sel[25]),
		.B2(I25[22]),
		.Z(O12[22])
	);
	AO_CELL inst_13_22(
		.A1(out_sel[26]),
		.A2(I26[22]),
		.B1(out_sel[27]),
		.B2(I27[22]),
		.Z(O13[22])
	);
	AO_CELL inst_14_22(
		.A1(out_sel[28]),
		.A2(I28[22]),
		.B1(out_sel[29]),
		.B2(I29[22]),
		.Z(O14[22])
	);
	AO_CELL inst_15_22(
		.A1(out_sel[30]),
		.A2(I30[22]),
		.B1(out_sel[31]),
		.B2(I31[22]),
		.Z(O15[22])
	);
	AO_CELL inst_16_22(
		.A1(out_sel[32]),
		.A2(I32[22]),
		.B1(out_sel[33]),
		.B2(I33[22]),
		.Z(O16[22])
	);
	AO_CELL inst_17_22(
		.A1(out_sel[34]),
		.A2(I34[22]),
		.B1(out_sel[35]),
		.B2(I35[22]),
		.Z(O17[22])
	);
	AO_CELL inst_18_22(
		.A1(out_sel[36]),
		.A2(I36[22]),
		.B1(out_sel[37]),
		.B2(I37[22]),
		.Z(O18[22])
	);
	AO_CELL inst_19_22(
		.A1(out_sel[38]),
		.A2(I38[22]),
		.B1(out_sel[39]),
		.B2(I39[22]),
		.Z(O19[22])
	);
	AO_CELL inst_20_22(
		.A1(out_sel[40]),
		.A2(I40[22]),
		.B1(out_sel[41]),
		.B2(I41[22]),
		.Z(O20[22])
	);
	AO_CELL inst_21_22(
		.A1(out_sel[42]),
		.A2(I42[22]),
		.B1(out_sel[43]),
		.B2(I43[22]),
		.Z(O21[22])
	);
	AO_CELL inst_22_22(
		.A1(out_sel[44]),
		.A2(I44[22]),
		.B1(out_sel[45]),
		.B2(I45[22]),
		.Z(O22[22])
	);
	AN_CELL inst_and_22(
		.A1(out_sel[46]),
		.A2(I46[22]),
		.Z(O23[22])
	);
	AO_CELL inst_0_23(
		.A1(out_sel[0]),
		.A2(I0[23]),
		.B1(out_sel[1]),
		.B2(I1[23]),
		.Z(O0[23])
	);
	AO_CELL inst_1_23(
		.A1(out_sel[2]),
		.A2(I2[23]),
		.B1(out_sel[3]),
		.B2(I3[23]),
		.Z(O1[23])
	);
	AO_CELL inst_2_23(
		.A1(out_sel[4]),
		.A2(I4[23]),
		.B1(out_sel[5]),
		.B2(I5[23]),
		.Z(O2[23])
	);
	AO_CELL inst_3_23(
		.A1(out_sel[6]),
		.A2(I6[23]),
		.B1(out_sel[7]),
		.B2(I7[23]),
		.Z(O3[23])
	);
	AO_CELL inst_4_23(
		.A1(out_sel[8]),
		.A2(I8[23]),
		.B1(out_sel[9]),
		.B2(I9[23]),
		.Z(O4[23])
	);
	AO_CELL inst_5_23(
		.A1(out_sel[10]),
		.A2(I10[23]),
		.B1(out_sel[11]),
		.B2(I11[23]),
		.Z(O5[23])
	);
	AO_CELL inst_6_23(
		.A1(out_sel[12]),
		.A2(I12[23]),
		.B1(out_sel[13]),
		.B2(I13[23]),
		.Z(O6[23])
	);
	AO_CELL inst_7_23(
		.A1(out_sel[14]),
		.A2(I14[23]),
		.B1(out_sel[15]),
		.B2(I15[23]),
		.Z(O7[23])
	);
	AO_CELL inst_8_23(
		.A1(out_sel[16]),
		.A2(I16[23]),
		.B1(out_sel[17]),
		.B2(I17[23]),
		.Z(O8[23])
	);
	AO_CELL inst_9_23(
		.A1(out_sel[18]),
		.A2(I18[23]),
		.B1(out_sel[19]),
		.B2(I19[23]),
		.Z(O9[23])
	);
	AO_CELL inst_10_23(
		.A1(out_sel[20]),
		.A2(I20[23]),
		.B1(out_sel[21]),
		.B2(I21[23]),
		.Z(O10[23])
	);
	AO_CELL inst_11_23(
		.A1(out_sel[22]),
		.A2(I22[23]),
		.B1(out_sel[23]),
		.B2(I23[23]),
		.Z(O11[23])
	);
	AO_CELL inst_12_23(
		.A1(out_sel[24]),
		.A2(I24[23]),
		.B1(out_sel[25]),
		.B2(I25[23]),
		.Z(O12[23])
	);
	AO_CELL inst_13_23(
		.A1(out_sel[26]),
		.A2(I26[23]),
		.B1(out_sel[27]),
		.B2(I27[23]),
		.Z(O13[23])
	);
	AO_CELL inst_14_23(
		.A1(out_sel[28]),
		.A2(I28[23]),
		.B1(out_sel[29]),
		.B2(I29[23]),
		.Z(O14[23])
	);
	AO_CELL inst_15_23(
		.A1(out_sel[30]),
		.A2(I30[23]),
		.B1(out_sel[31]),
		.B2(I31[23]),
		.Z(O15[23])
	);
	AO_CELL inst_16_23(
		.A1(out_sel[32]),
		.A2(I32[23]),
		.B1(out_sel[33]),
		.B2(I33[23]),
		.Z(O16[23])
	);
	AO_CELL inst_17_23(
		.A1(out_sel[34]),
		.A2(I34[23]),
		.B1(out_sel[35]),
		.B2(I35[23]),
		.Z(O17[23])
	);
	AO_CELL inst_18_23(
		.A1(out_sel[36]),
		.A2(I36[23]),
		.B1(out_sel[37]),
		.B2(I37[23]),
		.Z(O18[23])
	);
	AO_CELL inst_19_23(
		.A1(out_sel[38]),
		.A2(I38[23]),
		.B1(out_sel[39]),
		.B2(I39[23]),
		.Z(O19[23])
	);
	AO_CELL inst_20_23(
		.A1(out_sel[40]),
		.A2(I40[23]),
		.B1(out_sel[41]),
		.B2(I41[23]),
		.Z(O20[23])
	);
	AO_CELL inst_21_23(
		.A1(out_sel[42]),
		.A2(I42[23]),
		.B1(out_sel[43]),
		.B2(I43[23]),
		.Z(O21[23])
	);
	AO_CELL inst_22_23(
		.A1(out_sel[44]),
		.A2(I44[23]),
		.B1(out_sel[45]),
		.B2(I45[23]),
		.Z(O22[23])
	);
	AN_CELL inst_and_23(
		.A1(out_sel[46]),
		.A2(I46[23]),
		.Z(O23[23])
	);
	AO_CELL inst_0_24(
		.A1(out_sel[0]),
		.A2(I0[24]),
		.B1(out_sel[1]),
		.B2(I1[24]),
		.Z(O0[24])
	);
	AO_CELL inst_1_24(
		.A1(out_sel[2]),
		.A2(I2[24]),
		.B1(out_sel[3]),
		.B2(I3[24]),
		.Z(O1[24])
	);
	AO_CELL inst_2_24(
		.A1(out_sel[4]),
		.A2(I4[24]),
		.B1(out_sel[5]),
		.B2(I5[24]),
		.Z(O2[24])
	);
	AO_CELL inst_3_24(
		.A1(out_sel[6]),
		.A2(I6[24]),
		.B1(out_sel[7]),
		.B2(I7[24]),
		.Z(O3[24])
	);
	AO_CELL inst_4_24(
		.A1(out_sel[8]),
		.A2(I8[24]),
		.B1(out_sel[9]),
		.B2(I9[24]),
		.Z(O4[24])
	);
	AO_CELL inst_5_24(
		.A1(out_sel[10]),
		.A2(I10[24]),
		.B1(out_sel[11]),
		.B2(I11[24]),
		.Z(O5[24])
	);
	AO_CELL inst_6_24(
		.A1(out_sel[12]),
		.A2(I12[24]),
		.B1(out_sel[13]),
		.B2(I13[24]),
		.Z(O6[24])
	);
	AO_CELL inst_7_24(
		.A1(out_sel[14]),
		.A2(I14[24]),
		.B1(out_sel[15]),
		.B2(I15[24]),
		.Z(O7[24])
	);
	AO_CELL inst_8_24(
		.A1(out_sel[16]),
		.A2(I16[24]),
		.B1(out_sel[17]),
		.B2(I17[24]),
		.Z(O8[24])
	);
	AO_CELL inst_9_24(
		.A1(out_sel[18]),
		.A2(I18[24]),
		.B1(out_sel[19]),
		.B2(I19[24]),
		.Z(O9[24])
	);
	AO_CELL inst_10_24(
		.A1(out_sel[20]),
		.A2(I20[24]),
		.B1(out_sel[21]),
		.B2(I21[24]),
		.Z(O10[24])
	);
	AO_CELL inst_11_24(
		.A1(out_sel[22]),
		.A2(I22[24]),
		.B1(out_sel[23]),
		.B2(I23[24]),
		.Z(O11[24])
	);
	AO_CELL inst_12_24(
		.A1(out_sel[24]),
		.A2(I24[24]),
		.B1(out_sel[25]),
		.B2(I25[24]),
		.Z(O12[24])
	);
	AO_CELL inst_13_24(
		.A1(out_sel[26]),
		.A2(I26[24]),
		.B1(out_sel[27]),
		.B2(I27[24]),
		.Z(O13[24])
	);
	AO_CELL inst_14_24(
		.A1(out_sel[28]),
		.A2(I28[24]),
		.B1(out_sel[29]),
		.B2(I29[24]),
		.Z(O14[24])
	);
	AO_CELL inst_15_24(
		.A1(out_sel[30]),
		.A2(I30[24]),
		.B1(out_sel[31]),
		.B2(I31[24]),
		.Z(O15[24])
	);
	AO_CELL inst_16_24(
		.A1(out_sel[32]),
		.A2(I32[24]),
		.B1(out_sel[33]),
		.B2(I33[24]),
		.Z(O16[24])
	);
	AO_CELL inst_17_24(
		.A1(out_sel[34]),
		.A2(I34[24]),
		.B1(out_sel[35]),
		.B2(I35[24]),
		.Z(O17[24])
	);
	AO_CELL inst_18_24(
		.A1(out_sel[36]),
		.A2(I36[24]),
		.B1(out_sel[37]),
		.B2(I37[24]),
		.Z(O18[24])
	);
	AO_CELL inst_19_24(
		.A1(out_sel[38]),
		.A2(I38[24]),
		.B1(out_sel[39]),
		.B2(I39[24]),
		.Z(O19[24])
	);
	AO_CELL inst_20_24(
		.A1(out_sel[40]),
		.A2(I40[24]),
		.B1(out_sel[41]),
		.B2(I41[24]),
		.Z(O20[24])
	);
	AO_CELL inst_21_24(
		.A1(out_sel[42]),
		.A2(I42[24]),
		.B1(out_sel[43]),
		.B2(I43[24]),
		.Z(O21[24])
	);
	AO_CELL inst_22_24(
		.A1(out_sel[44]),
		.A2(I44[24]),
		.B1(out_sel[45]),
		.B2(I45[24]),
		.Z(O22[24])
	);
	AN_CELL inst_and_24(
		.A1(out_sel[46]),
		.A2(I46[24]),
		.Z(O23[24])
	);
	AO_CELL inst_0_25(
		.A1(out_sel[0]),
		.A2(I0[25]),
		.B1(out_sel[1]),
		.B2(I1[25]),
		.Z(O0[25])
	);
	AO_CELL inst_1_25(
		.A1(out_sel[2]),
		.A2(I2[25]),
		.B1(out_sel[3]),
		.B2(I3[25]),
		.Z(O1[25])
	);
	AO_CELL inst_2_25(
		.A1(out_sel[4]),
		.A2(I4[25]),
		.B1(out_sel[5]),
		.B2(I5[25]),
		.Z(O2[25])
	);
	AO_CELL inst_3_25(
		.A1(out_sel[6]),
		.A2(I6[25]),
		.B1(out_sel[7]),
		.B2(I7[25]),
		.Z(O3[25])
	);
	AO_CELL inst_4_25(
		.A1(out_sel[8]),
		.A2(I8[25]),
		.B1(out_sel[9]),
		.B2(I9[25]),
		.Z(O4[25])
	);
	AO_CELL inst_5_25(
		.A1(out_sel[10]),
		.A2(I10[25]),
		.B1(out_sel[11]),
		.B2(I11[25]),
		.Z(O5[25])
	);
	AO_CELL inst_6_25(
		.A1(out_sel[12]),
		.A2(I12[25]),
		.B1(out_sel[13]),
		.B2(I13[25]),
		.Z(O6[25])
	);
	AO_CELL inst_7_25(
		.A1(out_sel[14]),
		.A2(I14[25]),
		.B1(out_sel[15]),
		.B2(I15[25]),
		.Z(O7[25])
	);
	AO_CELL inst_8_25(
		.A1(out_sel[16]),
		.A2(I16[25]),
		.B1(out_sel[17]),
		.B2(I17[25]),
		.Z(O8[25])
	);
	AO_CELL inst_9_25(
		.A1(out_sel[18]),
		.A2(I18[25]),
		.B1(out_sel[19]),
		.B2(I19[25]),
		.Z(O9[25])
	);
	AO_CELL inst_10_25(
		.A1(out_sel[20]),
		.A2(I20[25]),
		.B1(out_sel[21]),
		.B2(I21[25]),
		.Z(O10[25])
	);
	AO_CELL inst_11_25(
		.A1(out_sel[22]),
		.A2(I22[25]),
		.B1(out_sel[23]),
		.B2(I23[25]),
		.Z(O11[25])
	);
	AO_CELL inst_12_25(
		.A1(out_sel[24]),
		.A2(I24[25]),
		.B1(out_sel[25]),
		.B2(I25[25]),
		.Z(O12[25])
	);
	AO_CELL inst_13_25(
		.A1(out_sel[26]),
		.A2(I26[25]),
		.B1(out_sel[27]),
		.B2(I27[25]),
		.Z(O13[25])
	);
	AO_CELL inst_14_25(
		.A1(out_sel[28]),
		.A2(I28[25]),
		.B1(out_sel[29]),
		.B2(I29[25]),
		.Z(O14[25])
	);
	AO_CELL inst_15_25(
		.A1(out_sel[30]),
		.A2(I30[25]),
		.B1(out_sel[31]),
		.B2(I31[25]),
		.Z(O15[25])
	);
	AO_CELL inst_16_25(
		.A1(out_sel[32]),
		.A2(I32[25]),
		.B1(out_sel[33]),
		.B2(I33[25]),
		.Z(O16[25])
	);
	AO_CELL inst_17_25(
		.A1(out_sel[34]),
		.A2(I34[25]),
		.B1(out_sel[35]),
		.B2(I35[25]),
		.Z(O17[25])
	);
	AO_CELL inst_18_25(
		.A1(out_sel[36]),
		.A2(I36[25]),
		.B1(out_sel[37]),
		.B2(I37[25]),
		.Z(O18[25])
	);
	AO_CELL inst_19_25(
		.A1(out_sel[38]),
		.A2(I38[25]),
		.B1(out_sel[39]),
		.B2(I39[25]),
		.Z(O19[25])
	);
	AO_CELL inst_20_25(
		.A1(out_sel[40]),
		.A2(I40[25]),
		.B1(out_sel[41]),
		.B2(I41[25]),
		.Z(O20[25])
	);
	AO_CELL inst_21_25(
		.A1(out_sel[42]),
		.A2(I42[25]),
		.B1(out_sel[43]),
		.B2(I43[25]),
		.Z(O21[25])
	);
	AO_CELL inst_22_25(
		.A1(out_sel[44]),
		.A2(I44[25]),
		.B1(out_sel[45]),
		.B2(I45[25]),
		.Z(O22[25])
	);
	AN_CELL inst_and_25(
		.A1(out_sel[46]),
		.A2(I46[25]),
		.Z(O23[25])
	);
	AO_CELL inst_0_26(
		.A1(out_sel[0]),
		.A2(I0[26]),
		.B1(out_sel[1]),
		.B2(I1[26]),
		.Z(O0[26])
	);
	AO_CELL inst_1_26(
		.A1(out_sel[2]),
		.A2(I2[26]),
		.B1(out_sel[3]),
		.B2(I3[26]),
		.Z(O1[26])
	);
	AO_CELL inst_2_26(
		.A1(out_sel[4]),
		.A2(I4[26]),
		.B1(out_sel[5]),
		.B2(I5[26]),
		.Z(O2[26])
	);
	AO_CELL inst_3_26(
		.A1(out_sel[6]),
		.A2(I6[26]),
		.B1(out_sel[7]),
		.B2(I7[26]),
		.Z(O3[26])
	);
	AO_CELL inst_4_26(
		.A1(out_sel[8]),
		.A2(I8[26]),
		.B1(out_sel[9]),
		.B2(I9[26]),
		.Z(O4[26])
	);
	AO_CELL inst_5_26(
		.A1(out_sel[10]),
		.A2(I10[26]),
		.B1(out_sel[11]),
		.B2(I11[26]),
		.Z(O5[26])
	);
	AO_CELL inst_6_26(
		.A1(out_sel[12]),
		.A2(I12[26]),
		.B1(out_sel[13]),
		.B2(I13[26]),
		.Z(O6[26])
	);
	AO_CELL inst_7_26(
		.A1(out_sel[14]),
		.A2(I14[26]),
		.B1(out_sel[15]),
		.B2(I15[26]),
		.Z(O7[26])
	);
	AO_CELL inst_8_26(
		.A1(out_sel[16]),
		.A2(I16[26]),
		.B1(out_sel[17]),
		.B2(I17[26]),
		.Z(O8[26])
	);
	AO_CELL inst_9_26(
		.A1(out_sel[18]),
		.A2(I18[26]),
		.B1(out_sel[19]),
		.B2(I19[26]),
		.Z(O9[26])
	);
	AO_CELL inst_10_26(
		.A1(out_sel[20]),
		.A2(I20[26]),
		.B1(out_sel[21]),
		.B2(I21[26]),
		.Z(O10[26])
	);
	AO_CELL inst_11_26(
		.A1(out_sel[22]),
		.A2(I22[26]),
		.B1(out_sel[23]),
		.B2(I23[26]),
		.Z(O11[26])
	);
	AO_CELL inst_12_26(
		.A1(out_sel[24]),
		.A2(I24[26]),
		.B1(out_sel[25]),
		.B2(I25[26]),
		.Z(O12[26])
	);
	AO_CELL inst_13_26(
		.A1(out_sel[26]),
		.A2(I26[26]),
		.B1(out_sel[27]),
		.B2(I27[26]),
		.Z(O13[26])
	);
	AO_CELL inst_14_26(
		.A1(out_sel[28]),
		.A2(I28[26]),
		.B1(out_sel[29]),
		.B2(I29[26]),
		.Z(O14[26])
	);
	AO_CELL inst_15_26(
		.A1(out_sel[30]),
		.A2(I30[26]),
		.B1(out_sel[31]),
		.B2(I31[26]),
		.Z(O15[26])
	);
	AO_CELL inst_16_26(
		.A1(out_sel[32]),
		.A2(I32[26]),
		.B1(out_sel[33]),
		.B2(I33[26]),
		.Z(O16[26])
	);
	AO_CELL inst_17_26(
		.A1(out_sel[34]),
		.A2(I34[26]),
		.B1(out_sel[35]),
		.B2(I35[26]),
		.Z(O17[26])
	);
	AO_CELL inst_18_26(
		.A1(out_sel[36]),
		.A2(I36[26]),
		.B1(out_sel[37]),
		.B2(I37[26]),
		.Z(O18[26])
	);
	AO_CELL inst_19_26(
		.A1(out_sel[38]),
		.A2(I38[26]),
		.B1(out_sel[39]),
		.B2(I39[26]),
		.Z(O19[26])
	);
	AO_CELL inst_20_26(
		.A1(out_sel[40]),
		.A2(I40[26]),
		.B1(out_sel[41]),
		.B2(I41[26]),
		.Z(O20[26])
	);
	AO_CELL inst_21_26(
		.A1(out_sel[42]),
		.A2(I42[26]),
		.B1(out_sel[43]),
		.B2(I43[26]),
		.Z(O21[26])
	);
	AO_CELL inst_22_26(
		.A1(out_sel[44]),
		.A2(I44[26]),
		.B1(out_sel[45]),
		.B2(I45[26]),
		.Z(O22[26])
	);
	AN_CELL inst_and_26(
		.A1(out_sel[46]),
		.A2(I46[26]),
		.Z(O23[26])
	);
	AO_CELL inst_0_27(
		.A1(out_sel[0]),
		.A2(I0[27]),
		.B1(out_sel[1]),
		.B2(I1[27]),
		.Z(O0[27])
	);
	AO_CELL inst_1_27(
		.A1(out_sel[2]),
		.A2(I2[27]),
		.B1(out_sel[3]),
		.B2(I3[27]),
		.Z(O1[27])
	);
	AO_CELL inst_2_27(
		.A1(out_sel[4]),
		.A2(I4[27]),
		.B1(out_sel[5]),
		.B2(I5[27]),
		.Z(O2[27])
	);
	AO_CELL inst_3_27(
		.A1(out_sel[6]),
		.A2(I6[27]),
		.B1(out_sel[7]),
		.B2(I7[27]),
		.Z(O3[27])
	);
	AO_CELL inst_4_27(
		.A1(out_sel[8]),
		.A2(I8[27]),
		.B1(out_sel[9]),
		.B2(I9[27]),
		.Z(O4[27])
	);
	AO_CELL inst_5_27(
		.A1(out_sel[10]),
		.A2(I10[27]),
		.B1(out_sel[11]),
		.B2(I11[27]),
		.Z(O5[27])
	);
	AO_CELL inst_6_27(
		.A1(out_sel[12]),
		.A2(I12[27]),
		.B1(out_sel[13]),
		.B2(I13[27]),
		.Z(O6[27])
	);
	AO_CELL inst_7_27(
		.A1(out_sel[14]),
		.A2(I14[27]),
		.B1(out_sel[15]),
		.B2(I15[27]),
		.Z(O7[27])
	);
	AO_CELL inst_8_27(
		.A1(out_sel[16]),
		.A2(I16[27]),
		.B1(out_sel[17]),
		.B2(I17[27]),
		.Z(O8[27])
	);
	AO_CELL inst_9_27(
		.A1(out_sel[18]),
		.A2(I18[27]),
		.B1(out_sel[19]),
		.B2(I19[27]),
		.Z(O9[27])
	);
	AO_CELL inst_10_27(
		.A1(out_sel[20]),
		.A2(I20[27]),
		.B1(out_sel[21]),
		.B2(I21[27]),
		.Z(O10[27])
	);
	AO_CELL inst_11_27(
		.A1(out_sel[22]),
		.A2(I22[27]),
		.B1(out_sel[23]),
		.B2(I23[27]),
		.Z(O11[27])
	);
	AO_CELL inst_12_27(
		.A1(out_sel[24]),
		.A2(I24[27]),
		.B1(out_sel[25]),
		.B2(I25[27]),
		.Z(O12[27])
	);
	AO_CELL inst_13_27(
		.A1(out_sel[26]),
		.A2(I26[27]),
		.B1(out_sel[27]),
		.B2(I27[27]),
		.Z(O13[27])
	);
	AO_CELL inst_14_27(
		.A1(out_sel[28]),
		.A2(I28[27]),
		.B1(out_sel[29]),
		.B2(I29[27]),
		.Z(O14[27])
	);
	AO_CELL inst_15_27(
		.A1(out_sel[30]),
		.A2(I30[27]),
		.B1(out_sel[31]),
		.B2(I31[27]),
		.Z(O15[27])
	);
	AO_CELL inst_16_27(
		.A1(out_sel[32]),
		.A2(I32[27]),
		.B1(out_sel[33]),
		.B2(I33[27]),
		.Z(O16[27])
	);
	AO_CELL inst_17_27(
		.A1(out_sel[34]),
		.A2(I34[27]),
		.B1(out_sel[35]),
		.B2(I35[27]),
		.Z(O17[27])
	);
	AO_CELL inst_18_27(
		.A1(out_sel[36]),
		.A2(I36[27]),
		.B1(out_sel[37]),
		.B2(I37[27]),
		.Z(O18[27])
	);
	AO_CELL inst_19_27(
		.A1(out_sel[38]),
		.A2(I38[27]),
		.B1(out_sel[39]),
		.B2(I39[27]),
		.Z(O19[27])
	);
	AO_CELL inst_20_27(
		.A1(out_sel[40]),
		.A2(I40[27]),
		.B1(out_sel[41]),
		.B2(I41[27]),
		.Z(O20[27])
	);
	AO_CELL inst_21_27(
		.A1(out_sel[42]),
		.A2(I42[27]),
		.B1(out_sel[43]),
		.B2(I43[27]),
		.Z(O21[27])
	);
	AO_CELL inst_22_27(
		.A1(out_sel[44]),
		.A2(I44[27]),
		.B1(out_sel[45]),
		.B2(I45[27]),
		.Z(O22[27])
	);
	AN_CELL inst_and_27(
		.A1(out_sel[46]),
		.A2(I46[27]),
		.Z(O23[27])
	);
	AO_CELL inst_0_28(
		.A1(out_sel[0]),
		.A2(I0[28]),
		.B1(out_sel[1]),
		.B2(I1[28]),
		.Z(O0[28])
	);
	AO_CELL inst_1_28(
		.A1(out_sel[2]),
		.A2(I2[28]),
		.B1(out_sel[3]),
		.B2(I3[28]),
		.Z(O1[28])
	);
	AO_CELL inst_2_28(
		.A1(out_sel[4]),
		.A2(I4[28]),
		.B1(out_sel[5]),
		.B2(I5[28]),
		.Z(O2[28])
	);
	AO_CELL inst_3_28(
		.A1(out_sel[6]),
		.A2(I6[28]),
		.B1(out_sel[7]),
		.B2(I7[28]),
		.Z(O3[28])
	);
	AO_CELL inst_4_28(
		.A1(out_sel[8]),
		.A2(I8[28]),
		.B1(out_sel[9]),
		.B2(I9[28]),
		.Z(O4[28])
	);
	AO_CELL inst_5_28(
		.A1(out_sel[10]),
		.A2(I10[28]),
		.B1(out_sel[11]),
		.B2(I11[28]),
		.Z(O5[28])
	);
	AO_CELL inst_6_28(
		.A1(out_sel[12]),
		.A2(I12[28]),
		.B1(out_sel[13]),
		.B2(I13[28]),
		.Z(O6[28])
	);
	AO_CELL inst_7_28(
		.A1(out_sel[14]),
		.A2(I14[28]),
		.B1(out_sel[15]),
		.B2(I15[28]),
		.Z(O7[28])
	);
	AO_CELL inst_8_28(
		.A1(out_sel[16]),
		.A2(I16[28]),
		.B1(out_sel[17]),
		.B2(I17[28]),
		.Z(O8[28])
	);
	AO_CELL inst_9_28(
		.A1(out_sel[18]),
		.A2(I18[28]),
		.B1(out_sel[19]),
		.B2(I19[28]),
		.Z(O9[28])
	);
	AO_CELL inst_10_28(
		.A1(out_sel[20]),
		.A2(I20[28]),
		.B1(out_sel[21]),
		.B2(I21[28]),
		.Z(O10[28])
	);
	AO_CELL inst_11_28(
		.A1(out_sel[22]),
		.A2(I22[28]),
		.B1(out_sel[23]),
		.B2(I23[28]),
		.Z(O11[28])
	);
	AO_CELL inst_12_28(
		.A1(out_sel[24]),
		.A2(I24[28]),
		.B1(out_sel[25]),
		.B2(I25[28]),
		.Z(O12[28])
	);
	AO_CELL inst_13_28(
		.A1(out_sel[26]),
		.A2(I26[28]),
		.B1(out_sel[27]),
		.B2(I27[28]),
		.Z(O13[28])
	);
	AO_CELL inst_14_28(
		.A1(out_sel[28]),
		.A2(I28[28]),
		.B1(out_sel[29]),
		.B2(I29[28]),
		.Z(O14[28])
	);
	AO_CELL inst_15_28(
		.A1(out_sel[30]),
		.A2(I30[28]),
		.B1(out_sel[31]),
		.B2(I31[28]),
		.Z(O15[28])
	);
	AO_CELL inst_16_28(
		.A1(out_sel[32]),
		.A2(I32[28]),
		.B1(out_sel[33]),
		.B2(I33[28]),
		.Z(O16[28])
	);
	AO_CELL inst_17_28(
		.A1(out_sel[34]),
		.A2(I34[28]),
		.B1(out_sel[35]),
		.B2(I35[28]),
		.Z(O17[28])
	);
	AO_CELL inst_18_28(
		.A1(out_sel[36]),
		.A2(I36[28]),
		.B1(out_sel[37]),
		.B2(I37[28]),
		.Z(O18[28])
	);
	AO_CELL inst_19_28(
		.A1(out_sel[38]),
		.A2(I38[28]),
		.B1(out_sel[39]),
		.B2(I39[28]),
		.Z(O19[28])
	);
	AO_CELL inst_20_28(
		.A1(out_sel[40]),
		.A2(I40[28]),
		.B1(out_sel[41]),
		.B2(I41[28]),
		.Z(O20[28])
	);
	AO_CELL inst_21_28(
		.A1(out_sel[42]),
		.A2(I42[28]),
		.B1(out_sel[43]),
		.B2(I43[28]),
		.Z(O21[28])
	);
	AO_CELL inst_22_28(
		.A1(out_sel[44]),
		.A2(I44[28]),
		.B1(out_sel[45]),
		.B2(I45[28]),
		.Z(O22[28])
	);
	AN_CELL inst_and_28(
		.A1(out_sel[46]),
		.A2(I46[28]),
		.Z(O23[28])
	);
	AO_CELL inst_0_29(
		.A1(out_sel[0]),
		.A2(I0[29]),
		.B1(out_sel[1]),
		.B2(I1[29]),
		.Z(O0[29])
	);
	AO_CELL inst_1_29(
		.A1(out_sel[2]),
		.A2(I2[29]),
		.B1(out_sel[3]),
		.B2(I3[29]),
		.Z(O1[29])
	);
	AO_CELL inst_2_29(
		.A1(out_sel[4]),
		.A2(I4[29]),
		.B1(out_sel[5]),
		.B2(I5[29]),
		.Z(O2[29])
	);
	AO_CELL inst_3_29(
		.A1(out_sel[6]),
		.A2(I6[29]),
		.B1(out_sel[7]),
		.B2(I7[29]),
		.Z(O3[29])
	);
	AO_CELL inst_4_29(
		.A1(out_sel[8]),
		.A2(I8[29]),
		.B1(out_sel[9]),
		.B2(I9[29]),
		.Z(O4[29])
	);
	AO_CELL inst_5_29(
		.A1(out_sel[10]),
		.A2(I10[29]),
		.B1(out_sel[11]),
		.B2(I11[29]),
		.Z(O5[29])
	);
	AO_CELL inst_6_29(
		.A1(out_sel[12]),
		.A2(I12[29]),
		.B1(out_sel[13]),
		.B2(I13[29]),
		.Z(O6[29])
	);
	AO_CELL inst_7_29(
		.A1(out_sel[14]),
		.A2(I14[29]),
		.B1(out_sel[15]),
		.B2(I15[29]),
		.Z(O7[29])
	);
	AO_CELL inst_8_29(
		.A1(out_sel[16]),
		.A2(I16[29]),
		.B1(out_sel[17]),
		.B2(I17[29]),
		.Z(O8[29])
	);
	AO_CELL inst_9_29(
		.A1(out_sel[18]),
		.A2(I18[29]),
		.B1(out_sel[19]),
		.B2(I19[29]),
		.Z(O9[29])
	);
	AO_CELL inst_10_29(
		.A1(out_sel[20]),
		.A2(I20[29]),
		.B1(out_sel[21]),
		.B2(I21[29]),
		.Z(O10[29])
	);
	AO_CELL inst_11_29(
		.A1(out_sel[22]),
		.A2(I22[29]),
		.B1(out_sel[23]),
		.B2(I23[29]),
		.Z(O11[29])
	);
	AO_CELL inst_12_29(
		.A1(out_sel[24]),
		.A2(I24[29]),
		.B1(out_sel[25]),
		.B2(I25[29]),
		.Z(O12[29])
	);
	AO_CELL inst_13_29(
		.A1(out_sel[26]),
		.A2(I26[29]),
		.B1(out_sel[27]),
		.B2(I27[29]),
		.Z(O13[29])
	);
	AO_CELL inst_14_29(
		.A1(out_sel[28]),
		.A2(I28[29]),
		.B1(out_sel[29]),
		.B2(I29[29]),
		.Z(O14[29])
	);
	AO_CELL inst_15_29(
		.A1(out_sel[30]),
		.A2(I30[29]),
		.B1(out_sel[31]),
		.B2(I31[29]),
		.Z(O15[29])
	);
	AO_CELL inst_16_29(
		.A1(out_sel[32]),
		.A2(I32[29]),
		.B1(out_sel[33]),
		.B2(I33[29]),
		.Z(O16[29])
	);
	AO_CELL inst_17_29(
		.A1(out_sel[34]),
		.A2(I34[29]),
		.B1(out_sel[35]),
		.B2(I35[29]),
		.Z(O17[29])
	);
	AO_CELL inst_18_29(
		.A1(out_sel[36]),
		.A2(I36[29]),
		.B1(out_sel[37]),
		.B2(I37[29]),
		.Z(O18[29])
	);
	AO_CELL inst_19_29(
		.A1(out_sel[38]),
		.A2(I38[29]),
		.B1(out_sel[39]),
		.B2(I39[29]),
		.Z(O19[29])
	);
	AO_CELL inst_20_29(
		.A1(out_sel[40]),
		.A2(I40[29]),
		.B1(out_sel[41]),
		.B2(I41[29]),
		.Z(O20[29])
	);
	AO_CELL inst_21_29(
		.A1(out_sel[42]),
		.A2(I42[29]),
		.B1(out_sel[43]),
		.B2(I43[29]),
		.Z(O21[29])
	);
	AO_CELL inst_22_29(
		.A1(out_sel[44]),
		.A2(I44[29]),
		.B1(out_sel[45]),
		.B2(I45[29]),
		.Z(O22[29])
	);
	AN_CELL inst_and_29(
		.A1(out_sel[46]),
		.A2(I46[29]),
		.Z(O23[29])
	);
	AO_CELL inst_0_30(
		.A1(out_sel[0]),
		.A2(I0[30]),
		.B1(out_sel[1]),
		.B2(I1[30]),
		.Z(O0[30])
	);
	AO_CELL inst_1_30(
		.A1(out_sel[2]),
		.A2(I2[30]),
		.B1(out_sel[3]),
		.B2(I3[30]),
		.Z(O1[30])
	);
	AO_CELL inst_2_30(
		.A1(out_sel[4]),
		.A2(I4[30]),
		.B1(out_sel[5]),
		.B2(I5[30]),
		.Z(O2[30])
	);
	AO_CELL inst_3_30(
		.A1(out_sel[6]),
		.A2(I6[30]),
		.B1(out_sel[7]),
		.B2(I7[30]),
		.Z(O3[30])
	);
	AO_CELL inst_4_30(
		.A1(out_sel[8]),
		.A2(I8[30]),
		.B1(out_sel[9]),
		.B2(I9[30]),
		.Z(O4[30])
	);
	AO_CELL inst_5_30(
		.A1(out_sel[10]),
		.A2(I10[30]),
		.B1(out_sel[11]),
		.B2(I11[30]),
		.Z(O5[30])
	);
	AO_CELL inst_6_30(
		.A1(out_sel[12]),
		.A2(I12[30]),
		.B1(out_sel[13]),
		.B2(I13[30]),
		.Z(O6[30])
	);
	AO_CELL inst_7_30(
		.A1(out_sel[14]),
		.A2(I14[30]),
		.B1(out_sel[15]),
		.B2(I15[30]),
		.Z(O7[30])
	);
	AO_CELL inst_8_30(
		.A1(out_sel[16]),
		.A2(I16[30]),
		.B1(out_sel[17]),
		.B2(I17[30]),
		.Z(O8[30])
	);
	AO_CELL inst_9_30(
		.A1(out_sel[18]),
		.A2(I18[30]),
		.B1(out_sel[19]),
		.B2(I19[30]),
		.Z(O9[30])
	);
	AO_CELL inst_10_30(
		.A1(out_sel[20]),
		.A2(I20[30]),
		.B1(out_sel[21]),
		.B2(I21[30]),
		.Z(O10[30])
	);
	AO_CELL inst_11_30(
		.A1(out_sel[22]),
		.A2(I22[30]),
		.B1(out_sel[23]),
		.B2(I23[30]),
		.Z(O11[30])
	);
	AO_CELL inst_12_30(
		.A1(out_sel[24]),
		.A2(I24[30]),
		.B1(out_sel[25]),
		.B2(I25[30]),
		.Z(O12[30])
	);
	AO_CELL inst_13_30(
		.A1(out_sel[26]),
		.A2(I26[30]),
		.B1(out_sel[27]),
		.B2(I27[30]),
		.Z(O13[30])
	);
	AO_CELL inst_14_30(
		.A1(out_sel[28]),
		.A2(I28[30]),
		.B1(out_sel[29]),
		.B2(I29[30]),
		.Z(O14[30])
	);
	AO_CELL inst_15_30(
		.A1(out_sel[30]),
		.A2(I30[30]),
		.B1(out_sel[31]),
		.B2(I31[30]),
		.Z(O15[30])
	);
	AO_CELL inst_16_30(
		.A1(out_sel[32]),
		.A2(I32[30]),
		.B1(out_sel[33]),
		.B2(I33[30]),
		.Z(O16[30])
	);
	AO_CELL inst_17_30(
		.A1(out_sel[34]),
		.A2(I34[30]),
		.B1(out_sel[35]),
		.B2(I35[30]),
		.Z(O17[30])
	);
	AO_CELL inst_18_30(
		.A1(out_sel[36]),
		.A2(I36[30]),
		.B1(out_sel[37]),
		.B2(I37[30]),
		.Z(O18[30])
	);
	AO_CELL inst_19_30(
		.A1(out_sel[38]),
		.A2(I38[30]),
		.B1(out_sel[39]),
		.B2(I39[30]),
		.Z(O19[30])
	);
	AO_CELL inst_20_30(
		.A1(out_sel[40]),
		.A2(I40[30]),
		.B1(out_sel[41]),
		.B2(I41[30]),
		.Z(O20[30])
	);
	AO_CELL inst_21_30(
		.A1(out_sel[42]),
		.A2(I42[30]),
		.B1(out_sel[43]),
		.B2(I43[30]),
		.Z(O21[30])
	);
	AO_CELL inst_22_30(
		.A1(out_sel[44]),
		.A2(I44[30]),
		.B1(out_sel[45]),
		.B2(I45[30]),
		.Z(O22[30])
	);
	AN_CELL inst_and_30(
		.A1(out_sel[46]),
		.A2(I46[30]),
		.Z(O23[30])
	);
	AO_CELL inst_0_31(
		.A1(out_sel[0]),
		.A2(I0[31]),
		.B1(out_sel[1]),
		.B2(I1[31]),
		.Z(O0[31])
	);
	AO_CELL inst_1_31(
		.A1(out_sel[2]),
		.A2(I2[31]),
		.B1(out_sel[3]),
		.B2(I3[31]),
		.Z(O1[31])
	);
	AO_CELL inst_2_31(
		.A1(out_sel[4]),
		.A2(I4[31]),
		.B1(out_sel[5]),
		.B2(I5[31]),
		.Z(O2[31])
	);
	AO_CELL inst_3_31(
		.A1(out_sel[6]),
		.A2(I6[31]),
		.B1(out_sel[7]),
		.B2(I7[31]),
		.Z(O3[31])
	);
	AO_CELL inst_4_31(
		.A1(out_sel[8]),
		.A2(I8[31]),
		.B1(out_sel[9]),
		.B2(I9[31]),
		.Z(O4[31])
	);
	AO_CELL inst_5_31(
		.A1(out_sel[10]),
		.A2(I10[31]),
		.B1(out_sel[11]),
		.B2(I11[31]),
		.Z(O5[31])
	);
	AO_CELL inst_6_31(
		.A1(out_sel[12]),
		.A2(I12[31]),
		.B1(out_sel[13]),
		.B2(I13[31]),
		.Z(O6[31])
	);
	AO_CELL inst_7_31(
		.A1(out_sel[14]),
		.A2(I14[31]),
		.B1(out_sel[15]),
		.B2(I15[31]),
		.Z(O7[31])
	);
	AO_CELL inst_8_31(
		.A1(out_sel[16]),
		.A2(I16[31]),
		.B1(out_sel[17]),
		.B2(I17[31]),
		.Z(O8[31])
	);
	AO_CELL inst_9_31(
		.A1(out_sel[18]),
		.A2(I18[31]),
		.B1(out_sel[19]),
		.B2(I19[31]),
		.Z(O9[31])
	);
	AO_CELL inst_10_31(
		.A1(out_sel[20]),
		.A2(I20[31]),
		.B1(out_sel[21]),
		.B2(I21[31]),
		.Z(O10[31])
	);
	AO_CELL inst_11_31(
		.A1(out_sel[22]),
		.A2(I22[31]),
		.B1(out_sel[23]),
		.B2(I23[31]),
		.Z(O11[31])
	);
	AO_CELL inst_12_31(
		.A1(out_sel[24]),
		.A2(I24[31]),
		.B1(out_sel[25]),
		.B2(I25[31]),
		.Z(O12[31])
	);
	AO_CELL inst_13_31(
		.A1(out_sel[26]),
		.A2(I26[31]),
		.B1(out_sel[27]),
		.B2(I27[31]),
		.Z(O13[31])
	);
	AO_CELL inst_14_31(
		.A1(out_sel[28]),
		.A2(I28[31]),
		.B1(out_sel[29]),
		.B2(I29[31]),
		.Z(O14[31])
	);
	AO_CELL inst_15_31(
		.A1(out_sel[30]),
		.A2(I30[31]),
		.B1(out_sel[31]),
		.B2(I31[31]),
		.Z(O15[31])
	);
	AO_CELL inst_16_31(
		.A1(out_sel[32]),
		.A2(I32[31]),
		.B1(out_sel[33]),
		.B2(I33[31]),
		.Z(O16[31])
	);
	AO_CELL inst_17_31(
		.A1(out_sel[34]),
		.A2(I34[31]),
		.B1(out_sel[35]),
		.B2(I35[31]),
		.Z(O17[31])
	);
	AO_CELL inst_18_31(
		.A1(out_sel[36]),
		.A2(I36[31]),
		.B1(out_sel[37]),
		.B2(I37[31]),
		.Z(O18[31])
	);
	AO_CELL inst_19_31(
		.A1(out_sel[38]),
		.A2(I38[31]),
		.B1(out_sel[39]),
		.B2(I39[31]),
		.Z(O19[31])
	);
	AO_CELL inst_20_31(
		.A1(out_sel[40]),
		.A2(I40[31]),
		.B1(out_sel[41]),
		.B2(I41[31]),
		.Z(O20[31])
	);
	AO_CELL inst_21_31(
		.A1(out_sel[42]),
		.A2(I42[31]),
		.B1(out_sel[43]),
		.B2(I43[31]),
		.Z(O21[31])
	);
	AO_CELL inst_22_31(
		.A1(out_sel[44]),
		.A2(I44[31]),
		.B1(out_sel[45]),
		.B2(I45[31]),
		.Z(O22[31])
	);
	AN_CELL inst_and_31(
		.A1(out_sel[46]),
		.A2(I46[31]),
		.Z(O23[31])
	);
endmodule
module mux_aoi_2_32 (
	I,
	S,
	out_sel,
	O
);
	input wire [63:0] I;
	input wire S;
	output wire [1:0] out_sel;
	output wire [31:0] O;
	wire [31:0] O_int0;
	precoder_32_2 u_precoder(
		.S(S),
		.out_sel(out_sel)
	);
	mux_logic_32_2 u_mux_logic(
		.I0(I[0+:32]),
		.I1(I[32+:32]),
		.out_sel(out_sel),
		.O0(O_int0)
	);
	assign O = O_int0;
endmodule
module precoder_32_2 (
	S,
	out_sel
);
	input wire [0:0] S;
	output reg [1:0] out_sel;
	always @(*) begin : mux_sel
		case (S)
			1'd0: out_sel = 2'b01;
			1'd1: out_sel = 2'b10;
			default: out_sel = 2'b00;
		endcase
	end
endmodule
module mux_logic_32_2 (
	out_sel,
	I0,
	I1,
	O0
);
	input wire [1:0] out_sel;
	input wire [31:0] I0;
	input wire [31:0] I1;
	output wire [31:0] O0;
	AO_CELL inst_0_0(
		.A1(out_sel[0]),
		.A2(I0[0]),
		.B1(out_sel[1]),
		.B2(I1[0]),
		.Z(O0[0])
	);
	AO_CELL inst_0_1(
		.A1(out_sel[0]),
		.A2(I0[1]),
		.B1(out_sel[1]),
		.B2(I1[1]),
		.Z(O0[1])
	);
	AO_CELL inst_0_2(
		.A1(out_sel[0]),
		.A2(I0[2]),
		.B1(out_sel[1]),
		.B2(I1[2]),
		.Z(O0[2])
	);
	AO_CELL inst_0_3(
		.A1(out_sel[0]),
		.A2(I0[3]),
		.B1(out_sel[1]),
		.B2(I1[3]),
		.Z(O0[3])
	);
	AO_CELL inst_0_4(
		.A1(out_sel[0]),
		.A2(I0[4]),
		.B1(out_sel[1]),
		.B2(I1[4]),
		.Z(O0[4])
	);
	AO_CELL inst_0_5(
		.A1(out_sel[0]),
		.A2(I0[5]),
		.B1(out_sel[1]),
		.B2(I1[5]),
		.Z(O0[5])
	);
	AO_CELL inst_0_6(
		.A1(out_sel[0]),
		.A2(I0[6]),
		.B1(out_sel[1]),
		.B2(I1[6]),
		.Z(O0[6])
	);
	AO_CELL inst_0_7(
		.A1(out_sel[0]),
		.A2(I0[7]),
		.B1(out_sel[1]),
		.B2(I1[7]),
		.Z(O0[7])
	);
	AO_CELL inst_0_8(
		.A1(out_sel[0]),
		.A2(I0[8]),
		.B1(out_sel[1]),
		.B2(I1[8]),
		.Z(O0[8])
	);
	AO_CELL inst_0_9(
		.A1(out_sel[0]),
		.A2(I0[9]),
		.B1(out_sel[1]),
		.B2(I1[9]),
		.Z(O0[9])
	);
	AO_CELL inst_0_10(
		.A1(out_sel[0]),
		.A2(I0[10]),
		.B1(out_sel[1]),
		.B2(I1[10]),
		.Z(O0[10])
	);
	AO_CELL inst_0_11(
		.A1(out_sel[0]),
		.A2(I0[11]),
		.B1(out_sel[1]),
		.B2(I1[11]),
		.Z(O0[11])
	);
	AO_CELL inst_0_12(
		.A1(out_sel[0]),
		.A2(I0[12]),
		.B1(out_sel[1]),
		.B2(I1[12]),
		.Z(O0[12])
	);
	AO_CELL inst_0_13(
		.A1(out_sel[0]),
		.A2(I0[13]),
		.B1(out_sel[1]),
		.B2(I1[13]),
		.Z(O0[13])
	);
	AO_CELL inst_0_14(
		.A1(out_sel[0]),
		.A2(I0[14]),
		.B1(out_sel[1]),
		.B2(I1[14]),
		.Z(O0[14])
	);
	AO_CELL inst_0_15(
		.A1(out_sel[0]),
		.A2(I0[15]),
		.B1(out_sel[1]),
		.B2(I1[15]),
		.Z(O0[15])
	);
	AO_CELL inst_0_16(
		.A1(out_sel[0]),
		.A2(I0[16]),
		.B1(out_sel[1]),
		.B2(I1[16]),
		.Z(O0[16])
	);
	AO_CELL inst_0_17(
		.A1(out_sel[0]),
		.A2(I0[17]),
		.B1(out_sel[1]),
		.B2(I1[17]),
		.Z(O0[17])
	);
	AO_CELL inst_0_18(
		.A1(out_sel[0]),
		.A2(I0[18]),
		.B1(out_sel[1]),
		.B2(I1[18]),
		.Z(O0[18])
	);
	AO_CELL inst_0_19(
		.A1(out_sel[0]),
		.A2(I0[19]),
		.B1(out_sel[1]),
		.B2(I1[19]),
		.Z(O0[19])
	);
	AO_CELL inst_0_20(
		.A1(out_sel[0]),
		.A2(I0[20]),
		.B1(out_sel[1]),
		.B2(I1[20]),
		.Z(O0[20])
	);
	AO_CELL inst_0_21(
		.A1(out_sel[0]),
		.A2(I0[21]),
		.B1(out_sel[1]),
		.B2(I1[21]),
		.Z(O0[21])
	);
	AO_CELL inst_0_22(
		.A1(out_sel[0]),
		.A2(I0[22]),
		.B1(out_sel[1]),
		.B2(I1[22]),
		.Z(O0[22])
	);
	AO_CELL inst_0_23(
		.A1(out_sel[0]),
		.A2(I0[23]),
		.B1(out_sel[1]),
		.B2(I1[23]),
		.Z(O0[23])
	);
	AO_CELL inst_0_24(
		.A1(out_sel[0]),
		.A2(I0[24]),
		.B1(out_sel[1]),
		.B2(I1[24]),
		.Z(O0[24])
	);
	AO_CELL inst_0_25(
		.A1(out_sel[0]),
		.A2(I0[25]),
		.B1(out_sel[1]),
		.B2(I1[25]),
		.Z(O0[25])
	);
	AO_CELL inst_0_26(
		.A1(out_sel[0]),
		.A2(I0[26]),
		.B1(out_sel[1]),
		.B2(I1[26]),
		.Z(O0[26])
	);
	AO_CELL inst_0_27(
		.A1(out_sel[0]),
		.A2(I0[27]),
		.B1(out_sel[1]),
		.B2(I1[27]),
		.Z(O0[27])
	);
	AO_CELL inst_0_28(
		.A1(out_sel[0]),
		.A2(I0[28]),
		.B1(out_sel[1]),
		.B2(I1[28]),
		.Z(O0[28])
	);
	AO_CELL inst_0_29(
		.A1(out_sel[0]),
		.A2(I0[29]),
		.B1(out_sel[1]),
		.B2(I1[29]),
		.Z(O0[29])
	);
	AO_CELL inst_0_30(
		.A1(out_sel[0]),
		.A2(I0[30]),
		.B1(out_sel[1]),
		.B2(I1[30]),
		.Z(O0[30])
	);
	AO_CELL inst_0_31(
		.A1(out_sel[0]),
		.A2(I0[31]),
		.B1(out_sel[1]),
		.B2(I1[31]),
		.Z(O0[31])
	);
endmodule
module mux_aoi_18_32 (
	I,
	S,
	out_sel,
	O
);
	input wire [575:0] I;
	input wire [4:0] S;
	output wire [31:0] out_sel;
	output wire [31:0] O;
	wire [31:0] O_int0;
	wire [31:0] O_int1;
	wire [31:0] O_int2;
	wire [31:0] O_int3;
	wire [31:0] O_int4;
	wire [31:0] O_int5;
	wire [31:0] O_int6;
	wire [31:0] O_int7;
	wire [31:0] O_int8;
	precoder_32_18 u_precoder(
		.S(S),
		.out_sel(out_sel)
	);
	mux_logic_32_18 u_mux_logic(
		.I0(I[0+:32]),
		.I1(I[32+:32]),
		.I2(I[64+:32]),
		.I3(I[96+:32]),
		.I4(I[128+:32]),
		.I5(I[160+:32]),
		.I6(I[192+:32]),
		.I7(I[224+:32]),
		.I8(I[256+:32]),
		.I9(I[288+:32]),
		.I10(I[320+:32]),
		.I11(I[352+:32]),
		.I12(I[384+:32]),
		.I13(I[416+:32]),
		.I14(I[448+:32]),
		.I15(I[480+:32]),
		.I16(I[512+:32]),
		.I17(I[544+:32]),
		.out_sel(out_sel),
		.O0(O_int0),
		.O1(O_int1),
		.O2(O_int2),
		.O3(O_int3),
		.O4(O_int4),
		.O5(O_int5),
		.O6(O_int6),
		.O7(O_int7),
		.O8(O_int8)
	);
	assign O = (((((((O_int0 | O_int1) | O_int2) | O_int3) | O_int4) | O_int5) | O_int6) | O_int7) | O_int8;
endmodule
module precoder_32_18 (
	S,
	out_sel
);
	input wire [4:0] S;
	output reg [31:0] out_sel;
	always @(*) begin : mux_sel
		case (S)
			5'd0: out_sel = 32'b00000000000000000000000000000001;
			5'd1: out_sel = 32'b00000000000000000000000000000010;
			5'd2: out_sel = 32'b00000000000000000000000000000100;
			5'd3: out_sel = 32'b00000000000000000000000000001000;
			5'd4: out_sel = 32'b00000000000000000000000000010000;
			5'd5: out_sel = 32'b00000000000000000000000000100000;
			5'd6: out_sel = 32'b00000000000000000000000001000000;
			5'd7: out_sel = 32'b00000000000000000000000010000000;
			5'd8: out_sel = 32'b00000000000000000000000100000000;
			5'd9: out_sel = 32'b00000000000000000000001000000000;
			5'd10: out_sel = 32'b00000000000000000000010000000000;
			5'd11: out_sel = 32'b00000000000000000000100000000000;
			5'd12: out_sel = 32'b00000000000000000001000000000000;
			5'd13: out_sel = 32'b00000000000000000010000000000000;
			5'd14: out_sel = 32'b00000000000000000100000000000000;
			5'd15: out_sel = 32'b00000000000000001000000000000000;
			5'd16: out_sel = 32'b00000000000000010000000000000000;
			5'd17: out_sel = 32'b00000000000000100000000000000000;
			default: out_sel = 32'b00000000000000000000000000000000;
		endcase
	end
endmodule
module mux_logic_32_18 (
	out_sel,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	I9,
	I10,
	I11,
	I12,
	I13,
	I14,
	I15,
	I16,
	I17,
	O0,
	O1,
	O2,
	O3,
	O4,
	O5,
	O6,
	O7,
	O8
);
	input wire [31:0] out_sel;
	input wire [31:0] I0;
	input wire [31:0] I1;
	input wire [31:0] I2;
	input wire [31:0] I3;
	input wire [31:0] I4;
	input wire [31:0] I5;
	input wire [31:0] I6;
	input wire [31:0] I7;
	input wire [31:0] I8;
	input wire [31:0] I9;
	input wire [31:0] I10;
	input wire [31:0] I11;
	input wire [31:0] I12;
	input wire [31:0] I13;
	input wire [31:0] I14;
	input wire [31:0] I15;
	input wire [31:0] I16;
	input wire [31:0] I17;
	output wire [31:0] O0;
	output wire [31:0] O1;
	output wire [31:0] O2;
	output wire [31:0] O3;
	output wire [31:0] O4;
	output wire [31:0] O5;
	output wire [31:0] O6;
	output wire [31:0] O7;
	output wire [31:0] O8;
	AO_CELL inst_0_0(
		.A1(out_sel[0]),
		.A2(I0[0]),
		.B1(out_sel[1]),
		.B2(I1[0]),
		.Z(O0[0])
	);
	AO_CELL inst_1_0(
		.A1(out_sel[2]),
		.A2(I2[0]),
		.B1(out_sel[3]),
		.B2(I3[0]),
		.Z(O1[0])
	);
	AO_CELL inst_2_0(
		.A1(out_sel[4]),
		.A2(I4[0]),
		.B1(out_sel[5]),
		.B2(I5[0]),
		.Z(O2[0])
	);
	AO_CELL inst_3_0(
		.A1(out_sel[6]),
		.A2(I6[0]),
		.B1(out_sel[7]),
		.B2(I7[0]),
		.Z(O3[0])
	);
	AO_CELL inst_4_0(
		.A1(out_sel[8]),
		.A2(I8[0]),
		.B1(out_sel[9]),
		.B2(I9[0]),
		.Z(O4[0])
	);
	AO_CELL inst_5_0(
		.A1(out_sel[10]),
		.A2(I10[0]),
		.B1(out_sel[11]),
		.B2(I11[0]),
		.Z(O5[0])
	);
	AO_CELL inst_6_0(
		.A1(out_sel[12]),
		.A2(I12[0]),
		.B1(out_sel[13]),
		.B2(I13[0]),
		.Z(O6[0])
	);
	AO_CELL inst_7_0(
		.A1(out_sel[14]),
		.A2(I14[0]),
		.B1(out_sel[15]),
		.B2(I15[0]),
		.Z(O7[0])
	);
	AO_CELL inst_8_0(
		.A1(out_sel[16]),
		.A2(I16[0]),
		.B1(out_sel[17]),
		.B2(I17[0]),
		.Z(O8[0])
	);
	AO_CELL inst_0_1(
		.A1(out_sel[0]),
		.A2(I0[1]),
		.B1(out_sel[1]),
		.B2(I1[1]),
		.Z(O0[1])
	);
	AO_CELL inst_1_1(
		.A1(out_sel[2]),
		.A2(I2[1]),
		.B1(out_sel[3]),
		.B2(I3[1]),
		.Z(O1[1])
	);
	AO_CELL inst_2_1(
		.A1(out_sel[4]),
		.A2(I4[1]),
		.B1(out_sel[5]),
		.B2(I5[1]),
		.Z(O2[1])
	);
	AO_CELL inst_3_1(
		.A1(out_sel[6]),
		.A2(I6[1]),
		.B1(out_sel[7]),
		.B2(I7[1]),
		.Z(O3[1])
	);
	AO_CELL inst_4_1(
		.A1(out_sel[8]),
		.A2(I8[1]),
		.B1(out_sel[9]),
		.B2(I9[1]),
		.Z(O4[1])
	);
	AO_CELL inst_5_1(
		.A1(out_sel[10]),
		.A2(I10[1]),
		.B1(out_sel[11]),
		.B2(I11[1]),
		.Z(O5[1])
	);
	AO_CELL inst_6_1(
		.A1(out_sel[12]),
		.A2(I12[1]),
		.B1(out_sel[13]),
		.B2(I13[1]),
		.Z(O6[1])
	);
	AO_CELL inst_7_1(
		.A1(out_sel[14]),
		.A2(I14[1]),
		.B1(out_sel[15]),
		.B2(I15[1]),
		.Z(O7[1])
	);
	AO_CELL inst_8_1(
		.A1(out_sel[16]),
		.A2(I16[1]),
		.B1(out_sel[17]),
		.B2(I17[1]),
		.Z(O8[1])
	);
	AO_CELL inst_0_2(
		.A1(out_sel[0]),
		.A2(I0[2]),
		.B1(out_sel[1]),
		.B2(I1[2]),
		.Z(O0[2])
	);
	AO_CELL inst_1_2(
		.A1(out_sel[2]),
		.A2(I2[2]),
		.B1(out_sel[3]),
		.B2(I3[2]),
		.Z(O1[2])
	);
	AO_CELL inst_2_2(
		.A1(out_sel[4]),
		.A2(I4[2]),
		.B1(out_sel[5]),
		.B2(I5[2]),
		.Z(O2[2])
	);
	AO_CELL inst_3_2(
		.A1(out_sel[6]),
		.A2(I6[2]),
		.B1(out_sel[7]),
		.B2(I7[2]),
		.Z(O3[2])
	);
	AO_CELL inst_4_2(
		.A1(out_sel[8]),
		.A2(I8[2]),
		.B1(out_sel[9]),
		.B2(I9[2]),
		.Z(O4[2])
	);
	AO_CELL inst_5_2(
		.A1(out_sel[10]),
		.A2(I10[2]),
		.B1(out_sel[11]),
		.B2(I11[2]),
		.Z(O5[2])
	);
	AO_CELL inst_6_2(
		.A1(out_sel[12]),
		.A2(I12[2]),
		.B1(out_sel[13]),
		.B2(I13[2]),
		.Z(O6[2])
	);
	AO_CELL inst_7_2(
		.A1(out_sel[14]),
		.A2(I14[2]),
		.B1(out_sel[15]),
		.B2(I15[2]),
		.Z(O7[2])
	);
	AO_CELL inst_8_2(
		.A1(out_sel[16]),
		.A2(I16[2]),
		.B1(out_sel[17]),
		.B2(I17[2]),
		.Z(O8[2])
	);
	AO_CELL inst_0_3(
		.A1(out_sel[0]),
		.A2(I0[3]),
		.B1(out_sel[1]),
		.B2(I1[3]),
		.Z(O0[3])
	);
	AO_CELL inst_1_3(
		.A1(out_sel[2]),
		.A2(I2[3]),
		.B1(out_sel[3]),
		.B2(I3[3]),
		.Z(O1[3])
	);
	AO_CELL inst_2_3(
		.A1(out_sel[4]),
		.A2(I4[3]),
		.B1(out_sel[5]),
		.B2(I5[3]),
		.Z(O2[3])
	);
	AO_CELL inst_3_3(
		.A1(out_sel[6]),
		.A2(I6[3]),
		.B1(out_sel[7]),
		.B2(I7[3]),
		.Z(O3[3])
	);
	AO_CELL inst_4_3(
		.A1(out_sel[8]),
		.A2(I8[3]),
		.B1(out_sel[9]),
		.B2(I9[3]),
		.Z(O4[3])
	);
	AO_CELL inst_5_3(
		.A1(out_sel[10]),
		.A2(I10[3]),
		.B1(out_sel[11]),
		.B2(I11[3]),
		.Z(O5[3])
	);
	AO_CELL inst_6_3(
		.A1(out_sel[12]),
		.A2(I12[3]),
		.B1(out_sel[13]),
		.B2(I13[3]),
		.Z(O6[3])
	);
	AO_CELL inst_7_3(
		.A1(out_sel[14]),
		.A2(I14[3]),
		.B1(out_sel[15]),
		.B2(I15[3]),
		.Z(O7[3])
	);
	AO_CELL inst_8_3(
		.A1(out_sel[16]),
		.A2(I16[3]),
		.B1(out_sel[17]),
		.B2(I17[3]),
		.Z(O8[3])
	);
	AO_CELL inst_0_4(
		.A1(out_sel[0]),
		.A2(I0[4]),
		.B1(out_sel[1]),
		.B2(I1[4]),
		.Z(O0[4])
	);
	AO_CELL inst_1_4(
		.A1(out_sel[2]),
		.A2(I2[4]),
		.B1(out_sel[3]),
		.B2(I3[4]),
		.Z(O1[4])
	);
	AO_CELL inst_2_4(
		.A1(out_sel[4]),
		.A2(I4[4]),
		.B1(out_sel[5]),
		.B2(I5[4]),
		.Z(O2[4])
	);
	AO_CELL inst_3_4(
		.A1(out_sel[6]),
		.A2(I6[4]),
		.B1(out_sel[7]),
		.B2(I7[4]),
		.Z(O3[4])
	);
	AO_CELL inst_4_4(
		.A1(out_sel[8]),
		.A2(I8[4]),
		.B1(out_sel[9]),
		.B2(I9[4]),
		.Z(O4[4])
	);
	AO_CELL inst_5_4(
		.A1(out_sel[10]),
		.A2(I10[4]),
		.B1(out_sel[11]),
		.B2(I11[4]),
		.Z(O5[4])
	);
	AO_CELL inst_6_4(
		.A1(out_sel[12]),
		.A2(I12[4]),
		.B1(out_sel[13]),
		.B2(I13[4]),
		.Z(O6[4])
	);
	AO_CELL inst_7_4(
		.A1(out_sel[14]),
		.A2(I14[4]),
		.B1(out_sel[15]),
		.B2(I15[4]),
		.Z(O7[4])
	);
	AO_CELL inst_8_4(
		.A1(out_sel[16]),
		.A2(I16[4]),
		.B1(out_sel[17]),
		.B2(I17[4]),
		.Z(O8[4])
	);
	AO_CELL inst_0_5(
		.A1(out_sel[0]),
		.A2(I0[5]),
		.B1(out_sel[1]),
		.B2(I1[5]),
		.Z(O0[5])
	);
	AO_CELL inst_1_5(
		.A1(out_sel[2]),
		.A2(I2[5]),
		.B1(out_sel[3]),
		.B2(I3[5]),
		.Z(O1[5])
	);
	AO_CELL inst_2_5(
		.A1(out_sel[4]),
		.A2(I4[5]),
		.B1(out_sel[5]),
		.B2(I5[5]),
		.Z(O2[5])
	);
	AO_CELL inst_3_5(
		.A1(out_sel[6]),
		.A2(I6[5]),
		.B1(out_sel[7]),
		.B2(I7[5]),
		.Z(O3[5])
	);
	AO_CELL inst_4_5(
		.A1(out_sel[8]),
		.A2(I8[5]),
		.B1(out_sel[9]),
		.B2(I9[5]),
		.Z(O4[5])
	);
	AO_CELL inst_5_5(
		.A1(out_sel[10]),
		.A2(I10[5]),
		.B1(out_sel[11]),
		.B2(I11[5]),
		.Z(O5[5])
	);
	AO_CELL inst_6_5(
		.A1(out_sel[12]),
		.A2(I12[5]),
		.B1(out_sel[13]),
		.B2(I13[5]),
		.Z(O6[5])
	);
	AO_CELL inst_7_5(
		.A1(out_sel[14]),
		.A2(I14[5]),
		.B1(out_sel[15]),
		.B2(I15[5]),
		.Z(O7[5])
	);
	AO_CELL inst_8_5(
		.A1(out_sel[16]),
		.A2(I16[5]),
		.B1(out_sel[17]),
		.B2(I17[5]),
		.Z(O8[5])
	);
	AO_CELL inst_0_6(
		.A1(out_sel[0]),
		.A2(I0[6]),
		.B1(out_sel[1]),
		.B2(I1[6]),
		.Z(O0[6])
	);
	AO_CELL inst_1_6(
		.A1(out_sel[2]),
		.A2(I2[6]),
		.B1(out_sel[3]),
		.B2(I3[6]),
		.Z(O1[6])
	);
	AO_CELL inst_2_6(
		.A1(out_sel[4]),
		.A2(I4[6]),
		.B1(out_sel[5]),
		.B2(I5[6]),
		.Z(O2[6])
	);
	AO_CELL inst_3_6(
		.A1(out_sel[6]),
		.A2(I6[6]),
		.B1(out_sel[7]),
		.B2(I7[6]),
		.Z(O3[6])
	);
	AO_CELL inst_4_6(
		.A1(out_sel[8]),
		.A2(I8[6]),
		.B1(out_sel[9]),
		.B2(I9[6]),
		.Z(O4[6])
	);
	AO_CELL inst_5_6(
		.A1(out_sel[10]),
		.A2(I10[6]),
		.B1(out_sel[11]),
		.B2(I11[6]),
		.Z(O5[6])
	);
	AO_CELL inst_6_6(
		.A1(out_sel[12]),
		.A2(I12[6]),
		.B1(out_sel[13]),
		.B2(I13[6]),
		.Z(O6[6])
	);
	AO_CELL inst_7_6(
		.A1(out_sel[14]),
		.A2(I14[6]),
		.B1(out_sel[15]),
		.B2(I15[6]),
		.Z(O7[6])
	);
	AO_CELL inst_8_6(
		.A1(out_sel[16]),
		.A2(I16[6]),
		.B1(out_sel[17]),
		.B2(I17[6]),
		.Z(O8[6])
	);
	AO_CELL inst_0_7(
		.A1(out_sel[0]),
		.A2(I0[7]),
		.B1(out_sel[1]),
		.B2(I1[7]),
		.Z(O0[7])
	);
	AO_CELL inst_1_7(
		.A1(out_sel[2]),
		.A2(I2[7]),
		.B1(out_sel[3]),
		.B2(I3[7]),
		.Z(O1[7])
	);
	AO_CELL inst_2_7(
		.A1(out_sel[4]),
		.A2(I4[7]),
		.B1(out_sel[5]),
		.B2(I5[7]),
		.Z(O2[7])
	);
	AO_CELL inst_3_7(
		.A1(out_sel[6]),
		.A2(I6[7]),
		.B1(out_sel[7]),
		.B2(I7[7]),
		.Z(O3[7])
	);
	AO_CELL inst_4_7(
		.A1(out_sel[8]),
		.A2(I8[7]),
		.B1(out_sel[9]),
		.B2(I9[7]),
		.Z(O4[7])
	);
	AO_CELL inst_5_7(
		.A1(out_sel[10]),
		.A2(I10[7]),
		.B1(out_sel[11]),
		.B2(I11[7]),
		.Z(O5[7])
	);
	AO_CELL inst_6_7(
		.A1(out_sel[12]),
		.A2(I12[7]),
		.B1(out_sel[13]),
		.B2(I13[7]),
		.Z(O6[7])
	);
	AO_CELL inst_7_7(
		.A1(out_sel[14]),
		.A2(I14[7]),
		.B1(out_sel[15]),
		.B2(I15[7]),
		.Z(O7[7])
	);
	AO_CELL inst_8_7(
		.A1(out_sel[16]),
		.A2(I16[7]),
		.B1(out_sel[17]),
		.B2(I17[7]),
		.Z(O8[7])
	);
	AO_CELL inst_0_8(
		.A1(out_sel[0]),
		.A2(I0[8]),
		.B1(out_sel[1]),
		.B2(I1[8]),
		.Z(O0[8])
	);
	AO_CELL inst_1_8(
		.A1(out_sel[2]),
		.A2(I2[8]),
		.B1(out_sel[3]),
		.B2(I3[8]),
		.Z(O1[8])
	);
	AO_CELL inst_2_8(
		.A1(out_sel[4]),
		.A2(I4[8]),
		.B1(out_sel[5]),
		.B2(I5[8]),
		.Z(O2[8])
	);
	AO_CELL inst_3_8(
		.A1(out_sel[6]),
		.A2(I6[8]),
		.B1(out_sel[7]),
		.B2(I7[8]),
		.Z(O3[8])
	);
	AO_CELL inst_4_8(
		.A1(out_sel[8]),
		.A2(I8[8]),
		.B1(out_sel[9]),
		.B2(I9[8]),
		.Z(O4[8])
	);
	AO_CELL inst_5_8(
		.A1(out_sel[10]),
		.A2(I10[8]),
		.B1(out_sel[11]),
		.B2(I11[8]),
		.Z(O5[8])
	);
	AO_CELL inst_6_8(
		.A1(out_sel[12]),
		.A2(I12[8]),
		.B1(out_sel[13]),
		.B2(I13[8]),
		.Z(O6[8])
	);
	AO_CELL inst_7_8(
		.A1(out_sel[14]),
		.A2(I14[8]),
		.B1(out_sel[15]),
		.B2(I15[8]),
		.Z(O7[8])
	);
	AO_CELL inst_8_8(
		.A1(out_sel[16]),
		.A2(I16[8]),
		.B1(out_sel[17]),
		.B2(I17[8]),
		.Z(O8[8])
	);
	AO_CELL inst_0_9(
		.A1(out_sel[0]),
		.A2(I0[9]),
		.B1(out_sel[1]),
		.B2(I1[9]),
		.Z(O0[9])
	);
	AO_CELL inst_1_9(
		.A1(out_sel[2]),
		.A2(I2[9]),
		.B1(out_sel[3]),
		.B2(I3[9]),
		.Z(O1[9])
	);
	AO_CELL inst_2_9(
		.A1(out_sel[4]),
		.A2(I4[9]),
		.B1(out_sel[5]),
		.B2(I5[9]),
		.Z(O2[9])
	);
	AO_CELL inst_3_9(
		.A1(out_sel[6]),
		.A2(I6[9]),
		.B1(out_sel[7]),
		.B2(I7[9]),
		.Z(O3[9])
	);
	AO_CELL inst_4_9(
		.A1(out_sel[8]),
		.A2(I8[9]),
		.B1(out_sel[9]),
		.B2(I9[9]),
		.Z(O4[9])
	);
	AO_CELL inst_5_9(
		.A1(out_sel[10]),
		.A2(I10[9]),
		.B1(out_sel[11]),
		.B2(I11[9]),
		.Z(O5[9])
	);
	AO_CELL inst_6_9(
		.A1(out_sel[12]),
		.A2(I12[9]),
		.B1(out_sel[13]),
		.B2(I13[9]),
		.Z(O6[9])
	);
	AO_CELL inst_7_9(
		.A1(out_sel[14]),
		.A2(I14[9]),
		.B1(out_sel[15]),
		.B2(I15[9]),
		.Z(O7[9])
	);
	AO_CELL inst_8_9(
		.A1(out_sel[16]),
		.A2(I16[9]),
		.B1(out_sel[17]),
		.B2(I17[9]),
		.Z(O8[9])
	);
	AO_CELL inst_0_10(
		.A1(out_sel[0]),
		.A2(I0[10]),
		.B1(out_sel[1]),
		.B2(I1[10]),
		.Z(O0[10])
	);
	AO_CELL inst_1_10(
		.A1(out_sel[2]),
		.A2(I2[10]),
		.B1(out_sel[3]),
		.B2(I3[10]),
		.Z(O1[10])
	);
	AO_CELL inst_2_10(
		.A1(out_sel[4]),
		.A2(I4[10]),
		.B1(out_sel[5]),
		.B2(I5[10]),
		.Z(O2[10])
	);
	AO_CELL inst_3_10(
		.A1(out_sel[6]),
		.A2(I6[10]),
		.B1(out_sel[7]),
		.B2(I7[10]),
		.Z(O3[10])
	);
	AO_CELL inst_4_10(
		.A1(out_sel[8]),
		.A2(I8[10]),
		.B1(out_sel[9]),
		.B2(I9[10]),
		.Z(O4[10])
	);
	AO_CELL inst_5_10(
		.A1(out_sel[10]),
		.A2(I10[10]),
		.B1(out_sel[11]),
		.B2(I11[10]),
		.Z(O5[10])
	);
	AO_CELL inst_6_10(
		.A1(out_sel[12]),
		.A2(I12[10]),
		.B1(out_sel[13]),
		.B2(I13[10]),
		.Z(O6[10])
	);
	AO_CELL inst_7_10(
		.A1(out_sel[14]),
		.A2(I14[10]),
		.B1(out_sel[15]),
		.B2(I15[10]),
		.Z(O7[10])
	);
	AO_CELL inst_8_10(
		.A1(out_sel[16]),
		.A2(I16[10]),
		.B1(out_sel[17]),
		.B2(I17[10]),
		.Z(O8[10])
	);
	AO_CELL inst_0_11(
		.A1(out_sel[0]),
		.A2(I0[11]),
		.B1(out_sel[1]),
		.B2(I1[11]),
		.Z(O0[11])
	);
	AO_CELL inst_1_11(
		.A1(out_sel[2]),
		.A2(I2[11]),
		.B1(out_sel[3]),
		.B2(I3[11]),
		.Z(O1[11])
	);
	AO_CELL inst_2_11(
		.A1(out_sel[4]),
		.A2(I4[11]),
		.B1(out_sel[5]),
		.B2(I5[11]),
		.Z(O2[11])
	);
	AO_CELL inst_3_11(
		.A1(out_sel[6]),
		.A2(I6[11]),
		.B1(out_sel[7]),
		.B2(I7[11]),
		.Z(O3[11])
	);
	AO_CELL inst_4_11(
		.A1(out_sel[8]),
		.A2(I8[11]),
		.B1(out_sel[9]),
		.B2(I9[11]),
		.Z(O4[11])
	);
	AO_CELL inst_5_11(
		.A1(out_sel[10]),
		.A2(I10[11]),
		.B1(out_sel[11]),
		.B2(I11[11]),
		.Z(O5[11])
	);
	AO_CELL inst_6_11(
		.A1(out_sel[12]),
		.A2(I12[11]),
		.B1(out_sel[13]),
		.B2(I13[11]),
		.Z(O6[11])
	);
	AO_CELL inst_7_11(
		.A1(out_sel[14]),
		.A2(I14[11]),
		.B1(out_sel[15]),
		.B2(I15[11]),
		.Z(O7[11])
	);
	AO_CELL inst_8_11(
		.A1(out_sel[16]),
		.A2(I16[11]),
		.B1(out_sel[17]),
		.B2(I17[11]),
		.Z(O8[11])
	);
	AO_CELL inst_0_12(
		.A1(out_sel[0]),
		.A2(I0[12]),
		.B1(out_sel[1]),
		.B2(I1[12]),
		.Z(O0[12])
	);
	AO_CELL inst_1_12(
		.A1(out_sel[2]),
		.A2(I2[12]),
		.B1(out_sel[3]),
		.B2(I3[12]),
		.Z(O1[12])
	);
	AO_CELL inst_2_12(
		.A1(out_sel[4]),
		.A2(I4[12]),
		.B1(out_sel[5]),
		.B2(I5[12]),
		.Z(O2[12])
	);
	AO_CELL inst_3_12(
		.A1(out_sel[6]),
		.A2(I6[12]),
		.B1(out_sel[7]),
		.B2(I7[12]),
		.Z(O3[12])
	);
	AO_CELL inst_4_12(
		.A1(out_sel[8]),
		.A2(I8[12]),
		.B1(out_sel[9]),
		.B2(I9[12]),
		.Z(O4[12])
	);
	AO_CELL inst_5_12(
		.A1(out_sel[10]),
		.A2(I10[12]),
		.B1(out_sel[11]),
		.B2(I11[12]),
		.Z(O5[12])
	);
	AO_CELL inst_6_12(
		.A1(out_sel[12]),
		.A2(I12[12]),
		.B1(out_sel[13]),
		.B2(I13[12]),
		.Z(O6[12])
	);
	AO_CELL inst_7_12(
		.A1(out_sel[14]),
		.A2(I14[12]),
		.B1(out_sel[15]),
		.B2(I15[12]),
		.Z(O7[12])
	);
	AO_CELL inst_8_12(
		.A1(out_sel[16]),
		.A2(I16[12]),
		.B1(out_sel[17]),
		.B2(I17[12]),
		.Z(O8[12])
	);
	AO_CELL inst_0_13(
		.A1(out_sel[0]),
		.A2(I0[13]),
		.B1(out_sel[1]),
		.B2(I1[13]),
		.Z(O0[13])
	);
	AO_CELL inst_1_13(
		.A1(out_sel[2]),
		.A2(I2[13]),
		.B1(out_sel[3]),
		.B2(I3[13]),
		.Z(O1[13])
	);
	AO_CELL inst_2_13(
		.A1(out_sel[4]),
		.A2(I4[13]),
		.B1(out_sel[5]),
		.B2(I5[13]),
		.Z(O2[13])
	);
	AO_CELL inst_3_13(
		.A1(out_sel[6]),
		.A2(I6[13]),
		.B1(out_sel[7]),
		.B2(I7[13]),
		.Z(O3[13])
	);
	AO_CELL inst_4_13(
		.A1(out_sel[8]),
		.A2(I8[13]),
		.B1(out_sel[9]),
		.B2(I9[13]),
		.Z(O4[13])
	);
	AO_CELL inst_5_13(
		.A1(out_sel[10]),
		.A2(I10[13]),
		.B1(out_sel[11]),
		.B2(I11[13]),
		.Z(O5[13])
	);
	AO_CELL inst_6_13(
		.A1(out_sel[12]),
		.A2(I12[13]),
		.B1(out_sel[13]),
		.B2(I13[13]),
		.Z(O6[13])
	);
	AO_CELL inst_7_13(
		.A1(out_sel[14]),
		.A2(I14[13]),
		.B1(out_sel[15]),
		.B2(I15[13]),
		.Z(O7[13])
	);
	AO_CELL inst_8_13(
		.A1(out_sel[16]),
		.A2(I16[13]),
		.B1(out_sel[17]),
		.B2(I17[13]),
		.Z(O8[13])
	);
	AO_CELL inst_0_14(
		.A1(out_sel[0]),
		.A2(I0[14]),
		.B1(out_sel[1]),
		.B2(I1[14]),
		.Z(O0[14])
	);
	AO_CELL inst_1_14(
		.A1(out_sel[2]),
		.A2(I2[14]),
		.B1(out_sel[3]),
		.B2(I3[14]),
		.Z(O1[14])
	);
	AO_CELL inst_2_14(
		.A1(out_sel[4]),
		.A2(I4[14]),
		.B1(out_sel[5]),
		.B2(I5[14]),
		.Z(O2[14])
	);
	AO_CELL inst_3_14(
		.A1(out_sel[6]),
		.A2(I6[14]),
		.B1(out_sel[7]),
		.B2(I7[14]),
		.Z(O3[14])
	);
	AO_CELL inst_4_14(
		.A1(out_sel[8]),
		.A2(I8[14]),
		.B1(out_sel[9]),
		.B2(I9[14]),
		.Z(O4[14])
	);
	AO_CELL inst_5_14(
		.A1(out_sel[10]),
		.A2(I10[14]),
		.B1(out_sel[11]),
		.B2(I11[14]),
		.Z(O5[14])
	);
	AO_CELL inst_6_14(
		.A1(out_sel[12]),
		.A2(I12[14]),
		.B1(out_sel[13]),
		.B2(I13[14]),
		.Z(O6[14])
	);
	AO_CELL inst_7_14(
		.A1(out_sel[14]),
		.A2(I14[14]),
		.B1(out_sel[15]),
		.B2(I15[14]),
		.Z(O7[14])
	);
	AO_CELL inst_8_14(
		.A1(out_sel[16]),
		.A2(I16[14]),
		.B1(out_sel[17]),
		.B2(I17[14]),
		.Z(O8[14])
	);
	AO_CELL inst_0_15(
		.A1(out_sel[0]),
		.A2(I0[15]),
		.B1(out_sel[1]),
		.B2(I1[15]),
		.Z(O0[15])
	);
	AO_CELL inst_1_15(
		.A1(out_sel[2]),
		.A2(I2[15]),
		.B1(out_sel[3]),
		.B2(I3[15]),
		.Z(O1[15])
	);
	AO_CELL inst_2_15(
		.A1(out_sel[4]),
		.A2(I4[15]),
		.B1(out_sel[5]),
		.B2(I5[15]),
		.Z(O2[15])
	);
	AO_CELL inst_3_15(
		.A1(out_sel[6]),
		.A2(I6[15]),
		.B1(out_sel[7]),
		.B2(I7[15]),
		.Z(O3[15])
	);
	AO_CELL inst_4_15(
		.A1(out_sel[8]),
		.A2(I8[15]),
		.B1(out_sel[9]),
		.B2(I9[15]),
		.Z(O4[15])
	);
	AO_CELL inst_5_15(
		.A1(out_sel[10]),
		.A2(I10[15]),
		.B1(out_sel[11]),
		.B2(I11[15]),
		.Z(O5[15])
	);
	AO_CELL inst_6_15(
		.A1(out_sel[12]),
		.A2(I12[15]),
		.B1(out_sel[13]),
		.B2(I13[15]),
		.Z(O6[15])
	);
	AO_CELL inst_7_15(
		.A1(out_sel[14]),
		.A2(I14[15]),
		.B1(out_sel[15]),
		.B2(I15[15]),
		.Z(O7[15])
	);
	AO_CELL inst_8_15(
		.A1(out_sel[16]),
		.A2(I16[15]),
		.B1(out_sel[17]),
		.B2(I17[15]),
		.Z(O8[15])
	);
	AO_CELL inst_0_16(
		.A1(out_sel[0]),
		.A2(I0[16]),
		.B1(out_sel[1]),
		.B2(I1[16]),
		.Z(O0[16])
	);
	AO_CELL inst_1_16(
		.A1(out_sel[2]),
		.A2(I2[16]),
		.B1(out_sel[3]),
		.B2(I3[16]),
		.Z(O1[16])
	);
	AO_CELL inst_2_16(
		.A1(out_sel[4]),
		.A2(I4[16]),
		.B1(out_sel[5]),
		.B2(I5[16]),
		.Z(O2[16])
	);
	AO_CELL inst_3_16(
		.A1(out_sel[6]),
		.A2(I6[16]),
		.B1(out_sel[7]),
		.B2(I7[16]),
		.Z(O3[16])
	);
	AO_CELL inst_4_16(
		.A1(out_sel[8]),
		.A2(I8[16]),
		.B1(out_sel[9]),
		.B2(I9[16]),
		.Z(O4[16])
	);
	AO_CELL inst_5_16(
		.A1(out_sel[10]),
		.A2(I10[16]),
		.B1(out_sel[11]),
		.B2(I11[16]),
		.Z(O5[16])
	);
	AO_CELL inst_6_16(
		.A1(out_sel[12]),
		.A2(I12[16]),
		.B1(out_sel[13]),
		.B2(I13[16]),
		.Z(O6[16])
	);
	AO_CELL inst_7_16(
		.A1(out_sel[14]),
		.A2(I14[16]),
		.B1(out_sel[15]),
		.B2(I15[16]),
		.Z(O7[16])
	);
	AO_CELL inst_8_16(
		.A1(out_sel[16]),
		.A2(I16[16]),
		.B1(out_sel[17]),
		.B2(I17[16]),
		.Z(O8[16])
	);
	AO_CELL inst_0_17(
		.A1(out_sel[0]),
		.A2(I0[17]),
		.B1(out_sel[1]),
		.B2(I1[17]),
		.Z(O0[17])
	);
	AO_CELL inst_1_17(
		.A1(out_sel[2]),
		.A2(I2[17]),
		.B1(out_sel[3]),
		.B2(I3[17]),
		.Z(O1[17])
	);
	AO_CELL inst_2_17(
		.A1(out_sel[4]),
		.A2(I4[17]),
		.B1(out_sel[5]),
		.B2(I5[17]),
		.Z(O2[17])
	);
	AO_CELL inst_3_17(
		.A1(out_sel[6]),
		.A2(I6[17]),
		.B1(out_sel[7]),
		.B2(I7[17]),
		.Z(O3[17])
	);
	AO_CELL inst_4_17(
		.A1(out_sel[8]),
		.A2(I8[17]),
		.B1(out_sel[9]),
		.B2(I9[17]),
		.Z(O4[17])
	);
	AO_CELL inst_5_17(
		.A1(out_sel[10]),
		.A2(I10[17]),
		.B1(out_sel[11]),
		.B2(I11[17]),
		.Z(O5[17])
	);
	AO_CELL inst_6_17(
		.A1(out_sel[12]),
		.A2(I12[17]),
		.B1(out_sel[13]),
		.B2(I13[17]),
		.Z(O6[17])
	);
	AO_CELL inst_7_17(
		.A1(out_sel[14]),
		.A2(I14[17]),
		.B1(out_sel[15]),
		.B2(I15[17]),
		.Z(O7[17])
	);
	AO_CELL inst_8_17(
		.A1(out_sel[16]),
		.A2(I16[17]),
		.B1(out_sel[17]),
		.B2(I17[17]),
		.Z(O8[17])
	);
	AO_CELL inst_0_18(
		.A1(out_sel[0]),
		.A2(I0[18]),
		.B1(out_sel[1]),
		.B2(I1[18]),
		.Z(O0[18])
	);
	AO_CELL inst_1_18(
		.A1(out_sel[2]),
		.A2(I2[18]),
		.B1(out_sel[3]),
		.B2(I3[18]),
		.Z(O1[18])
	);
	AO_CELL inst_2_18(
		.A1(out_sel[4]),
		.A2(I4[18]),
		.B1(out_sel[5]),
		.B2(I5[18]),
		.Z(O2[18])
	);
	AO_CELL inst_3_18(
		.A1(out_sel[6]),
		.A2(I6[18]),
		.B1(out_sel[7]),
		.B2(I7[18]),
		.Z(O3[18])
	);
	AO_CELL inst_4_18(
		.A1(out_sel[8]),
		.A2(I8[18]),
		.B1(out_sel[9]),
		.B2(I9[18]),
		.Z(O4[18])
	);
	AO_CELL inst_5_18(
		.A1(out_sel[10]),
		.A2(I10[18]),
		.B1(out_sel[11]),
		.B2(I11[18]),
		.Z(O5[18])
	);
	AO_CELL inst_6_18(
		.A1(out_sel[12]),
		.A2(I12[18]),
		.B1(out_sel[13]),
		.B2(I13[18]),
		.Z(O6[18])
	);
	AO_CELL inst_7_18(
		.A1(out_sel[14]),
		.A2(I14[18]),
		.B1(out_sel[15]),
		.B2(I15[18]),
		.Z(O7[18])
	);
	AO_CELL inst_8_18(
		.A1(out_sel[16]),
		.A2(I16[18]),
		.B1(out_sel[17]),
		.B2(I17[18]),
		.Z(O8[18])
	);
	AO_CELL inst_0_19(
		.A1(out_sel[0]),
		.A2(I0[19]),
		.B1(out_sel[1]),
		.B2(I1[19]),
		.Z(O0[19])
	);
	AO_CELL inst_1_19(
		.A1(out_sel[2]),
		.A2(I2[19]),
		.B1(out_sel[3]),
		.B2(I3[19]),
		.Z(O1[19])
	);
	AO_CELL inst_2_19(
		.A1(out_sel[4]),
		.A2(I4[19]),
		.B1(out_sel[5]),
		.B2(I5[19]),
		.Z(O2[19])
	);
	AO_CELL inst_3_19(
		.A1(out_sel[6]),
		.A2(I6[19]),
		.B1(out_sel[7]),
		.B2(I7[19]),
		.Z(O3[19])
	);
	AO_CELL inst_4_19(
		.A1(out_sel[8]),
		.A2(I8[19]),
		.B1(out_sel[9]),
		.B2(I9[19]),
		.Z(O4[19])
	);
	AO_CELL inst_5_19(
		.A1(out_sel[10]),
		.A2(I10[19]),
		.B1(out_sel[11]),
		.B2(I11[19]),
		.Z(O5[19])
	);
	AO_CELL inst_6_19(
		.A1(out_sel[12]),
		.A2(I12[19]),
		.B1(out_sel[13]),
		.B2(I13[19]),
		.Z(O6[19])
	);
	AO_CELL inst_7_19(
		.A1(out_sel[14]),
		.A2(I14[19]),
		.B1(out_sel[15]),
		.B2(I15[19]),
		.Z(O7[19])
	);
	AO_CELL inst_8_19(
		.A1(out_sel[16]),
		.A2(I16[19]),
		.B1(out_sel[17]),
		.B2(I17[19]),
		.Z(O8[19])
	);
	AO_CELL inst_0_20(
		.A1(out_sel[0]),
		.A2(I0[20]),
		.B1(out_sel[1]),
		.B2(I1[20]),
		.Z(O0[20])
	);
	AO_CELL inst_1_20(
		.A1(out_sel[2]),
		.A2(I2[20]),
		.B1(out_sel[3]),
		.B2(I3[20]),
		.Z(O1[20])
	);
	AO_CELL inst_2_20(
		.A1(out_sel[4]),
		.A2(I4[20]),
		.B1(out_sel[5]),
		.B2(I5[20]),
		.Z(O2[20])
	);
	AO_CELL inst_3_20(
		.A1(out_sel[6]),
		.A2(I6[20]),
		.B1(out_sel[7]),
		.B2(I7[20]),
		.Z(O3[20])
	);
	AO_CELL inst_4_20(
		.A1(out_sel[8]),
		.A2(I8[20]),
		.B1(out_sel[9]),
		.B2(I9[20]),
		.Z(O4[20])
	);
	AO_CELL inst_5_20(
		.A1(out_sel[10]),
		.A2(I10[20]),
		.B1(out_sel[11]),
		.B2(I11[20]),
		.Z(O5[20])
	);
	AO_CELL inst_6_20(
		.A1(out_sel[12]),
		.A2(I12[20]),
		.B1(out_sel[13]),
		.B2(I13[20]),
		.Z(O6[20])
	);
	AO_CELL inst_7_20(
		.A1(out_sel[14]),
		.A2(I14[20]),
		.B1(out_sel[15]),
		.B2(I15[20]),
		.Z(O7[20])
	);
	AO_CELL inst_8_20(
		.A1(out_sel[16]),
		.A2(I16[20]),
		.B1(out_sel[17]),
		.B2(I17[20]),
		.Z(O8[20])
	);
	AO_CELL inst_0_21(
		.A1(out_sel[0]),
		.A2(I0[21]),
		.B1(out_sel[1]),
		.B2(I1[21]),
		.Z(O0[21])
	);
	AO_CELL inst_1_21(
		.A1(out_sel[2]),
		.A2(I2[21]),
		.B1(out_sel[3]),
		.B2(I3[21]),
		.Z(O1[21])
	);
	AO_CELL inst_2_21(
		.A1(out_sel[4]),
		.A2(I4[21]),
		.B1(out_sel[5]),
		.B2(I5[21]),
		.Z(O2[21])
	);
	AO_CELL inst_3_21(
		.A1(out_sel[6]),
		.A2(I6[21]),
		.B1(out_sel[7]),
		.B2(I7[21]),
		.Z(O3[21])
	);
	AO_CELL inst_4_21(
		.A1(out_sel[8]),
		.A2(I8[21]),
		.B1(out_sel[9]),
		.B2(I9[21]),
		.Z(O4[21])
	);
	AO_CELL inst_5_21(
		.A1(out_sel[10]),
		.A2(I10[21]),
		.B1(out_sel[11]),
		.B2(I11[21]),
		.Z(O5[21])
	);
	AO_CELL inst_6_21(
		.A1(out_sel[12]),
		.A2(I12[21]),
		.B1(out_sel[13]),
		.B2(I13[21]),
		.Z(O6[21])
	);
	AO_CELL inst_7_21(
		.A1(out_sel[14]),
		.A2(I14[21]),
		.B1(out_sel[15]),
		.B2(I15[21]),
		.Z(O7[21])
	);
	AO_CELL inst_8_21(
		.A1(out_sel[16]),
		.A2(I16[21]),
		.B1(out_sel[17]),
		.B2(I17[21]),
		.Z(O8[21])
	);
	AO_CELL inst_0_22(
		.A1(out_sel[0]),
		.A2(I0[22]),
		.B1(out_sel[1]),
		.B2(I1[22]),
		.Z(O0[22])
	);
	AO_CELL inst_1_22(
		.A1(out_sel[2]),
		.A2(I2[22]),
		.B1(out_sel[3]),
		.B2(I3[22]),
		.Z(O1[22])
	);
	AO_CELL inst_2_22(
		.A1(out_sel[4]),
		.A2(I4[22]),
		.B1(out_sel[5]),
		.B2(I5[22]),
		.Z(O2[22])
	);
	AO_CELL inst_3_22(
		.A1(out_sel[6]),
		.A2(I6[22]),
		.B1(out_sel[7]),
		.B2(I7[22]),
		.Z(O3[22])
	);
	AO_CELL inst_4_22(
		.A1(out_sel[8]),
		.A2(I8[22]),
		.B1(out_sel[9]),
		.B2(I9[22]),
		.Z(O4[22])
	);
	AO_CELL inst_5_22(
		.A1(out_sel[10]),
		.A2(I10[22]),
		.B1(out_sel[11]),
		.B2(I11[22]),
		.Z(O5[22])
	);
	AO_CELL inst_6_22(
		.A1(out_sel[12]),
		.A2(I12[22]),
		.B1(out_sel[13]),
		.B2(I13[22]),
		.Z(O6[22])
	);
	AO_CELL inst_7_22(
		.A1(out_sel[14]),
		.A2(I14[22]),
		.B1(out_sel[15]),
		.B2(I15[22]),
		.Z(O7[22])
	);
	AO_CELL inst_8_22(
		.A1(out_sel[16]),
		.A2(I16[22]),
		.B1(out_sel[17]),
		.B2(I17[22]),
		.Z(O8[22])
	);
	AO_CELL inst_0_23(
		.A1(out_sel[0]),
		.A2(I0[23]),
		.B1(out_sel[1]),
		.B2(I1[23]),
		.Z(O0[23])
	);
	AO_CELL inst_1_23(
		.A1(out_sel[2]),
		.A2(I2[23]),
		.B1(out_sel[3]),
		.B2(I3[23]),
		.Z(O1[23])
	);
	AO_CELL inst_2_23(
		.A1(out_sel[4]),
		.A2(I4[23]),
		.B1(out_sel[5]),
		.B2(I5[23]),
		.Z(O2[23])
	);
	AO_CELL inst_3_23(
		.A1(out_sel[6]),
		.A2(I6[23]),
		.B1(out_sel[7]),
		.B2(I7[23]),
		.Z(O3[23])
	);
	AO_CELL inst_4_23(
		.A1(out_sel[8]),
		.A2(I8[23]),
		.B1(out_sel[9]),
		.B2(I9[23]),
		.Z(O4[23])
	);
	AO_CELL inst_5_23(
		.A1(out_sel[10]),
		.A2(I10[23]),
		.B1(out_sel[11]),
		.B2(I11[23]),
		.Z(O5[23])
	);
	AO_CELL inst_6_23(
		.A1(out_sel[12]),
		.A2(I12[23]),
		.B1(out_sel[13]),
		.B2(I13[23]),
		.Z(O6[23])
	);
	AO_CELL inst_7_23(
		.A1(out_sel[14]),
		.A2(I14[23]),
		.B1(out_sel[15]),
		.B2(I15[23]),
		.Z(O7[23])
	);
	AO_CELL inst_8_23(
		.A1(out_sel[16]),
		.A2(I16[23]),
		.B1(out_sel[17]),
		.B2(I17[23]),
		.Z(O8[23])
	);
	AO_CELL inst_0_24(
		.A1(out_sel[0]),
		.A2(I0[24]),
		.B1(out_sel[1]),
		.B2(I1[24]),
		.Z(O0[24])
	);
	AO_CELL inst_1_24(
		.A1(out_sel[2]),
		.A2(I2[24]),
		.B1(out_sel[3]),
		.B2(I3[24]),
		.Z(O1[24])
	);
	AO_CELL inst_2_24(
		.A1(out_sel[4]),
		.A2(I4[24]),
		.B1(out_sel[5]),
		.B2(I5[24]),
		.Z(O2[24])
	);
	AO_CELL inst_3_24(
		.A1(out_sel[6]),
		.A2(I6[24]),
		.B1(out_sel[7]),
		.B2(I7[24]),
		.Z(O3[24])
	);
	AO_CELL inst_4_24(
		.A1(out_sel[8]),
		.A2(I8[24]),
		.B1(out_sel[9]),
		.B2(I9[24]),
		.Z(O4[24])
	);
	AO_CELL inst_5_24(
		.A1(out_sel[10]),
		.A2(I10[24]),
		.B1(out_sel[11]),
		.B2(I11[24]),
		.Z(O5[24])
	);
	AO_CELL inst_6_24(
		.A1(out_sel[12]),
		.A2(I12[24]),
		.B1(out_sel[13]),
		.B2(I13[24]),
		.Z(O6[24])
	);
	AO_CELL inst_7_24(
		.A1(out_sel[14]),
		.A2(I14[24]),
		.B1(out_sel[15]),
		.B2(I15[24]),
		.Z(O7[24])
	);
	AO_CELL inst_8_24(
		.A1(out_sel[16]),
		.A2(I16[24]),
		.B1(out_sel[17]),
		.B2(I17[24]),
		.Z(O8[24])
	);
	AO_CELL inst_0_25(
		.A1(out_sel[0]),
		.A2(I0[25]),
		.B1(out_sel[1]),
		.B2(I1[25]),
		.Z(O0[25])
	);
	AO_CELL inst_1_25(
		.A1(out_sel[2]),
		.A2(I2[25]),
		.B1(out_sel[3]),
		.B2(I3[25]),
		.Z(O1[25])
	);
	AO_CELL inst_2_25(
		.A1(out_sel[4]),
		.A2(I4[25]),
		.B1(out_sel[5]),
		.B2(I5[25]),
		.Z(O2[25])
	);
	AO_CELL inst_3_25(
		.A1(out_sel[6]),
		.A2(I6[25]),
		.B1(out_sel[7]),
		.B2(I7[25]),
		.Z(O3[25])
	);
	AO_CELL inst_4_25(
		.A1(out_sel[8]),
		.A2(I8[25]),
		.B1(out_sel[9]),
		.B2(I9[25]),
		.Z(O4[25])
	);
	AO_CELL inst_5_25(
		.A1(out_sel[10]),
		.A2(I10[25]),
		.B1(out_sel[11]),
		.B2(I11[25]),
		.Z(O5[25])
	);
	AO_CELL inst_6_25(
		.A1(out_sel[12]),
		.A2(I12[25]),
		.B1(out_sel[13]),
		.B2(I13[25]),
		.Z(O6[25])
	);
	AO_CELL inst_7_25(
		.A1(out_sel[14]),
		.A2(I14[25]),
		.B1(out_sel[15]),
		.B2(I15[25]),
		.Z(O7[25])
	);
	AO_CELL inst_8_25(
		.A1(out_sel[16]),
		.A2(I16[25]),
		.B1(out_sel[17]),
		.B2(I17[25]),
		.Z(O8[25])
	);
	AO_CELL inst_0_26(
		.A1(out_sel[0]),
		.A2(I0[26]),
		.B1(out_sel[1]),
		.B2(I1[26]),
		.Z(O0[26])
	);
	AO_CELL inst_1_26(
		.A1(out_sel[2]),
		.A2(I2[26]),
		.B1(out_sel[3]),
		.B2(I3[26]),
		.Z(O1[26])
	);
	AO_CELL inst_2_26(
		.A1(out_sel[4]),
		.A2(I4[26]),
		.B1(out_sel[5]),
		.B2(I5[26]),
		.Z(O2[26])
	);
	AO_CELL inst_3_26(
		.A1(out_sel[6]),
		.A2(I6[26]),
		.B1(out_sel[7]),
		.B2(I7[26]),
		.Z(O3[26])
	);
	AO_CELL inst_4_26(
		.A1(out_sel[8]),
		.A2(I8[26]),
		.B1(out_sel[9]),
		.B2(I9[26]),
		.Z(O4[26])
	);
	AO_CELL inst_5_26(
		.A1(out_sel[10]),
		.A2(I10[26]),
		.B1(out_sel[11]),
		.B2(I11[26]),
		.Z(O5[26])
	);
	AO_CELL inst_6_26(
		.A1(out_sel[12]),
		.A2(I12[26]),
		.B1(out_sel[13]),
		.B2(I13[26]),
		.Z(O6[26])
	);
	AO_CELL inst_7_26(
		.A1(out_sel[14]),
		.A2(I14[26]),
		.B1(out_sel[15]),
		.B2(I15[26]),
		.Z(O7[26])
	);
	AO_CELL inst_8_26(
		.A1(out_sel[16]),
		.A2(I16[26]),
		.B1(out_sel[17]),
		.B2(I17[26]),
		.Z(O8[26])
	);
	AO_CELL inst_0_27(
		.A1(out_sel[0]),
		.A2(I0[27]),
		.B1(out_sel[1]),
		.B2(I1[27]),
		.Z(O0[27])
	);
	AO_CELL inst_1_27(
		.A1(out_sel[2]),
		.A2(I2[27]),
		.B1(out_sel[3]),
		.B2(I3[27]),
		.Z(O1[27])
	);
	AO_CELL inst_2_27(
		.A1(out_sel[4]),
		.A2(I4[27]),
		.B1(out_sel[5]),
		.B2(I5[27]),
		.Z(O2[27])
	);
	AO_CELL inst_3_27(
		.A1(out_sel[6]),
		.A2(I6[27]),
		.B1(out_sel[7]),
		.B2(I7[27]),
		.Z(O3[27])
	);
	AO_CELL inst_4_27(
		.A1(out_sel[8]),
		.A2(I8[27]),
		.B1(out_sel[9]),
		.B2(I9[27]),
		.Z(O4[27])
	);
	AO_CELL inst_5_27(
		.A1(out_sel[10]),
		.A2(I10[27]),
		.B1(out_sel[11]),
		.B2(I11[27]),
		.Z(O5[27])
	);
	AO_CELL inst_6_27(
		.A1(out_sel[12]),
		.A2(I12[27]),
		.B1(out_sel[13]),
		.B2(I13[27]),
		.Z(O6[27])
	);
	AO_CELL inst_7_27(
		.A1(out_sel[14]),
		.A2(I14[27]),
		.B1(out_sel[15]),
		.B2(I15[27]),
		.Z(O7[27])
	);
	AO_CELL inst_8_27(
		.A1(out_sel[16]),
		.A2(I16[27]),
		.B1(out_sel[17]),
		.B2(I17[27]),
		.Z(O8[27])
	);
	AO_CELL inst_0_28(
		.A1(out_sel[0]),
		.A2(I0[28]),
		.B1(out_sel[1]),
		.B2(I1[28]),
		.Z(O0[28])
	);
	AO_CELL inst_1_28(
		.A1(out_sel[2]),
		.A2(I2[28]),
		.B1(out_sel[3]),
		.B2(I3[28]),
		.Z(O1[28])
	);
	AO_CELL inst_2_28(
		.A1(out_sel[4]),
		.A2(I4[28]),
		.B1(out_sel[5]),
		.B2(I5[28]),
		.Z(O2[28])
	);
	AO_CELL inst_3_28(
		.A1(out_sel[6]),
		.A2(I6[28]),
		.B1(out_sel[7]),
		.B2(I7[28]),
		.Z(O3[28])
	);
	AO_CELL inst_4_28(
		.A1(out_sel[8]),
		.A2(I8[28]),
		.B1(out_sel[9]),
		.B2(I9[28]),
		.Z(O4[28])
	);
	AO_CELL inst_5_28(
		.A1(out_sel[10]),
		.A2(I10[28]),
		.B1(out_sel[11]),
		.B2(I11[28]),
		.Z(O5[28])
	);
	AO_CELL inst_6_28(
		.A1(out_sel[12]),
		.A2(I12[28]),
		.B1(out_sel[13]),
		.B2(I13[28]),
		.Z(O6[28])
	);
	AO_CELL inst_7_28(
		.A1(out_sel[14]),
		.A2(I14[28]),
		.B1(out_sel[15]),
		.B2(I15[28]),
		.Z(O7[28])
	);
	AO_CELL inst_8_28(
		.A1(out_sel[16]),
		.A2(I16[28]),
		.B1(out_sel[17]),
		.B2(I17[28]),
		.Z(O8[28])
	);
	AO_CELL inst_0_29(
		.A1(out_sel[0]),
		.A2(I0[29]),
		.B1(out_sel[1]),
		.B2(I1[29]),
		.Z(O0[29])
	);
	AO_CELL inst_1_29(
		.A1(out_sel[2]),
		.A2(I2[29]),
		.B1(out_sel[3]),
		.B2(I3[29]),
		.Z(O1[29])
	);
	AO_CELL inst_2_29(
		.A1(out_sel[4]),
		.A2(I4[29]),
		.B1(out_sel[5]),
		.B2(I5[29]),
		.Z(O2[29])
	);
	AO_CELL inst_3_29(
		.A1(out_sel[6]),
		.A2(I6[29]),
		.B1(out_sel[7]),
		.B2(I7[29]),
		.Z(O3[29])
	);
	AO_CELL inst_4_29(
		.A1(out_sel[8]),
		.A2(I8[29]),
		.B1(out_sel[9]),
		.B2(I9[29]),
		.Z(O4[29])
	);
	AO_CELL inst_5_29(
		.A1(out_sel[10]),
		.A2(I10[29]),
		.B1(out_sel[11]),
		.B2(I11[29]),
		.Z(O5[29])
	);
	AO_CELL inst_6_29(
		.A1(out_sel[12]),
		.A2(I12[29]),
		.B1(out_sel[13]),
		.B2(I13[29]),
		.Z(O6[29])
	);
	AO_CELL inst_7_29(
		.A1(out_sel[14]),
		.A2(I14[29]),
		.B1(out_sel[15]),
		.B2(I15[29]),
		.Z(O7[29])
	);
	AO_CELL inst_8_29(
		.A1(out_sel[16]),
		.A2(I16[29]),
		.B1(out_sel[17]),
		.B2(I17[29]),
		.Z(O8[29])
	);
	AO_CELL inst_0_30(
		.A1(out_sel[0]),
		.A2(I0[30]),
		.B1(out_sel[1]),
		.B2(I1[30]),
		.Z(O0[30])
	);
	AO_CELL inst_1_30(
		.A1(out_sel[2]),
		.A2(I2[30]),
		.B1(out_sel[3]),
		.B2(I3[30]),
		.Z(O1[30])
	);
	AO_CELL inst_2_30(
		.A1(out_sel[4]),
		.A2(I4[30]),
		.B1(out_sel[5]),
		.B2(I5[30]),
		.Z(O2[30])
	);
	AO_CELL inst_3_30(
		.A1(out_sel[6]),
		.A2(I6[30]),
		.B1(out_sel[7]),
		.B2(I7[30]),
		.Z(O3[30])
	);
	AO_CELL inst_4_30(
		.A1(out_sel[8]),
		.A2(I8[30]),
		.B1(out_sel[9]),
		.B2(I9[30]),
		.Z(O4[30])
	);
	AO_CELL inst_5_30(
		.A1(out_sel[10]),
		.A2(I10[30]),
		.B1(out_sel[11]),
		.B2(I11[30]),
		.Z(O5[30])
	);
	AO_CELL inst_6_30(
		.A1(out_sel[12]),
		.A2(I12[30]),
		.B1(out_sel[13]),
		.B2(I13[30]),
		.Z(O6[30])
	);
	AO_CELL inst_7_30(
		.A1(out_sel[14]),
		.A2(I14[30]),
		.B1(out_sel[15]),
		.B2(I15[30]),
		.Z(O7[30])
	);
	AO_CELL inst_8_30(
		.A1(out_sel[16]),
		.A2(I16[30]),
		.B1(out_sel[17]),
		.B2(I17[30]),
		.Z(O8[30])
	);
	AO_CELL inst_0_31(
		.A1(out_sel[0]),
		.A2(I0[31]),
		.B1(out_sel[1]),
		.B2(I1[31]),
		.Z(O0[31])
	);
	AO_CELL inst_1_31(
		.A1(out_sel[2]),
		.A2(I2[31]),
		.B1(out_sel[3]),
		.B2(I3[31]),
		.Z(O1[31])
	);
	AO_CELL inst_2_31(
		.A1(out_sel[4]),
		.A2(I4[31]),
		.B1(out_sel[5]),
		.B2(I5[31]),
		.Z(O2[31])
	);
	AO_CELL inst_3_31(
		.A1(out_sel[6]),
		.A2(I6[31]),
		.B1(out_sel[7]),
		.B2(I7[31]),
		.Z(O3[31])
	);
	AO_CELL inst_4_31(
		.A1(out_sel[8]),
		.A2(I8[31]),
		.B1(out_sel[9]),
		.B2(I9[31]),
		.Z(O4[31])
	);
	AO_CELL inst_5_31(
		.A1(out_sel[10]),
		.A2(I10[31]),
		.B1(out_sel[11]),
		.B2(I11[31]),
		.Z(O5[31])
	);
	AO_CELL inst_6_31(
		.A1(out_sel[12]),
		.A2(I12[31]),
		.B1(out_sel[13]),
		.B2(I13[31]),
		.Z(O6[31])
	);
	AO_CELL inst_7_31(
		.A1(out_sel[14]),
		.A2(I14[31]),
		.B1(out_sel[15]),
		.B2(I15[31]),
		.Z(O7[31])
	);
	AO_CELL inst_8_31(
		.A1(out_sel[16]),
		.A2(I16[31]),
		.B1(out_sel[17]),
		.B2(I17[31]),
		.Z(O8[31])
	);
endmodule
module mux_aoi_16_32 (
	I,
	S,
	out_sel,
	O
);
	input wire [511:0] I;
	input wire [3:0] S;
	output wire [15:0] out_sel;
	output wire [31:0] O;
	wire [31:0] O_int0;
	wire [31:0] O_int1;
	wire [31:0] O_int2;
	wire [31:0] O_int3;
	wire [31:0] O_int4;
	wire [31:0] O_int5;
	wire [31:0] O_int6;
	wire [31:0] O_int7;
	precoder_32_16 u_precoder(
		.S(S),
		.out_sel(out_sel)
	);
	mux_logic_32_16 u_mux_logic(
		.I0(I[0+:32]),
		.I1(I[32+:32]),
		.I2(I[64+:32]),
		.I3(I[96+:32]),
		.I4(I[128+:32]),
		.I5(I[160+:32]),
		.I6(I[192+:32]),
		.I7(I[224+:32]),
		.I8(I[256+:32]),
		.I9(I[288+:32]),
		.I10(I[320+:32]),
		.I11(I[352+:32]),
		.I12(I[384+:32]),
		.I13(I[416+:32]),
		.I14(I[448+:32]),
		.I15(I[480+:32]),
		.out_sel(out_sel),
		.O0(O_int0),
		.O1(O_int1),
		.O2(O_int2),
		.O3(O_int3),
		.O4(O_int4),
		.O5(O_int5),
		.O6(O_int6),
		.O7(O_int7)
	);
	assign O = ((((((O_int0 | O_int1) | O_int2) | O_int3) | O_int4) | O_int5) | O_int6) | O_int7;
endmodule
module precoder_32_16 (
	S,
	out_sel
);
	input wire [3:0] S;
	output reg [15:0] out_sel;
	always @(*) begin : mux_sel
		case (S)
			4'd0: out_sel = 16'b0000000000000001;
			4'd1: out_sel = 16'b0000000000000010;
			4'd2: out_sel = 16'b0000000000000100;
			4'd3: out_sel = 16'b0000000000001000;
			4'd4: out_sel = 16'b0000000000010000;
			4'd5: out_sel = 16'b0000000000100000;
			4'd6: out_sel = 16'b0000000001000000;
			4'd7: out_sel = 16'b0000000010000000;
			4'd8: out_sel = 16'b0000000100000000;
			4'd9: out_sel = 16'b0000001000000000;
			4'd10: out_sel = 16'b0000010000000000;
			4'd11: out_sel = 16'b0000100000000000;
			4'd12: out_sel = 16'b0001000000000000;
			4'd13: out_sel = 16'b0010000000000000;
			4'd14: out_sel = 16'b0100000000000000;
			4'd15: out_sel = 16'b1000000000000000;
			default: out_sel = 16'b0000000000000000;
		endcase
	end
endmodule
module mux_logic_32_16 (
	out_sel,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	I9,
	I10,
	I11,
	I12,
	I13,
	I14,
	I15,
	O0,
	O1,
	O2,
	O3,
	O4,
	O5,
	O6,
	O7
);
	input wire [15:0] out_sel;
	input wire [31:0] I0;
	input wire [31:0] I1;
	input wire [31:0] I2;
	input wire [31:0] I3;
	input wire [31:0] I4;
	input wire [31:0] I5;
	input wire [31:0] I6;
	input wire [31:0] I7;
	input wire [31:0] I8;
	input wire [31:0] I9;
	input wire [31:0] I10;
	input wire [31:0] I11;
	input wire [31:0] I12;
	input wire [31:0] I13;
	input wire [31:0] I14;
	input wire [31:0] I15;
	output wire [31:0] O0;
	output wire [31:0] O1;
	output wire [31:0] O2;
	output wire [31:0] O3;
	output wire [31:0] O4;
	output wire [31:0] O5;
	output wire [31:0] O6;
	output wire [31:0] O7;
	AO_CELL inst_0_0(
		.A1(out_sel[0]),
		.A2(I0[0]),
		.B1(out_sel[1]),
		.B2(I1[0]),
		.Z(O0[0])
	);
	AO_CELL inst_1_0(
		.A1(out_sel[2]),
		.A2(I2[0]),
		.B1(out_sel[3]),
		.B2(I3[0]),
		.Z(O1[0])
	);
	AO_CELL inst_2_0(
		.A1(out_sel[4]),
		.A2(I4[0]),
		.B1(out_sel[5]),
		.B2(I5[0]),
		.Z(O2[0])
	);
	AO_CELL inst_3_0(
		.A1(out_sel[6]),
		.A2(I6[0]),
		.B1(out_sel[7]),
		.B2(I7[0]),
		.Z(O3[0])
	);
	AO_CELL inst_4_0(
		.A1(out_sel[8]),
		.A2(I8[0]),
		.B1(out_sel[9]),
		.B2(I9[0]),
		.Z(O4[0])
	);
	AO_CELL inst_5_0(
		.A1(out_sel[10]),
		.A2(I10[0]),
		.B1(out_sel[11]),
		.B2(I11[0]),
		.Z(O5[0])
	);
	AO_CELL inst_6_0(
		.A1(out_sel[12]),
		.A2(I12[0]),
		.B1(out_sel[13]),
		.B2(I13[0]),
		.Z(O6[0])
	);
	AO_CELL inst_7_0(
		.A1(out_sel[14]),
		.A2(I14[0]),
		.B1(out_sel[15]),
		.B2(I15[0]),
		.Z(O7[0])
	);
	AO_CELL inst_0_1(
		.A1(out_sel[0]),
		.A2(I0[1]),
		.B1(out_sel[1]),
		.B2(I1[1]),
		.Z(O0[1])
	);
	AO_CELL inst_1_1(
		.A1(out_sel[2]),
		.A2(I2[1]),
		.B1(out_sel[3]),
		.B2(I3[1]),
		.Z(O1[1])
	);
	AO_CELL inst_2_1(
		.A1(out_sel[4]),
		.A2(I4[1]),
		.B1(out_sel[5]),
		.B2(I5[1]),
		.Z(O2[1])
	);
	AO_CELL inst_3_1(
		.A1(out_sel[6]),
		.A2(I6[1]),
		.B1(out_sel[7]),
		.B2(I7[1]),
		.Z(O3[1])
	);
	AO_CELL inst_4_1(
		.A1(out_sel[8]),
		.A2(I8[1]),
		.B1(out_sel[9]),
		.B2(I9[1]),
		.Z(O4[1])
	);
	AO_CELL inst_5_1(
		.A1(out_sel[10]),
		.A2(I10[1]),
		.B1(out_sel[11]),
		.B2(I11[1]),
		.Z(O5[1])
	);
	AO_CELL inst_6_1(
		.A1(out_sel[12]),
		.A2(I12[1]),
		.B1(out_sel[13]),
		.B2(I13[1]),
		.Z(O6[1])
	);
	AO_CELL inst_7_1(
		.A1(out_sel[14]),
		.A2(I14[1]),
		.B1(out_sel[15]),
		.B2(I15[1]),
		.Z(O7[1])
	);
	AO_CELL inst_0_2(
		.A1(out_sel[0]),
		.A2(I0[2]),
		.B1(out_sel[1]),
		.B2(I1[2]),
		.Z(O0[2])
	);
	AO_CELL inst_1_2(
		.A1(out_sel[2]),
		.A2(I2[2]),
		.B1(out_sel[3]),
		.B2(I3[2]),
		.Z(O1[2])
	);
	AO_CELL inst_2_2(
		.A1(out_sel[4]),
		.A2(I4[2]),
		.B1(out_sel[5]),
		.B2(I5[2]),
		.Z(O2[2])
	);
	AO_CELL inst_3_2(
		.A1(out_sel[6]),
		.A2(I6[2]),
		.B1(out_sel[7]),
		.B2(I7[2]),
		.Z(O3[2])
	);
	AO_CELL inst_4_2(
		.A1(out_sel[8]),
		.A2(I8[2]),
		.B1(out_sel[9]),
		.B2(I9[2]),
		.Z(O4[2])
	);
	AO_CELL inst_5_2(
		.A1(out_sel[10]),
		.A2(I10[2]),
		.B1(out_sel[11]),
		.B2(I11[2]),
		.Z(O5[2])
	);
	AO_CELL inst_6_2(
		.A1(out_sel[12]),
		.A2(I12[2]),
		.B1(out_sel[13]),
		.B2(I13[2]),
		.Z(O6[2])
	);
	AO_CELL inst_7_2(
		.A1(out_sel[14]),
		.A2(I14[2]),
		.B1(out_sel[15]),
		.B2(I15[2]),
		.Z(O7[2])
	);
	AO_CELL inst_0_3(
		.A1(out_sel[0]),
		.A2(I0[3]),
		.B1(out_sel[1]),
		.B2(I1[3]),
		.Z(O0[3])
	);
	AO_CELL inst_1_3(
		.A1(out_sel[2]),
		.A2(I2[3]),
		.B1(out_sel[3]),
		.B2(I3[3]),
		.Z(O1[3])
	);
	AO_CELL inst_2_3(
		.A1(out_sel[4]),
		.A2(I4[3]),
		.B1(out_sel[5]),
		.B2(I5[3]),
		.Z(O2[3])
	);
	AO_CELL inst_3_3(
		.A1(out_sel[6]),
		.A2(I6[3]),
		.B1(out_sel[7]),
		.B2(I7[3]),
		.Z(O3[3])
	);
	AO_CELL inst_4_3(
		.A1(out_sel[8]),
		.A2(I8[3]),
		.B1(out_sel[9]),
		.B2(I9[3]),
		.Z(O4[3])
	);
	AO_CELL inst_5_3(
		.A1(out_sel[10]),
		.A2(I10[3]),
		.B1(out_sel[11]),
		.B2(I11[3]),
		.Z(O5[3])
	);
	AO_CELL inst_6_3(
		.A1(out_sel[12]),
		.A2(I12[3]),
		.B1(out_sel[13]),
		.B2(I13[3]),
		.Z(O6[3])
	);
	AO_CELL inst_7_3(
		.A1(out_sel[14]),
		.A2(I14[3]),
		.B1(out_sel[15]),
		.B2(I15[3]),
		.Z(O7[3])
	);
	AO_CELL inst_0_4(
		.A1(out_sel[0]),
		.A2(I0[4]),
		.B1(out_sel[1]),
		.B2(I1[4]),
		.Z(O0[4])
	);
	AO_CELL inst_1_4(
		.A1(out_sel[2]),
		.A2(I2[4]),
		.B1(out_sel[3]),
		.B2(I3[4]),
		.Z(O1[4])
	);
	AO_CELL inst_2_4(
		.A1(out_sel[4]),
		.A2(I4[4]),
		.B1(out_sel[5]),
		.B2(I5[4]),
		.Z(O2[4])
	);
	AO_CELL inst_3_4(
		.A1(out_sel[6]),
		.A2(I6[4]),
		.B1(out_sel[7]),
		.B2(I7[4]),
		.Z(O3[4])
	);
	AO_CELL inst_4_4(
		.A1(out_sel[8]),
		.A2(I8[4]),
		.B1(out_sel[9]),
		.B2(I9[4]),
		.Z(O4[4])
	);
	AO_CELL inst_5_4(
		.A1(out_sel[10]),
		.A2(I10[4]),
		.B1(out_sel[11]),
		.B2(I11[4]),
		.Z(O5[4])
	);
	AO_CELL inst_6_4(
		.A1(out_sel[12]),
		.A2(I12[4]),
		.B1(out_sel[13]),
		.B2(I13[4]),
		.Z(O6[4])
	);
	AO_CELL inst_7_4(
		.A1(out_sel[14]),
		.A2(I14[4]),
		.B1(out_sel[15]),
		.B2(I15[4]),
		.Z(O7[4])
	);
	AO_CELL inst_0_5(
		.A1(out_sel[0]),
		.A2(I0[5]),
		.B1(out_sel[1]),
		.B2(I1[5]),
		.Z(O0[5])
	);
	AO_CELL inst_1_5(
		.A1(out_sel[2]),
		.A2(I2[5]),
		.B1(out_sel[3]),
		.B2(I3[5]),
		.Z(O1[5])
	);
	AO_CELL inst_2_5(
		.A1(out_sel[4]),
		.A2(I4[5]),
		.B1(out_sel[5]),
		.B2(I5[5]),
		.Z(O2[5])
	);
	AO_CELL inst_3_5(
		.A1(out_sel[6]),
		.A2(I6[5]),
		.B1(out_sel[7]),
		.B2(I7[5]),
		.Z(O3[5])
	);
	AO_CELL inst_4_5(
		.A1(out_sel[8]),
		.A2(I8[5]),
		.B1(out_sel[9]),
		.B2(I9[5]),
		.Z(O4[5])
	);
	AO_CELL inst_5_5(
		.A1(out_sel[10]),
		.A2(I10[5]),
		.B1(out_sel[11]),
		.B2(I11[5]),
		.Z(O5[5])
	);
	AO_CELL inst_6_5(
		.A1(out_sel[12]),
		.A2(I12[5]),
		.B1(out_sel[13]),
		.B2(I13[5]),
		.Z(O6[5])
	);
	AO_CELL inst_7_5(
		.A1(out_sel[14]),
		.A2(I14[5]),
		.B1(out_sel[15]),
		.B2(I15[5]),
		.Z(O7[5])
	);
	AO_CELL inst_0_6(
		.A1(out_sel[0]),
		.A2(I0[6]),
		.B1(out_sel[1]),
		.B2(I1[6]),
		.Z(O0[6])
	);
	AO_CELL inst_1_6(
		.A1(out_sel[2]),
		.A2(I2[6]),
		.B1(out_sel[3]),
		.B2(I3[6]),
		.Z(O1[6])
	);
	AO_CELL inst_2_6(
		.A1(out_sel[4]),
		.A2(I4[6]),
		.B1(out_sel[5]),
		.B2(I5[6]),
		.Z(O2[6])
	);
	AO_CELL inst_3_6(
		.A1(out_sel[6]),
		.A2(I6[6]),
		.B1(out_sel[7]),
		.B2(I7[6]),
		.Z(O3[6])
	);
	AO_CELL inst_4_6(
		.A1(out_sel[8]),
		.A2(I8[6]),
		.B1(out_sel[9]),
		.B2(I9[6]),
		.Z(O4[6])
	);
	AO_CELL inst_5_6(
		.A1(out_sel[10]),
		.A2(I10[6]),
		.B1(out_sel[11]),
		.B2(I11[6]),
		.Z(O5[6])
	);
	AO_CELL inst_6_6(
		.A1(out_sel[12]),
		.A2(I12[6]),
		.B1(out_sel[13]),
		.B2(I13[6]),
		.Z(O6[6])
	);
	AO_CELL inst_7_6(
		.A1(out_sel[14]),
		.A2(I14[6]),
		.B1(out_sel[15]),
		.B2(I15[6]),
		.Z(O7[6])
	);
	AO_CELL inst_0_7(
		.A1(out_sel[0]),
		.A2(I0[7]),
		.B1(out_sel[1]),
		.B2(I1[7]),
		.Z(O0[7])
	);
	AO_CELL inst_1_7(
		.A1(out_sel[2]),
		.A2(I2[7]),
		.B1(out_sel[3]),
		.B2(I3[7]),
		.Z(O1[7])
	);
	AO_CELL inst_2_7(
		.A1(out_sel[4]),
		.A2(I4[7]),
		.B1(out_sel[5]),
		.B2(I5[7]),
		.Z(O2[7])
	);
	AO_CELL inst_3_7(
		.A1(out_sel[6]),
		.A2(I6[7]),
		.B1(out_sel[7]),
		.B2(I7[7]),
		.Z(O3[7])
	);
	AO_CELL inst_4_7(
		.A1(out_sel[8]),
		.A2(I8[7]),
		.B1(out_sel[9]),
		.B2(I9[7]),
		.Z(O4[7])
	);
	AO_CELL inst_5_7(
		.A1(out_sel[10]),
		.A2(I10[7]),
		.B1(out_sel[11]),
		.B2(I11[7]),
		.Z(O5[7])
	);
	AO_CELL inst_6_7(
		.A1(out_sel[12]),
		.A2(I12[7]),
		.B1(out_sel[13]),
		.B2(I13[7]),
		.Z(O6[7])
	);
	AO_CELL inst_7_7(
		.A1(out_sel[14]),
		.A2(I14[7]),
		.B1(out_sel[15]),
		.B2(I15[7]),
		.Z(O7[7])
	);
	AO_CELL inst_0_8(
		.A1(out_sel[0]),
		.A2(I0[8]),
		.B1(out_sel[1]),
		.B2(I1[8]),
		.Z(O0[8])
	);
	AO_CELL inst_1_8(
		.A1(out_sel[2]),
		.A2(I2[8]),
		.B1(out_sel[3]),
		.B2(I3[8]),
		.Z(O1[8])
	);
	AO_CELL inst_2_8(
		.A1(out_sel[4]),
		.A2(I4[8]),
		.B1(out_sel[5]),
		.B2(I5[8]),
		.Z(O2[8])
	);
	AO_CELL inst_3_8(
		.A1(out_sel[6]),
		.A2(I6[8]),
		.B1(out_sel[7]),
		.B2(I7[8]),
		.Z(O3[8])
	);
	AO_CELL inst_4_8(
		.A1(out_sel[8]),
		.A2(I8[8]),
		.B1(out_sel[9]),
		.B2(I9[8]),
		.Z(O4[8])
	);
	AO_CELL inst_5_8(
		.A1(out_sel[10]),
		.A2(I10[8]),
		.B1(out_sel[11]),
		.B2(I11[8]),
		.Z(O5[8])
	);
	AO_CELL inst_6_8(
		.A1(out_sel[12]),
		.A2(I12[8]),
		.B1(out_sel[13]),
		.B2(I13[8]),
		.Z(O6[8])
	);
	AO_CELL inst_7_8(
		.A1(out_sel[14]),
		.A2(I14[8]),
		.B1(out_sel[15]),
		.B2(I15[8]),
		.Z(O7[8])
	);
	AO_CELL inst_0_9(
		.A1(out_sel[0]),
		.A2(I0[9]),
		.B1(out_sel[1]),
		.B2(I1[9]),
		.Z(O0[9])
	);
	AO_CELL inst_1_9(
		.A1(out_sel[2]),
		.A2(I2[9]),
		.B1(out_sel[3]),
		.B2(I3[9]),
		.Z(O1[9])
	);
	AO_CELL inst_2_9(
		.A1(out_sel[4]),
		.A2(I4[9]),
		.B1(out_sel[5]),
		.B2(I5[9]),
		.Z(O2[9])
	);
	AO_CELL inst_3_9(
		.A1(out_sel[6]),
		.A2(I6[9]),
		.B1(out_sel[7]),
		.B2(I7[9]),
		.Z(O3[9])
	);
	AO_CELL inst_4_9(
		.A1(out_sel[8]),
		.A2(I8[9]),
		.B1(out_sel[9]),
		.B2(I9[9]),
		.Z(O4[9])
	);
	AO_CELL inst_5_9(
		.A1(out_sel[10]),
		.A2(I10[9]),
		.B1(out_sel[11]),
		.B2(I11[9]),
		.Z(O5[9])
	);
	AO_CELL inst_6_9(
		.A1(out_sel[12]),
		.A2(I12[9]),
		.B1(out_sel[13]),
		.B2(I13[9]),
		.Z(O6[9])
	);
	AO_CELL inst_7_9(
		.A1(out_sel[14]),
		.A2(I14[9]),
		.B1(out_sel[15]),
		.B2(I15[9]),
		.Z(O7[9])
	);
	AO_CELL inst_0_10(
		.A1(out_sel[0]),
		.A2(I0[10]),
		.B1(out_sel[1]),
		.B2(I1[10]),
		.Z(O0[10])
	);
	AO_CELL inst_1_10(
		.A1(out_sel[2]),
		.A2(I2[10]),
		.B1(out_sel[3]),
		.B2(I3[10]),
		.Z(O1[10])
	);
	AO_CELL inst_2_10(
		.A1(out_sel[4]),
		.A2(I4[10]),
		.B1(out_sel[5]),
		.B2(I5[10]),
		.Z(O2[10])
	);
	AO_CELL inst_3_10(
		.A1(out_sel[6]),
		.A2(I6[10]),
		.B1(out_sel[7]),
		.B2(I7[10]),
		.Z(O3[10])
	);
	AO_CELL inst_4_10(
		.A1(out_sel[8]),
		.A2(I8[10]),
		.B1(out_sel[9]),
		.B2(I9[10]),
		.Z(O4[10])
	);
	AO_CELL inst_5_10(
		.A1(out_sel[10]),
		.A2(I10[10]),
		.B1(out_sel[11]),
		.B2(I11[10]),
		.Z(O5[10])
	);
	AO_CELL inst_6_10(
		.A1(out_sel[12]),
		.A2(I12[10]),
		.B1(out_sel[13]),
		.B2(I13[10]),
		.Z(O6[10])
	);
	AO_CELL inst_7_10(
		.A1(out_sel[14]),
		.A2(I14[10]),
		.B1(out_sel[15]),
		.B2(I15[10]),
		.Z(O7[10])
	);
	AO_CELL inst_0_11(
		.A1(out_sel[0]),
		.A2(I0[11]),
		.B1(out_sel[1]),
		.B2(I1[11]),
		.Z(O0[11])
	);
	AO_CELL inst_1_11(
		.A1(out_sel[2]),
		.A2(I2[11]),
		.B1(out_sel[3]),
		.B2(I3[11]),
		.Z(O1[11])
	);
	AO_CELL inst_2_11(
		.A1(out_sel[4]),
		.A2(I4[11]),
		.B1(out_sel[5]),
		.B2(I5[11]),
		.Z(O2[11])
	);
	AO_CELL inst_3_11(
		.A1(out_sel[6]),
		.A2(I6[11]),
		.B1(out_sel[7]),
		.B2(I7[11]),
		.Z(O3[11])
	);
	AO_CELL inst_4_11(
		.A1(out_sel[8]),
		.A2(I8[11]),
		.B1(out_sel[9]),
		.B2(I9[11]),
		.Z(O4[11])
	);
	AO_CELL inst_5_11(
		.A1(out_sel[10]),
		.A2(I10[11]),
		.B1(out_sel[11]),
		.B2(I11[11]),
		.Z(O5[11])
	);
	AO_CELL inst_6_11(
		.A1(out_sel[12]),
		.A2(I12[11]),
		.B1(out_sel[13]),
		.B2(I13[11]),
		.Z(O6[11])
	);
	AO_CELL inst_7_11(
		.A1(out_sel[14]),
		.A2(I14[11]),
		.B1(out_sel[15]),
		.B2(I15[11]),
		.Z(O7[11])
	);
	AO_CELL inst_0_12(
		.A1(out_sel[0]),
		.A2(I0[12]),
		.B1(out_sel[1]),
		.B2(I1[12]),
		.Z(O0[12])
	);
	AO_CELL inst_1_12(
		.A1(out_sel[2]),
		.A2(I2[12]),
		.B1(out_sel[3]),
		.B2(I3[12]),
		.Z(O1[12])
	);
	AO_CELL inst_2_12(
		.A1(out_sel[4]),
		.A2(I4[12]),
		.B1(out_sel[5]),
		.B2(I5[12]),
		.Z(O2[12])
	);
	AO_CELL inst_3_12(
		.A1(out_sel[6]),
		.A2(I6[12]),
		.B1(out_sel[7]),
		.B2(I7[12]),
		.Z(O3[12])
	);
	AO_CELL inst_4_12(
		.A1(out_sel[8]),
		.A2(I8[12]),
		.B1(out_sel[9]),
		.B2(I9[12]),
		.Z(O4[12])
	);
	AO_CELL inst_5_12(
		.A1(out_sel[10]),
		.A2(I10[12]),
		.B1(out_sel[11]),
		.B2(I11[12]),
		.Z(O5[12])
	);
	AO_CELL inst_6_12(
		.A1(out_sel[12]),
		.A2(I12[12]),
		.B1(out_sel[13]),
		.B2(I13[12]),
		.Z(O6[12])
	);
	AO_CELL inst_7_12(
		.A1(out_sel[14]),
		.A2(I14[12]),
		.B1(out_sel[15]),
		.B2(I15[12]),
		.Z(O7[12])
	);
	AO_CELL inst_0_13(
		.A1(out_sel[0]),
		.A2(I0[13]),
		.B1(out_sel[1]),
		.B2(I1[13]),
		.Z(O0[13])
	);
	AO_CELL inst_1_13(
		.A1(out_sel[2]),
		.A2(I2[13]),
		.B1(out_sel[3]),
		.B2(I3[13]),
		.Z(O1[13])
	);
	AO_CELL inst_2_13(
		.A1(out_sel[4]),
		.A2(I4[13]),
		.B1(out_sel[5]),
		.B2(I5[13]),
		.Z(O2[13])
	);
	AO_CELL inst_3_13(
		.A1(out_sel[6]),
		.A2(I6[13]),
		.B1(out_sel[7]),
		.B2(I7[13]),
		.Z(O3[13])
	);
	AO_CELL inst_4_13(
		.A1(out_sel[8]),
		.A2(I8[13]),
		.B1(out_sel[9]),
		.B2(I9[13]),
		.Z(O4[13])
	);
	AO_CELL inst_5_13(
		.A1(out_sel[10]),
		.A2(I10[13]),
		.B1(out_sel[11]),
		.B2(I11[13]),
		.Z(O5[13])
	);
	AO_CELL inst_6_13(
		.A1(out_sel[12]),
		.A2(I12[13]),
		.B1(out_sel[13]),
		.B2(I13[13]),
		.Z(O6[13])
	);
	AO_CELL inst_7_13(
		.A1(out_sel[14]),
		.A2(I14[13]),
		.B1(out_sel[15]),
		.B2(I15[13]),
		.Z(O7[13])
	);
	AO_CELL inst_0_14(
		.A1(out_sel[0]),
		.A2(I0[14]),
		.B1(out_sel[1]),
		.B2(I1[14]),
		.Z(O0[14])
	);
	AO_CELL inst_1_14(
		.A1(out_sel[2]),
		.A2(I2[14]),
		.B1(out_sel[3]),
		.B2(I3[14]),
		.Z(O1[14])
	);
	AO_CELL inst_2_14(
		.A1(out_sel[4]),
		.A2(I4[14]),
		.B1(out_sel[5]),
		.B2(I5[14]),
		.Z(O2[14])
	);
	AO_CELL inst_3_14(
		.A1(out_sel[6]),
		.A2(I6[14]),
		.B1(out_sel[7]),
		.B2(I7[14]),
		.Z(O3[14])
	);
	AO_CELL inst_4_14(
		.A1(out_sel[8]),
		.A2(I8[14]),
		.B1(out_sel[9]),
		.B2(I9[14]),
		.Z(O4[14])
	);
	AO_CELL inst_5_14(
		.A1(out_sel[10]),
		.A2(I10[14]),
		.B1(out_sel[11]),
		.B2(I11[14]),
		.Z(O5[14])
	);
	AO_CELL inst_6_14(
		.A1(out_sel[12]),
		.A2(I12[14]),
		.B1(out_sel[13]),
		.B2(I13[14]),
		.Z(O6[14])
	);
	AO_CELL inst_7_14(
		.A1(out_sel[14]),
		.A2(I14[14]),
		.B1(out_sel[15]),
		.B2(I15[14]),
		.Z(O7[14])
	);
	AO_CELL inst_0_15(
		.A1(out_sel[0]),
		.A2(I0[15]),
		.B1(out_sel[1]),
		.B2(I1[15]),
		.Z(O0[15])
	);
	AO_CELL inst_1_15(
		.A1(out_sel[2]),
		.A2(I2[15]),
		.B1(out_sel[3]),
		.B2(I3[15]),
		.Z(O1[15])
	);
	AO_CELL inst_2_15(
		.A1(out_sel[4]),
		.A2(I4[15]),
		.B1(out_sel[5]),
		.B2(I5[15]),
		.Z(O2[15])
	);
	AO_CELL inst_3_15(
		.A1(out_sel[6]),
		.A2(I6[15]),
		.B1(out_sel[7]),
		.B2(I7[15]),
		.Z(O3[15])
	);
	AO_CELL inst_4_15(
		.A1(out_sel[8]),
		.A2(I8[15]),
		.B1(out_sel[9]),
		.B2(I9[15]),
		.Z(O4[15])
	);
	AO_CELL inst_5_15(
		.A1(out_sel[10]),
		.A2(I10[15]),
		.B1(out_sel[11]),
		.B2(I11[15]),
		.Z(O5[15])
	);
	AO_CELL inst_6_15(
		.A1(out_sel[12]),
		.A2(I12[15]),
		.B1(out_sel[13]),
		.B2(I13[15]),
		.Z(O6[15])
	);
	AO_CELL inst_7_15(
		.A1(out_sel[14]),
		.A2(I14[15]),
		.B1(out_sel[15]),
		.B2(I15[15]),
		.Z(O7[15])
	);
	AO_CELL inst_0_16(
		.A1(out_sel[0]),
		.A2(I0[16]),
		.B1(out_sel[1]),
		.B2(I1[16]),
		.Z(O0[16])
	);
	AO_CELL inst_1_16(
		.A1(out_sel[2]),
		.A2(I2[16]),
		.B1(out_sel[3]),
		.B2(I3[16]),
		.Z(O1[16])
	);
	AO_CELL inst_2_16(
		.A1(out_sel[4]),
		.A2(I4[16]),
		.B1(out_sel[5]),
		.B2(I5[16]),
		.Z(O2[16])
	);
	AO_CELL inst_3_16(
		.A1(out_sel[6]),
		.A2(I6[16]),
		.B1(out_sel[7]),
		.B2(I7[16]),
		.Z(O3[16])
	);
	AO_CELL inst_4_16(
		.A1(out_sel[8]),
		.A2(I8[16]),
		.B1(out_sel[9]),
		.B2(I9[16]),
		.Z(O4[16])
	);
	AO_CELL inst_5_16(
		.A1(out_sel[10]),
		.A2(I10[16]),
		.B1(out_sel[11]),
		.B2(I11[16]),
		.Z(O5[16])
	);
	AO_CELL inst_6_16(
		.A1(out_sel[12]),
		.A2(I12[16]),
		.B1(out_sel[13]),
		.B2(I13[16]),
		.Z(O6[16])
	);
	AO_CELL inst_7_16(
		.A1(out_sel[14]),
		.A2(I14[16]),
		.B1(out_sel[15]),
		.B2(I15[16]),
		.Z(O7[16])
	);
	AO_CELL inst_0_17(
		.A1(out_sel[0]),
		.A2(I0[17]),
		.B1(out_sel[1]),
		.B2(I1[17]),
		.Z(O0[17])
	);
	AO_CELL inst_1_17(
		.A1(out_sel[2]),
		.A2(I2[17]),
		.B1(out_sel[3]),
		.B2(I3[17]),
		.Z(O1[17])
	);
	AO_CELL inst_2_17(
		.A1(out_sel[4]),
		.A2(I4[17]),
		.B1(out_sel[5]),
		.B2(I5[17]),
		.Z(O2[17])
	);
	AO_CELL inst_3_17(
		.A1(out_sel[6]),
		.A2(I6[17]),
		.B1(out_sel[7]),
		.B2(I7[17]),
		.Z(O3[17])
	);
	AO_CELL inst_4_17(
		.A1(out_sel[8]),
		.A2(I8[17]),
		.B1(out_sel[9]),
		.B2(I9[17]),
		.Z(O4[17])
	);
	AO_CELL inst_5_17(
		.A1(out_sel[10]),
		.A2(I10[17]),
		.B1(out_sel[11]),
		.B2(I11[17]),
		.Z(O5[17])
	);
	AO_CELL inst_6_17(
		.A1(out_sel[12]),
		.A2(I12[17]),
		.B1(out_sel[13]),
		.B2(I13[17]),
		.Z(O6[17])
	);
	AO_CELL inst_7_17(
		.A1(out_sel[14]),
		.A2(I14[17]),
		.B1(out_sel[15]),
		.B2(I15[17]),
		.Z(O7[17])
	);
	AO_CELL inst_0_18(
		.A1(out_sel[0]),
		.A2(I0[18]),
		.B1(out_sel[1]),
		.B2(I1[18]),
		.Z(O0[18])
	);
	AO_CELL inst_1_18(
		.A1(out_sel[2]),
		.A2(I2[18]),
		.B1(out_sel[3]),
		.B2(I3[18]),
		.Z(O1[18])
	);
	AO_CELL inst_2_18(
		.A1(out_sel[4]),
		.A2(I4[18]),
		.B1(out_sel[5]),
		.B2(I5[18]),
		.Z(O2[18])
	);
	AO_CELL inst_3_18(
		.A1(out_sel[6]),
		.A2(I6[18]),
		.B1(out_sel[7]),
		.B2(I7[18]),
		.Z(O3[18])
	);
	AO_CELL inst_4_18(
		.A1(out_sel[8]),
		.A2(I8[18]),
		.B1(out_sel[9]),
		.B2(I9[18]),
		.Z(O4[18])
	);
	AO_CELL inst_5_18(
		.A1(out_sel[10]),
		.A2(I10[18]),
		.B1(out_sel[11]),
		.B2(I11[18]),
		.Z(O5[18])
	);
	AO_CELL inst_6_18(
		.A1(out_sel[12]),
		.A2(I12[18]),
		.B1(out_sel[13]),
		.B2(I13[18]),
		.Z(O6[18])
	);
	AO_CELL inst_7_18(
		.A1(out_sel[14]),
		.A2(I14[18]),
		.B1(out_sel[15]),
		.B2(I15[18]),
		.Z(O7[18])
	);
	AO_CELL inst_0_19(
		.A1(out_sel[0]),
		.A2(I0[19]),
		.B1(out_sel[1]),
		.B2(I1[19]),
		.Z(O0[19])
	);
	AO_CELL inst_1_19(
		.A1(out_sel[2]),
		.A2(I2[19]),
		.B1(out_sel[3]),
		.B2(I3[19]),
		.Z(O1[19])
	);
	AO_CELL inst_2_19(
		.A1(out_sel[4]),
		.A2(I4[19]),
		.B1(out_sel[5]),
		.B2(I5[19]),
		.Z(O2[19])
	);
	AO_CELL inst_3_19(
		.A1(out_sel[6]),
		.A2(I6[19]),
		.B1(out_sel[7]),
		.B2(I7[19]),
		.Z(O3[19])
	);
	AO_CELL inst_4_19(
		.A1(out_sel[8]),
		.A2(I8[19]),
		.B1(out_sel[9]),
		.B2(I9[19]),
		.Z(O4[19])
	);
	AO_CELL inst_5_19(
		.A1(out_sel[10]),
		.A2(I10[19]),
		.B1(out_sel[11]),
		.B2(I11[19]),
		.Z(O5[19])
	);
	AO_CELL inst_6_19(
		.A1(out_sel[12]),
		.A2(I12[19]),
		.B1(out_sel[13]),
		.B2(I13[19]),
		.Z(O6[19])
	);
	AO_CELL inst_7_19(
		.A1(out_sel[14]),
		.A2(I14[19]),
		.B1(out_sel[15]),
		.B2(I15[19]),
		.Z(O7[19])
	);
	AO_CELL inst_0_20(
		.A1(out_sel[0]),
		.A2(I0[20]),
		.B1(out_sel[1]),
		.B2(I1[20]),
		.Z(O0[20])
	);
	AO_CELL inst_1_20(
		.A1(out_sel[2]),
		.A2(I2[20]),
		.B1(out_sel[3]),
		.B2(I3[20]),
		.Z(O1[20])
	);
	AO_CELL inst_2_20(
		.A1(out_sel[4]),
		.A2(I4[20]),
		.B1(out_sel[5]),
		.B2(I5[20]),
		.Z(O2[20])
	);
	AO_CELL inst_3_20(
		.A1(out_sel[6]),
		.A2(I6[20]),
		.B1(out_sel[7]),
		.B2(I7[20]),
		.Z(O3[20])
	);
	AO_CELL inst_4_20(
		.A1(out_sel[8]),
		.A2(I8[20]),
		.B1(out_sel[9]),
		.B2(I9[20]),
		.Z(O4[20])
	);
	AO_CELL inst_5_20(
		.A1(out_sel[10]),
		.A2(I10[20]),
		.B1(out_sel[11]),
		.B2(I11[20]),
		.Z(O5[20])
	);
	AO_CELL inst_6_20(
		.A1(out_sel[12]),
		.A2(I12[20]),
		.B1(out_sel[13]),
		.B2(I13[20]),
		.Z(O6[20])
	);
	AO_CELL inst_7_20(
		.A1(out_sel[14]),
		.A2(I14[20]),
		.B1(out_sel[15]),
		.B2(I15[20]),
		.Z(O7[20])
	);
	AO_CELL inst_0_21(
		.A1(out_sel[0]),
		.A2(I0[21]),
		.B1(out_sel[1]),
		.B2(I1[21]),
		.Z(O0[21])
	);
	AO_CELL inst_1_21(
		.A1(out_sel[2]),
		.A2(I2[21]),
		.B1(out_sel[3]),
		.B2(I3[21]),
		.Z(O1[21])
	);
	AO_CELL inst_2_21(
		.A1(out_sel[4]),
		.A2(I4[21]),
		.B1(out_sel[5]),
		.B2(I5[21]),
		.Z(O2[21])
	);
	AO_CELL inst_3_21(
		.A1(out_sel[6]),
		.A2(I6[21]),
		.B1(out_sel[7]),
		.B2(I7[21]),
		.Z(O3[21])
	);
	AO_CELL inst_4_21(
		.A1(out_sel[8]),
		.A2(I8[21]),
		.B1(out_sel[9]),
		.B2(I9[21]),
		.Z(O4[21])
	);
	AO_CELL inst_5_21(
		.A1(out_sel[10]),
		.A2(I10[21]),
		.B1(out_sel[11]),
		.B2(I11[21]),
		.Z(O5[21])
	);
	AO_CELL inst_6_21(
		.A1(out_sel[12]),
		.A2(I12[21]),
		.B1(out_sel[13]),
		.B2(I13[21]),
		.Z(O6[21])
	);
	AO_CELL inst_7_21(
		.A1(out_sel[14]),
		.A2(I14[21]),
		.B1(out_sel[15]),
		.B2(I15[21]),
		.Z(O7[21])
	);
	AO_CELL inst_0_22(
		.A1(out_sel[0]),
		.A2(I0[22]),
		.B1(out_sel[1]),
		.B2(I1[22]),
		.Z(O0[22])
	);
	AO_CELL inst_1_22(
		.A1(out_sel[2]),
		.A2(I2[22]),
		.B1(out_sel[3]),
		.B2(I3[22]),
		.Z(O1[22])
	);
	AO_CELL inst_2_22(
		.A1(out_sel[4]),
		.A2(I4[22]),
		.B1(out_sel[5]),
		.B2(I5[22]),
		.Z(O2[22])
	);
	AO_CELL inst_3_22(
		.A1(out_sel[6]),
		.A2(I6[22]),
		.B1(out_sel[7]),
		.B2(I7[22]),
		.Z(O3[22])
	);
	AO_CELL inst_4_22(
		.A1(out_sel[8]),
		.A2(I8[22]),
		.B1(out_sel[9]),
		.B2(I9[22]),
		.Z(O4[22])
	);
	AO_CELL inst_5_22(
		.A1(out_sel[10]),
		.A2(I10[22]),
		.B1(out_sel[11]),
		.B2(I11[22]),
		.Z(O5[22])
	);
	AO_CELL inst_6_22(
		.A1(out_sel[12]),
		.A2(I12[22]),
		.B1(out_sel[13]),
		.B2(I13[22]),
		.Z(O6[22])
	);
	AO_CELL inst_7_22(
		.A1(out_sel[14]),
		.A2(I14[22]),
		.B1(out_sel[15]),
		.B2(I15[22]),
		.Z(O7[22])
	);
	AO_CELL inst_0_23(
		.A1(out_sel[0]),
		.A2(I0[23]),
		.B1(out_sel[1]),
		.B2(I1[23]),
		.Z(O0[23])
	);
	AO_CELL inst_1_23(
		.A1(out_sel[2]),
		.A2(I2[23]),
		.B1(out_sel[3]),
		.B2(I3[23]),
		.Z(O1[23])
	);
	AO_CELL inst_2_23(
		.A1(out_sel[4]),
		.A2(I4[23]),
		.B1(out_sel[5]),
		.B2(I5[23]),
		.Z(O2[23])
	);
	AO_CELL inst_3_23(
		.A1(out_sel[6]),
		.A2(I6[23]),
		.B1(out_sel[7]),
		.B2(I7[23]),
		.Z(O3[23])
	);
	AO_CELL inst_4_23(
		.A1(out_sel[8]),
		.A2(I8[23]),
		.B1(out_sel[9]),
		.B2(I9[23]),
		.Z(O4[23])
	);
	AO_CELL inst_5_23(
		.A1(out_sel[10]),
		.A2(I10[23]),
		.B1(out_sel[11]),
		.B2(I11[23]),
		.Z(O5[23])
	);
	AO_CELL inst_6_23(
		.A1(out_sel[12]),
		.A2(I12[23]),
		.B1(out_sel[13]),
		.B2(I13[23]),
		.Z(O6[23])
	);
	AO_CELL inst_7_23(
		.A1(out_sel[14]),
		.A2(I14[23]),
		.B1(out_sel[15]),
		.B2(I15[23]),
		.Z(O7[23])
	);
	AO_CELL inst_0_24(
		.A1(out_sel[0]),
		.A2(I0[24]),
		.B1(out_sel[1]),
		.B2(I1[24]),
		.Z(O0[24])
	);
	AO_CELL inst_1_24(
		.A1(out_sel[2]),
		.A2(I2[24]),
		.B1(out_sel[3]),
		.B2(I3[24]),
		.Z(O1[24])
	);
	AO_CELL inst_2_24(
		.A1(out_sel[4]),
		.A2(I4[24]),
		.B1(out_sel[5]),
		.B2(I5[24]),
		.Z(O2[24])
	);
	AO_CELL inst_3_24(
		.A1(out_sel[6]),
		.A2(I6[24]),
		.B1(out_sel[7]),
		.B2(I7[24]),
		.Z(O3[24])
	);
	AO_CELL inst_4_24(
		.A1(out_sel[8]),
		.A2(I8[24]),
		.B1(out_sel[9]),
		.B2(I9[24]),
		.Z(O4[24])
	);
	AO_CELL inst_5_24(
		.A1(out_sel[10]),
		.A2(I10[24]),
		.B1(out_sel[11]),
		.B2(I11[24]),
		.Z(O5[24])
	);
	AO_CELL inst_6_24(
		.A1(out_sel[12]),
		.A2(I12[24]),
		.B1(out_sel[13]),
		.B2(I13[24]),
		.Z(O6[24])
	);
	AO_CELL inst_7_24(
		.A1(out_sel[14]),
		.A2(I14[24]),
		.B1(out_sel[15]),
		.B2(I15[24]),
		.Z(O7[24])
	);
	AO_CELL inst_0_25(
		.A1(out_sel[0]),
		.A2(I0[25]),
		.B1(out_sel[1]),
		.B2(I1[25]),
		.Z(O0[25])
	);
	AO_CELL inst_1_25(
		.A1(out_sel[2]),
		.A2(I2[25]),
		.B1(out_sel[3]),
		.B2(I3[25]),
		.Z(O1[25])
	);
	AO_CELL inst_2_25(
		.A1(out_sel[4]),
		.A2(I4[25]),
		.B1(out_sel[5]),
		.B2(I5[25]),
		.Z(O2[25])
	);
	AO_CELL inst_3_25(
		.A1(out_sel[6]),
		.A2(I6[25]),
		.B1(out_sel[7]),
		.B2(I7[25]),
		.Z(O3[25])
	);
	AO_CELL inst_4_25(
		.A1(out_sel[8]),
		.A2(I8[25]),
		.B1(out_sel[9]),
		.B2(I9[25]),
		.Z(O4[25])
	);
	AO_CELL inst_5_25(
		.A1(out_sel[10]),
		.A2(I10[25]),
		.B1(out_sel[11]),
		.B2(I11[25]),
		.Z(O5[25])
	);
	AO_CELL inst_6_25(
		.A1(out_sel[12]),
		.A2(I12[25]),
		.B1(out_sel[13]),
		.B2(I13[25]),
		.Z(O6[25])
	);
	AO_CELL inst_7_25(
		.A1(out_sel[14]),
		.A2(I14[25]),
		.B1(out_sel[15]),
		.B2(I15[25]),
		.Z(O7[25])
	);
	AO_CELL inst_0_26(
		.A1(out_sel[0]),
		.A2(I0[26]),
		.B1(out_sel[1]),
		.B2(I1[26]),
		.Z(O0[26])
	);
	AO_CELL inst_1_26(
		.A1(out_sel[2]),
		.A2(I2[26]),
		.B1(out_sel[3]),
		.B2(I3[26]),
		.Z(O1[26])
	);
	AO_CELL inst_2_26(
		.A1(out_sel[4]),
		.A2(I4[26]),
		.B1(out_sel[5]),
		.B2(I5[26]),
		.Z(O2[26])
	);
	AO_CELL inst_3_26(
		.A1(out_sel[6]),
		.A2(I6[26]),
		.B1(out_sel[7]),
		.B2(I7[26]),
		.Z(O3[26])
	);
	AO_CELL inst_4_26(
		.A1(out_sel[8]),
		.A2(I8[26]),
		.B1(out_sel[9]),
		.B2(I9[26]),
		.Z(O4[26])
	);
	AO_CELL inst_5_26(
		.A1(out_sel[10]),
		.A2(I10[26]),
		.B1(out_sel[11]),
		.B2(I11[26]),
		.Z(O5[26])
	);
	AO_CELL inst_6_26(
		.A1(out_sel[12]),
		.A2(I12[26]),
		.B1(out_sel[13]),
		.B2(I13[26]),
		.Z(O6[26])
	);
	AO_CELL inst_7_26(
		.A1(out_sel[14]),
		.A2(I14[26]),
		.B1(out_sel[15]),
		.B2(I15[26]),
		.Z(O7[26])
	);
	AO_CELL inst_0_27(
		.A1(out_sel[0]),
		.A2(I0[27]),
		.B1(out_sel[1]),
		.B2(I1[27]),
		.Z(O0[27])
	);
	AO_CELL inst_1_27(
		.A1(out_sel[2]),
		.A2(I2[27]),
		.B1(out_sel[3]),
		.B2(I3[27]),
		.Z(O1[27])
	);
	AO_CELL inst_2_27(
		.A1(out_sel[4]),
		.A2(I4[27]),
		.B1(out_sel[5]),
		.B2(I5[27]),
		.Z(O2[27])
	);
	AO_CELL inst_3_27(
		.A1(out_sel[6]),
		.A2(I6[27]),
		.B1(out_sel[7]),
		.B2(I7[27]),
		.Z(O3[27])
	);
	AO_CELL inst_4_27(
		.A1(out_sel[8]),
		.A2(I8[27]),
		.B1(out_sel[9]),
		.B2(I9[27]),
		.Z(O4[27])
	);
	AO_CELL inst_5_27(
		.A1(out_sel[10]),
		.A2(I10[27]),
		.B1(out_sel[11]),
		.B2(I11[27]),
		.Z(O5[27])
	);
	AO_CELL inst_6_27(
		.A1(out_sel[12]),
		.A2(I12[27]),
		.B1(out_sel[13]),
		.B2(I13[27]),
		.Z(O6[27])
	);
	AO_CELL inst_7_27(
		.A1(out_sel[14]),
		.A2(I14[27]),
		.B1(out_sel[15]),
		.B2(I15[27]),
		.Z(O7[27])
	);
	AO_CELL inst_0_28(
		.A1(out_sel[0]),
		.A2(I0[28]),
		.B1(out_sel[1]),
		.B2(I1[28]),
		.Z(O0[28])
	);
	AO_CELL inst_1_28(
		.A1(out_sel[2]),
		.A2(I2[28]),
		.B1(out_sel[3]),
		.B2(I3[28]),
		.Z(O1[28])
	);
	AO_CELL inst_2_28(
		.A1(out_sel[4]),
		.A2(I4[28]),
		.B1(out_sel[5]),
		.B2(I5[28]),
		.Z(O2[28])
	);
	AO_CELL inst_3_28(
		.A1(out_sel[6]),
		.A2(I6[28]),
		.B1(out_sel[7]),
		.B2(I7[28]),
		.Z(O3[28])
	);
	AO_CELL inst_4_28(
		.A1(out_sel[8]),
		.A2(I8[28]),
		.B1(out_sel[9]),
		.B2(I9[28]),
		.Z(O4[28])
	);
	AO_CELL inst_5_28(
		.A1(out_sel[10]),
		.A2(I10[28]),
		.B1(out_sel[11]),
		.B2(I11[28]),
		.Z(O5[28])
	);
	AO_CELL inst_6_28(
		.A1(out_sel[12]),
		.A2(I12[28]),
		.B1(out_sel[13]),
		.B2(I13[28]),
		.Z(O6[28])
	);
	AO_CELL inst_7_28(
		.A1(out_sel[14]),
		.A2(I14[28]),
		.B1(out_sel[15]),
		.B2(I15[28]),
		.Z(O7[28])
	);
	AO_CELL inst_0_29(
		.A1(out_sel[0]),
		.A2(I0[29]),
		.B1(out_sel[1]),
		.B2(I1[29]),
		.Z(O0[29])
	);
	AO_CELL inst_1_29(
		.A1(out_sel[2]),
		.A2(I2[29]),
		.B1(out_sel[3]),
		.B2(I3[29]),
		.Z(O1[29])
	);
	AO_CELL inst_2_29(
		.A1(out_sel[4]),
		.A2(I4[29]),
		.B1(out_sel[5]),
		.B2(I5[29]),
		.Z(O2[29])
	);
	AO_CELL inst_3_29(
		.A1(out_sel[6]),
		.A2(I6[29]),
		.B1(out_sel[7]),
		.B2(I7[29]),
		.Z(O3[29])
	);
	AO_CELL inst_4_29(
		.A1(out_sel[8]),
		.A2(I8[29]),
		.B1(out_sel[9]),
		.B2(I9[29]),
		.Z(O4[29])
	);
	AO_CELL inst_5_29(
		.A1(out_sel[10]),
		.A2(I10[29]),
		.B1(out_sel[11]),
		.B2(I11[29]),
		.Z(O5[29])
	);
	AO_CELL inst_6_29(
		.A1(out_sel[12]),
		.A2(I12[29]),
		.B1(out_sel[13]),
		.B2(I13[29]),
		.Z(O6[29])
	);
	AO_CELL inst_7_29(
		.A1(out_sel[14]),
		.A2(I14[29]),
		.B1(out_sel[15]),
		.B2(I15[29]),
		.Z(O7[29])
	);
	AO_CELL inst_0_30(
		.A1(out_sel[0]),
		.A2(I0[30]),
		.B1(out_sel[1]),
		.B2(I1[30]),
		.Z(O0[30])
	);
	AO_CELL inst_1_30(
		.A1(out_sel[2]),
		.A2(I2[30]),
		.B1(out_sel[3]),
		.B2(I3[30]),
		.Z(O1[30])
	);
	AO_CELL inst_2_30(
		.A1(out_sel[4]),
		.A2(I4[30]),
		.B1(out_sel[5]),
		.B2(I5[30]),
		.Z(O2[30])
	);
	AO_CELL inst_3_30(
		.A1(out_sel[6]),
		.A2(I6[30]),
		.B1(out_sel[7]),
		.B2(I7[30]),
		.Z(O3[30])
	);
	AO_CELL inst_4_30(
		.A1(out_sel[8]),
		.A2(I8[30]),
		.B1(out_sel[9]),
		.B2(I9[30]),
		.Z(O4[30])
	);
	AO_CELL inst_5_30(
		.A1(out_sel[10]),
		.A2(I10[30]),
		.B1(out_sel[11]),
		.B2(I11[30]),
		.Z(O5[30])
	);
	AO_CELL inst_6_30(
		.A1(out_sel[12]),
		.A2(I12[30]),
		.B1(out_sel[13]),
		.B2(I13[30]),
		.Z(O6[30])
	);
	AO_CELL inst_7_30(
		.A1(out_sel[14]),
		.A2(I14[30]),
		.B1(out_sel[15]),
		.B2(I15[30]),
		.Z(O7[30])
	);
	AO_CELL inst_0_31(
		.A1(out_sel[0]),
		.A2(I0[31]),
		.B1(out_sel[1]),
		.B2(I1[31]),
		.Z(O0[31])
	);
	AO_CELL inst_1_31(
		.A1(out_sel[2]),
		.A2(I2[31]),
		.B1(out_sel[3]),
		.B2(I3[31]),
		.Z(O1[31])
	);
	AO_CELL inst_2_31(
		.A1(out_sel[4]),
		.A2(I4[31]),
		.B1(out_sel[5]),
		.B2(I5[31]),
		.Z(O2[31])
	);
	AO_CELL inst_3_31(
		.A1(out_sel[6]),
		.A2(I6[31]),
		.B1(out_sel[7]),
		.B2(I7[31]),
		.Z(O3[31])
	);
	AO_CELL inst_4_31(
		.A1(out_sel[8]),
		.A2(I8[31]),
		.B1(out_sel[9]),
		.B2(I9[31]),
		.Z(O4[31])
	);
	AO_CELL inst_5_31(
		.A1(out_sel[10]),
		.A2(I10[31]),
		.B1(out_sel[11]),
		.B2(I11[31]),
		.Z(O5[31])
	);
	AO_CELL inst_6_31(
		.A1(out_sel[12]),
		.A2(I12[31]),
		.B1(out_sel[13]),
		.B2(I13[31]),
		.Z(O6[31])
	);
	AO_CELL inst_7_31(
		.A1(out_sel[14]),
		.A2(I14[31]),
		.B1(out_sel[15]),
		.B2(I15[31]),
		.Z(O7[31])
	);
endmodule
module mux_aoi_13_32 (
	I,
	S,
	out_sel,
	O
);
	input wire [415:0] I;
	input wire [3:0] S;
	output wire [15:0] out_sel;
	output wire [31:0] O;
	wire [31:0] O_int0;
	wire [31:0] O_int1;
	wire [31:0] O_int2;
	wire [31:0] O_int3;
	wire [31:0] O_int4;
	wire [31:0] O_int5;
	wire [31:0] O_int6;
	precoder_32_13 u_precoder(
		.S(S),
		.out_sel(out_sel)
	);
	mux_logic_32_13 u_mux_logic(
		.I0(I[0+:32]),
		.I1(I[32+:32]),
		.I2(I[64+:32]),
		.I3(I[96+:32]),
		.I4(I[128+:32]),
		.I5(I[160+:32]),
		.I6(I[192+:32]),
		.I7(I[224+:32]),
		.I8(I[256+:32]),
		.I9(I[288+:32]),
		.I10(I[320+:32]),
		.I11(I[352+:32]),
		.I12(I[384+:32]),
		.out_sel(out_sel),
		.O0(O_int0),
		.O1(O_int1),
		.O2(O_int2),
		.O3(O_int3),
		.O4(O_int4),
		.O5(O_int5),
		.O6(O_int6)
	);
	assign O = (((((O_int0 | O_int1) | O_int2) | O_int3) | O_int4) | O_int5) | O_int6;
endmodule
module precoder_32_13 (
	S,
	out_sel
);
	input wire [3:0] S;
	output reg [15:0] out_sel;
	always @(*) begin : mux_sel
		case (S)
			4'd0: out_sel = 16'b0000000000000001;
			4'd1: out_sel = 16'b0000000000000010;
			4'd2: out_sel = 16'b0000000000000100;
			4'd3: out_sel = 16'b0000000000001000;
			4'd4: out_sel = 16'b0000000000010000;
			4'd5: out_sel = 16'b0000000000100000;
			4'd6: out_sel = 16'b0000000001000000;
			4'd7: out_sel = 16'b0000000010000000;
			4'd8: out_sel = 16'b0000000100000000;
			4'd9: out_sel = 16'b0000001000000000;
			4'd10: out_sel = 16'b0000010000000000;
			4'd11: out_sel = 16'b0000100000000000;
			4'd12: out_sel = 16'b0001000000000000;
			default: out_sel = 16'b0000000000000000;
		endcase
	end
endmodule
module mux_logic_32_13 (
	out_sel,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	I9,
	I10,
	I11,
	I12,
	O0,
	O1,
	O2,
	O3,
	O4,
	O5,
	O6
);
	input wire [15:0] out_sel;
	input wire [31:0] I0;
	input wire [31:0] I1;
	input wire [31:0] I2;
	input wire [31:0] I3;
	input wire [31:0] I4;
	input wire [31:0] I5;
	input wire [31:0] I6;
	input wire [31:0] I7;
	input wire [31:0] I8;
	input wire [31:0] I9;
	input wire [31:0] I10;
	input wire [31:0] I11;
	input wire [31:0] I12;
	output wire [31:0] O0;
	output wire [31:0] O1;
	output wire [31:0] O2;
	output wire [31:0] O3;
	output wire [31:0] O4;
	output wire [31:0] O5;
	output wire [31:0] O6;
	AO_CELL inst_0_0(
		.A1(out_sel[0]),
		.A2(I0[0]),
		.B1(out_sel[1]),
		.B2(I1[0]),
		.Z(O0[0])
	);
	AO_CELL inst_1_0(
		.A1(out_sel[2]),
		.A2(I2[0]),
		.B1(out_sel[3]),
		.B2(I3[0]),
		.Z(O1[0])
	);
	AO_CELL inst_2_0(
		.A1(out_sel[4]),
		.A2(I4[0]),
		.B1(out_sel[5]),
		.B2(I5[0]),
		.Z(O2[0])
	);
	AO_CELL inst_3_0(
		.A1(out_sel[6]),
		.A2(I6[0]),
		.B1(out_sel[7]),
		.B2(I7[0]),
		.Z(O3[0])
	);
	AO_CELL inst_4_0(
		.A1(out_sel[8]),
		.A2(I8[0]),
		.B1(out_sel[9]),
		.B2(I9[0]),
		.Z(O4[0])
	);
	AO_CELL inst_5_0(
		.A1(out_sel[10]),
		.A2(I10[0]),
		.B1(out_sel[11]),
		.B2(I11[0]),
		.Z(O5[0])
	);
	AN_CELL inst_and_0(
		.A1(out_sel[12]),
		.A2(I12[0]),
		.Z(O6[0])
	);
	AO_CELL inst_0_1(
		.A1(out_sel[0]),
		.A2(I0[1]),
		.B1(out_sel[1]),
		.B2(I1[1]),
		.Z(O0[1])
	);
	AO_CELL inst_1_1(
		.A1(out_sel[2]),
		.A2(I2[1]),
		.B1(out_sel[3]),
		.B2(I3[1]),
		.Z(O1[1])
	);
	AO_CELL inst_2_1(
		.A1(out_sel[4]),
		.A2(I4[1]),
		.B1(out_sel[5]),
		.B2(I5[1]),
		.Z(O2[1])
	);
	AO_CELL inst_3_1(
		.A1(out_sel[6]),
		.A2(I6[1]),
		.B1(out_sel[7]),
		.B2(I7[1]),
		.Z(O3[1])
	);
	AO_CELL inst_4_1(
		.A1(out_sel[8]),
		.A2(I8[1]),
		.B1(out_sel[9]),
		.B2(I9[1]),
		.Z(O4[1])
	);
	AO_CELL inst_5_1(
		.A1(out_sel[10]),
		.A2(I10[1]),
		.B1(out_sel[11]),
		.B2(I11[1]),
		.Z(O5[1])
	);
	AN_CELL inst_and_1(
		.A1(out_sel[12]),
		.A2(I12[1]),
		.Z(O6[1])
	);
	AO_CELL inst_0_2(
		.A1(out_sel[0]),
		.A2(I0[2]),
		.B1(out_sel[1]),
		.B2(I1[2]),
		.Z(O0[2])
	);
	AO_CELL inst_1_2(
		.A1(out_sel[2]),
		.A2(I2[2]),
		.B1(out_sel[3]),
		.B2(I3[2]),
		.Z(O1[2])
	);
	AO_CELL inst_2_2(
		.A1(out_sel[4]),
		.A2(I4[2]),
		.B1(out_sel[5]),
		.B2(I5[2]),
		.Z(O2[2])
	);
	AO_CELL inst_3_2(
		.A1(out_sel[6]),
		.A2(I6[2]),
		.B1(out_sel[7]),
		.B2(I7[2]),
		.Z(O3[2])
	);
	AO_CELL inst_4_2(
		.A1(out_sel[8]),
		.A2(I8[2]),
		.B1(out_sel[9]),
		.B2(I9[2]),
		.Z(O4[2])
	);
	AO_CELL inst_5_2(
		.A1(out_sel[10]),
		.A2(I10[2]),
		.B1(out_sel[11]),
		.B2(I11[2]),
		.Z(O5[2])
	);
	AN_CELL inst_and_2(
		.A1(out_sel[12]),
		.A2(I12[2]),
		.Z(O6[2])
	);
	AO_CELL inst_0_3(
		.A1(out_sel[0]),
		.A2(I0[3]),
		.B1(out_sel[1]),
		.B2(I1[3]),
		.Z(O0[3])
	);
	AO_CELL inst_1_3(
		.A1(out_sel[2]),
		.A2(I2[3]),
		.B1(out_sel[3]),
		.B2(I3[3]),
		.Z(O1[3])
	);
	AO_CELL inst_2_3(
		.A1(out_sel[4]),
		.A2(I4[3]),
		.B1(out_sel[5]),
		.B2(I5[3]),
		.Z(O2[3])
	);
	AO_CELL inst_3_3(
		.A1(out_sel[6]),
		.A2(I6[3]),
		.B1(out_sel[7]),
		.B2(I7[3]),
		.Z(O3[3])
	);
	AO_CELL inst_4_3(
		.A1(out_sel[8]),
		.A2(I8[3]),
		.B1(out_sel[9]),
		.B2(I9[3]),
		.Z(O4[3])
	);
	AO_CELL inst_5_3(
		.A1(out_sel[10]),
		.A2(I10[3]),
		.B1(out_sel[11]),
		.B2(I11[3]),
		.Z(O5[3])
	);
	AN_CELL inst_and_3(
		.A1(out_sel[12]),
		.A2(I12[3]),
		.Z(O6[3])
	);
	AO_CELL inst_0_4(
		.A1(out_sel[0]),
		.A2(I0[4]),
		.B1(out_sel[1]),
		.B2(I1[4]),
		.Z(O0[4])
	);
	AO_CELL inst_1_4(
		.A1(out_sel[2]),
		.A2(I2[4]),
		.B1(out_sel[3]),
		.B2(I3[4]),
		.Z(O1[4])
	);
	AO_CELL inst_2_4(
		.A1(out_sel[4]),
		.A2(I4[4]),
		.B1(out_sel[5]),
		.B2(I5[4]),
		.Z(O2[4])
	);
	AO_CELL inst_3_4(
		.A1(out_sel[6]),
		.A2(I6[4]),
		.B1(out_sel[7]),
		.B2(I7[4]),
		.Z(O3[4])
	);
	AO_CELL inst_4_4(
		.A1(out_sel[8]),
		.A2(I8[4]),
		.B1(out_sel[9]),
		.B2(I9[4]),
		.Z(O4[4])
	);
	AO_CELL inst_5_4(
		.A1(out_sel[10]),
		.A2(I10[4]),
		.B1(out_sel[11]),
		.B2(I11[4]),
		.Z(O5[4])
	);
	AN_CELL inst_and_4(
		.A1(out_sel[12]),
		.A2(I12[4]),
		.Z(O6[4])
	);
	AO_CELL inst_0_5(
		.A1(out_sel[0]),
		.A2(I0[5]),
		.B1(out_sel[1]),
		.B2(I1[5]),
		.Z(O0[5])
	);
	AO_CELL inst_1_5(
		.A1(out_sel[2]),
		.A2(I2[5]),
		.B1(out_sel[3]),
		.B2(I3[5]),
		.Z(O1[5])
	);
	AO_CELL inst_2_5(
		.A1(out_sel[4]),
		.A2(I4[5]),
		.B1(out_sel[5]),
		.B2(I5[5]),
		.Z(O2[5])
	);
	AO_CELL inst_3_5(
		.A1(out_sel[6]),
		.A2(I6[5]),
		.B1(out_sel[7]),
		.B2(I7[5]),
		.Z(O3[5])
	);
	AO_CELL inst_4_5(
		.A1(out_sel[8]),
		.A2(I8[5]),
		.B1(out_sel[9]),
		.B2(I9[5]),
		.Z(O4[5])
	);
	AO_CELL inst_5_5(
		.A1(out_sel[10]),
		.A2(I10[5]),
		.B1(out_sel[11]),
		.B2(I11[5]),
		.Z(O5[5])
	);
	AN_CELL inst_and_5(
		.A1(out_sel[12]),
		.A2(I12[5]),
		.Z(O6[5])
	);
	AO_CELL inst_0_6(
		.A1(out_sel[0]),
		.A2(I0[6]),
		.B1(out_sel[1]),
		.B2(I1[6]),
		.Z(O0[6])
	);
	AO_CELL inst_1_6(
		.A1(out_sel[2]),
		.A2(I2[6]),
		.B1(out_sel[3]),
		.B2(I3[6]),
		.Z(O1[6])
	);
	AO_CELL inst_2_6(
		.A1(out_sel[4]),
		.A2(I4[6]),
		.B1(out_sel[5]),
		.B2(I5[6]),
		.Z(O2[6])
	);
	AO_CELL inst_3_6(
		.A1(out_sel[6]),
		.A2(I6[6]),
		.B1(out_sel[7]),
		.B2(I7[6]),
		.Z(O3[6])
	);
	AO_CELL inst_4_6(
		.A1(out_sel[8]),
		.A2(I8[6]),
		.B1(out_sel[9]),
		.B2(I9[6]),
		.Z(O4[6])
	);
	AO_CELL inst_5_6(
		.A1(out_sel[10]),
		.A2(I10[6]),
		.B1(out_sel[11]),
		.B2(I11[6]),
		.Z(O5[6])
	);
	AN_CELL inst_and_6(
		.A1(out_sel[12]),
		.A2(I12[6]),
		.Z(O6[6])
	);
	AO_CELL inst_0_7(
		.A1(out_sel[0]),
		.A2(I0[7]),
		.B1(out_sel[1]),
		.B2(I1[7]),
		.Z(O0[7])
	);
	AO_CELL inst_1_7(
		.A1(out_sel[2]),
		.A2(I2[7]),
		.B1(out_sel[3]),
		.B2(I3[7]),
		.Z(O1[7])
	);
	AO_CELL inst_2_7(
		.A1(out_sel[4]),
		.A2(I4[7]),
		.B1(out_sel[5]),
		.B2(I5[7]),
		.Z(O2[7])
	);
	AO_CELL inst_3_7(
		.A1(out_sel[6]),
		.A2(I6[7]),
		.B1(out_sel[7]),
		.B2(I7[7]),
		.Z(O3[7])
	);
	AO_CELL inst_4_7(
		.A1(out_sel[8]),
		.A2(I8[7]),
		.B1(out_sel[9]),
		.B2(I9[7]),
		.Z(O4[7])
	);
	AO_CELL inst_5_7(
		.A1(out_sel[10]),
		.A2(I10[7]),
		.B1(out_sel[11]),
		.B2(I11[7]),
		.Z(O5[7])
	);
	AN_CELL inst_and_7(
		.A1(out_sel[12]),
		.A2(I12[7]),
		.Z(O6[7])
	);
	AO_CELL inst_0_8(
		.A1(out_sel[0]),
		.A2(I0[8]),
		.B1(out_sel[1]),
		.B2(I1[8]),
		.Z(O0[8])
	);
	AO_CELL inst_1_8(
		.A1(out_sel[2]),
		.A2(I2[8]),
		.B1(out_sel[3]),
		.B2(I3[8]),
		.Z(O1[8])
	);
	AO_CELL inst_2_8(
		.A1(out_sel[4]),
		.A2(I4[8]),
		.B1(out_sel[5]),
		.B2(I5[8]),
		.Z(O2[8])
	);
	AO_CELL inst_3_8(
		.A1(out_sel[6]),
		.A2(I6[8]),
		.B1(out_sel[7]),
		.B2(I7[8]),
		.Z(O3[8])
	);
	AO_CELL inst_4_8(
		.A1(out_sel[8]),
		.A2(I8[8]),
		.B1(out_sel[9]),
		.B2(I9[8]),
		.Z(O4[8])
	);
	AO_CELL inst_5_8(
		.A1(out_sel[10]),
		.A2(I10[8]),
		.B1(out_sel[11]),
		.B2(I11[8]),
		.Z(O5[8])
	);
	AN_CELL inst_and_8(
		.A1(out_sel[12]),
		.A2(I12[8]),
		.Z(O6[8])
	);
	AO_CELL inst_0_9(
		.A1(out_sel[0]),
		.A2(I0[9]),
		.B1(out_sel[1]),
		.B2(I1[9]),
		.Z(O0[9])
	);
	AO_CELL inst_1_9(
		.A1(out_sel[2]),
		.A2(I2[9]),
		.B1(out_sel[3]),
		.B2(I3[9]),
		.Z(O1[9])
	);
	AO_CELL inst_2_9(
		.A1(out_sel[4]),
		.A2(I4[9]),
		.B1(out_sel[5]),
		.B2(I5[9]),
		.Z(O2[9])
	);
	AO_CELL inst_3_9(
		.A1(out_sel[6]),
		.A2(I6[9]),
		.B1(out_sel[7]),
		.B2(I7[9]),
		.Z(O3[9])
	);
	AO_CELL inst_4_9(
		.A1(out_sel[8]),
		.A2(I8[9]),
		.B1(out_sel[9]),
		.B2(I9[9]),
		.Z(O4[9])
	);
	AO_CELL inst_5_9(
		.A1(out_sel[10]),
		.A2(I10[9]),
		.B1(out_sel[11]),
		.B2(I11[9]),
		.Z(O5[9])
	);
	AN_CELL inst_and_9(
		.A1(out_sel[12]),
		.A2(I12[9]),
		.Z(O6[9])
	);
	AO_CELL inst_0_10(
		.A1(out_sel[0]),
		.A2(I0[10]),
		.B1(out_sel[1]),
		.B2(I1[10]),
		.Z(O0[10])
	);
	AO_CELL inst_1_10(
		.A1(out_sel[2]),
		.A2(I2[10]),
		.B1(out_sel[3]),
		.B2(I3[10]),
		.Z(O1[10])
	);
	AO_CELL inst_2_10(
		.A1(out_sel[4]),
		.A2(I4[10]),
		.B1(out_sel[5]),
		.B2(I5[10]),
		.Z(O2[10])
	);
	AO_CELL inst_3_10(
		.A1(out_sel[6]),
		.A2(I6[10]),
		.B1(out_sel[7]),
		.B2(I7[10]),
		.Z(O3[10])
	);
	AO_CELL inst_4_10(
		.A1(out_sel[8]),
		.A2(I8[10]),
		.B1(out_sel[9]),
		.B2(I9[10]),
		.Z(O4[10])
	);
	AO_CELL inst_5_10(
		.A1(out_sel[10]),
		.A2(I10[10]),
		.B1(out_sel[11]),
		.B2(I11[10]),
		.Z(O5[10])
	);
	AN_CELL inst_and_10(
		.A1(out_sel[12]),
		.A2(I12[10]),
		.Z(O6[10])
	);
	AO_CELL inst_0_11(
		.A1(out_sel[0]),
		.A2(I0[11]),
		.B1(out_sel[1]),
		.B2(I1[11]),
		.Z(O0[11])
	);
	AO_CELL inst_1_11(
		.A1(out_sel[2]),
		.A2(I2[11]),
		.B1(out_sel[3]),
		.B2(I3[11]),
		.Z(O1[11])
	);
	AO_CELL inst_2_11(
		.A1(out_sel[4]),
		.A2(I4[11]),
		.B1(out_sel[5]),
		.B2(I5[11]),
		.Z(O2[11])
	);
	AO_CELL inst_3_11(
		.A1(out_sel[6]),
		.A2(I6[11]),
		.B1(out_sel[7]),
		.B2(I7[11]),
		.Z(O3[11])
	);
	AO_CELL inst_4_11(
		.A1(out_sel[8]),
		.A2(I8[11]),
		.B1(out_sel[9]),
		.B2(I9[11]),
		.Z(O4[11])
	);
	AO_CELL inst_5_11(
		.A1(out_sel[10]),
		.A2(I10[11]),
		.B1(out_sel[11]),
		.B2(I11[11]),
		.Z(O5[11])
	);
	AN_CELL inst_and_11(
		.A1(out_sel[12]),
		.A2(I12[11]),
		.Z(O6[11])
	);
	AO_CELL inst_0_12(
		.A1(out_sel[0]),
		.A2(I0[12]),
		.B1(out_sel[1]),
		.B2(I1[12]),
		.Z(O0[12])
	);
	AO_CELL inst_1_12(
		.A1(out_sel[2]),
		.A2(I2[12]),
		.B1(out_sel[3]),
		.B2(I3[12]),
		.Z(O1[12])
	);
	AO_CELL inst_2_12(
		.A1(out_sel[4]),
		.A2(I4[12]),
		.B1(out_sel[5]),
		.B2(I5[12]),
		.Z(O2[12])
	);
	AO_CELL inst_3_12(
		.A1(out_sel[6]),
		.A2(I6[12]),
		.B1(out_sel[7]),
		.B2(I7[12]),
		.Z(O3[12])
	);
	AO_CELL inst_4_12(
		.A1(out_sel[8]),
		.A2(I8[12]),
		.B1(out_sel[9]),
		.B2(I9[12]),
		.Z(O4[12])
	);
	AO_CELL inst_5_12(
		.A1(out_sel[10]),
		.A2(I10[12]),
		.B1(out_sel[11]),
		.B2(I11[12]),
		.Z(O5[12])
	);
	AN_CELL inst_and_12(
		.A1(out_sel[12]),
		.A2(I12[12]),
		.Z(O6[12])
	);
	AO_CELL inst_0_13(
		.A1(out_sel[0]),
		.A2(I0[13]),
		.B1(out_sel[1]),
		.B2(I1[13]),
		.Z(O0[13])
	);
	AO_CELL inst_1_13(
		.A1(out_sel[2]),
		.A2(I2[13]),
		.B1(out_sel[3]),
		.B2(I3[13]),
		.Z(O1[13])
	);
	AO_CELL inst_2_13(
		.A1(out_sel[4]),
		.A2(I4[13]),
		.B1(out_sel[5]),
		.B2(I5[13]),
		.Z(O2[13])
	);
	AO_CELL inst_3_13(
		.A1(out_sel[6]),
		.A2(I6[13]),
		.B1(out_sel[7]),
		.B2(I7[13]),
		.Z(O3[13])
	);
	AO_CELL inst_4_13(
		.A1(out_sel[8]),
		.A2(I8[13]),
		.B1(out_sel[9]),
		.B2(I9[13]),
		.Z(O4[13])
	);
	AO_CELL inst_5_13(
		.A1(out_sel[10]),
		.A2(I10[13]),
		.B1(out_sel[11]),
		.B2(I11[13]),
		.Z(O5[13])
	);
	AN_CELL inst_and_13(
		.A1(out_sel[12]),
		.A2(I12[13]),
		.Z(O6[13])
	);
	AO_CELL inst_0_14(
		.A1(out_sel[0]),
		.A2(I0[14]),
		.B1(out_sel[1]),
		.B2(I1[14]),
		.Z(O0[14])
	);
	AO_CELL inst_1_14(
		.A1(out_sel[2]),
		.A2(I2[14]),
		.B1(out_sel[3]),
		.B2(I3[14]),
		.Z(O1[14])
	);
	AO_CELL inst_2_14(
		.A1(out_sel[4]),
		.A2(I4[14]),
		.B1(out_sel[5]),
		.B2(I5[14]),
		.Z(O2[14])
	);
	AO_CELL inst_3_14(
		.A1(out_sel[6]),
		.A2(I6[14]),
		.B1(out_sel[7]),
		.B2(I7[14]),
		.Z(O3[14])
	);
	AO_CELL inst_4_14(
		.A1(out_sel[8]),
		.A2(I8[14]),
		.B1(out_sel[9]),
		.B2(I9[14]),
		.Z(O4[14])
	);
	AO_CELL inst_5_14(
		.A1(out_sel[10]),
		.A2(I10[14]),
		.B1(out_sel[11]),
		.B2(I11[14]),
		.Z(O5[14])
	);
	AN_CELL inst_and_14(
		.A1(out_sel[12]),
		.A2(I12[14]),
		.Z(O6[14])
	);
	AO_CELL inst_0_15(
		.A1(out_sel[0]),
		.A2(I0[15]),
		.B1(out_sel[1]),
		.B2(I1[15]),
		.Z(O0[15])
	);
	AO_CELL inst_1_15(
		.A1(out_sel[2]),
		.A2(I2[15]),
		.B1(out_sel[3]),
		.B2(I3[15]),
		.Z(O1[15])
	);
	AO_CELL inst_2_15(
		.A1(out_sel[4]),
		.A2(I4[15]),
		.B1(out_sel[5]),
		.B2(I5[15]),
		.Z(O2[15])
	);
	AO_CELL inst_3_15(
		.A1(out_sel[6]),
		.A2(I6[15]),
		.B1(out_sel[7]),
		.B2(I7[15]),
		.Z(O3[15])
	);
	AO_CELL inst_4_15(
		.A1(out_sel[8]),
		.A2(I8[15]),
		.B1(out_sel[9]),
		.B2(I9[15]),
		.Z(O4[15])
	);
	AO_CELL inst_5_15(
		.A1(out_sel[10]),
		.A2(I10[15]),
		.B1(out_sel[11]),
		.B2(I11[15]),
		.Z(O5[15])
	);
	AN_CELL inst_and_15(
		.A1(out_sel[12]),
		.A2(I12[15]),
		.Z(O6[15])
	);
	AO_CELL inst_0_16(
		.A1(out_sel[0]),
		.A2(I0[16]),
		.B1(out_sel[1]),
		.B2(I1[16]),
		.Z(O0[16])
	);
	AO_CELL inst_1_16(
		.A1(out_sel[2]),
		.A2(I2[16]),
		.B1(out_sel[3]),
		.B2(I3[16]),
		.Z(O1[16])
	);
	AO_CELL inst_2_16(
		.A1(out_sel[4]),
		.A2(I4[16]),
		.B1(out_sel[5]),
		.B2(I5[16]),
		.Z(O2[16])
	);
	AO_CELL inst_3_16(
		.A1(out_sel[6]),
		.A2(I6[16]),
		.B1(out_sel[7]),
		.B2(I7[16]),
		.Z(O3[16])
	);
	AO_CELL inst_4_16(
		.A1(out_sel[8]),
		.A2(I8[16]),
		.B1(out_sel[9]),
		.B2(I9[16]),
		.Z(O4[16])
	);
	AO_CELL inst_5_16(
		.A1(out_sel[10]),
		.A2(I10[16]),
		.B1(out_sel[11]),
		.B2(I11[16]),
		.Z(O5[16])
	);
	AN_CELL inst_and_16(
		.A1(out_sel[12]),
		.A2(I12[16]),
		.Z(O6[16])
	);
	AO_CELL inst_0_17(
		.A1(out_sel[0]),
		.A2(I0[17]),
		.B1(out_sel[1]),
		.B2(I1[17]),
		.Z(O0[17])
	);
	AO_CELL inst_1_17(
		.A1(out_sel[2]),
		.A2(I2[17]),
		.B1(out_sel[3]),
		.B2(I3[17]),
		.Z(O1[17])
	);
	AO_CELL inst_2_17(
		.A1(out_sel[4]),
		.A2(I4[17]),
		.B1(out_sel[5]),
		.B2(I5[17]),
		.Z(O2[17])
	);
	AO_CELL inst_3_17(
		.A1(out_sel[6]),
		.A2(I6[17]),
		.B1(out_sel[7]),
		.B2(I7[17]),
		.Z(O3[17])
	);
	AO_CELL inst_4_17(
		.A1(out_sel[8]),
		.A2(I8[17]),
		.B1(out_sel[9]),
		.B2(I9[17]),
		.Z(O4[17])
	);
	AO_CELL inst_5_17(
		.A1(out_sel[10]),
		.A2(I10[17]),
		.B1(out_sel[11]),
		.B2(I11[17]),
		.Z(O5[17])
	);
	AN_CELL inst_and_17(
		.A1(out_sel[12]),
		.A2(I12[17]),
		.Z(O6[17])
	);
	AO_CELL inst_0_18(
		.A1(out_sel[0]),
		.A2(I0[18]),
		.B1(out_sel[1]),
		.B2(I1[18]),
		.Z(O0[18])
	);
	AO_CELL inst_1_18(
		.A1(out_sel[2]),
		.A2(I2[18]),
		.B1(out_sel[3]),
		.B2(I3[18]),
		.Z(O1[18])
	);
	AO_CELL inst_2_18(
		.A1(out_sel[4]),
		.A2(I4[18]),
		.B1(out_sel[5]),
		.B2(I5[18]),
		.Z(O2[18])
	);
	AO_CELL inst_3_18(
		.A1(out_sel[6]),
		.A2(I6[18]),
		.B1(out_sel[7]),
		.B2(I7[18]),
		.Z(O3[18])
	);
	AO_CELL inst_4_18(
		.A1(out_sel[8]),
		.A2(I8[18]),
		.B1(out_sel[9]),
		.B2(I9[18]),
		.Z(O4[18])
	);
	AO_CELL inst_5_18(
		.A1(out_sel[10]),
		.A2(I10[18]),
		.B1(out_sel[11]),
		.B2(I11[18]),
		.Z(O5[18])
	);
	AN_CELL inst_and_18(
		.A1(out_sel[12]),
		.A2(I12[18]),
		.Z(O6[18])
	);
	AO_CELL inst_0_19(
		.A1(out_sel[0]),
		.A2(I0[19]),
		.B1(out_sel[1]),
		.B2(I1[19]),
		.Z(O0[19])
	);
	AO_CELL inst_1_19(
		.A1(out_sel[2]),
		.A2(I2[19]),
		.B1(out_sel[3]),
		.B2(I3[19]),
		.Z(O1[19])
	);
	AO_CELL inst_2_19(
		.A1(out_sel[4]),
		.A2(I4[19]),
		.B1(out_sel[5]),
		.B2(I5[19]),
		.Z(O2[19])
	);
	AO_CELL inst_3_19(
		.A1(out_sel[6]),
		.A2(I6[19]),
		.B1(out_sel[7]),
		.B2(I7[19]),
		.Z(O3[19])
	);
	AO_CELL inst_4_19(
		.A1(out_sel[8]),
		.A2(I8[19]),
		.B1(out_sel[9]),
		.B2(I9[19]),
		.Z(O4[19])
	);
	AO_CELL inst_5_19(
		.A1(out_sel[10]),
		.A2(I10[19]),
		.B1(out_sel[11]),
		.B2(I11[19]),
		.Z(O5[19])
	);
	AN_CELL inst_and_19(
		.A1(out_sel[12]),
		.A2(I12[19]),
		.Z(O6[19])
	);
	AO_CELL inst_0_20(
		.A1(out_sel[0]),
		.A2(I0[20]),
		.B1(out_sel[1]),
		.B2(I1[20]),
		.Z(O0[20])
	);
	AO_CELL inst_1_20(
		.A1(out_sel[2]),
		.A2(I2[20]),
		.B1(out_sel[3]),
		.B2(I3[20]),
		.Z(O1[20])
	);
	AO_CELL inst_2_20(
		.A1(out_sel[4]),
		.A2(I4[20]),
		.B1(out_sel[5]),
		.B2(I5[20]),
		.Z(O2[20])
	);
	AO_CELL inst_3_20(
		.A1(out_sel[6]),
		.A2(I6[20]),
		.B1(out_sel[7]),
		.B2(I7[20]),
		.Z(O3[20])
	);
	AO_CELL inst_4_20(
		.A1(out_sel[8]),
		.A2(I8[20]),
		.B1(out_sel[9]),
		.B2(I9[20]),
		.Z(O4[20])
	);
	AO_CELL inst_5_20(
		.A1(out_sel[10]),
		.A2(I10[20]),
		.B1(out_sel[11]),
		.B2(I11[20]),
		.Z(O5[20])
	);
	AN_CELL inst_and_20(
		.A1(out_sel[12]),
		.A2(I12[20]),
		.Z(O6[20])
	);
	AO_CELL inst_0_21(
		.A1(out_sel[0]),
		.A2(I0[21]),
		.B1(out_sel[1]),
		.B2(I1[21]),
		.Z(O0[21])
	);
	AO_CELL inst_1_21(
		.A1(out_sel[2]),
		.A2(I2[21]),
		.B1(out_sel[3]),
		.B2(I3[21]),
		.Z(O1[21])
	);
	AO_CELL inst_2_21(
		.A1(out_sel[4]),
		.A2(I4[21]),
		.B1(out_sel[5]),
		.B2(I5[21]),
		.Z(O2[21])
	);
	AO_CELL inst_3_21(
		.A1(out_sel[6]),
		.A2(I6[21]),
		.B1(out_sel[7]),
		.B2(I7[21]),
		.Z(O3[21])
	);
	AO_CELL inst_4_21(
		.A1(out_sel[8]),
		.A2(I8[21]),
		.B1(out_sel[9]),
		.B2(I9[21]),
		.Z(O4[21])
	);
	AO_CELL inst_5_21(
		.A1(out_sel[10]),
		.A2(I10[21]),
		.B1(out_sel[11]),
		.B2(I11[21]),
		.Z(O5[21])
	);
	AN_CELL inst_and_21(
		.A1(out_sel[12]),
		.A2(I12[21]),
		.Z(O6[21])
	);
	AO_CELL inst_0_22(
		.A1(out_sel[0]),
		.A2(I0[22]),
		.B1(out_sel[1]),
		.B2(I1[22]),
		.Z(O0[22])
	);
	AO_CELL inst_1_22(
		.A1(out_sel[2]),
		.A2(I2[22]),
		.B1(out_sel[3]),
		.B2(I3[22]),
		.Z(O1[22])
	);
	AO_CELL inst_2_22(
		.A1(out_sel[4]),
		.A2(I4[22]),
		.B1(out_sel[5]),
		.B2(I5[22]),
		.Z(O2[22])
	);
	AO_CELL inst_3_22(
		.A1(out_sel[6]),
		.A2(I6[22]),
		.B1(out_sel[7]),
		.B2(I7[22]),
		.Z(O3[22])
	);
	AO_CELL inst_4_22(
		.A1(out_sel[8]),
		.A2(I8[22]),
		.B1(out_sel[9]),
		.B2(I9[22]),
		.Z(O4[22])
	);
	AO_CELL inst_5_22(
		.A1(out_sel[10]),
		.A2(I10[22]),
		.B1(out_sel[11]),
		.B2(I11[22]),
		.Z(O5[22])
	);
	AN_CELL inst_and_22(
		.A1(out_sel[12]),
		.A2(I12[22]),
		.Z(O6[22])
	);
	AO_CELL inst_0_23(
		.A1(out_sel[0]),
		.A2(I0[23]),
		.B1(out_sel[1]),
		.B2(I1[23]),
		.Z(O0[23])
	);
	AO_CELL inst_1_23(
		.A1(out_sel[2]),
		.A2(I2[23]),
		.B1(out_sel[3]),
		.B2(I3[23]),
		.Z(O1[23])
	);
	AO_CELL inst_2_23(
		.A1(out_sel[4]),
		.A2(I4[23]),
		.B1(out_sel[5]),
		.B2(I5[23]),
		.Z(O2[23])
	);
	AO_CELL inst_3_23(
		.A1(out_sel[6]),
		.A2(I6[23]),
		.B1(out_sel[7]),
		.B2(I7[23]),
		.Z(O3[23])
	);
	AO_CELL inst_4_23(
		.A1(out_sel[8]),
		.A2(I8[23]),
		.B1(out_sel[9]),
		.B2(I9[23]),
		.Z(O4[23])
	);
	AO_CELL inst_5_23(
		.A1(out_sel[10]),
		.A2(I10[23]),
		.B1(out_sel[11]),
		.B2(I11[23]),
		.Z(O5[23])
	);
	AN_CELL inst_and_23(
		.A1(out_sel[12]),
		.A2(I12[23]),
		.Z(O6[23])
	);
	AO_CELL inst_0_24(
		.A1(out_sel[0]),
		.A2(I0[24]),
		.B1(out_sel[1]),
		.B2(I1[24]),
		.Z(O0[24])
	);
	AO_CELL inst_1_24(
		.A1(out_sel[2]),
		.A2(I2[24]),
		.B1(out_sel[3]),
		.B2(I3[24]),
		.Z(O1[24])
	);
	AO_CELL inst_2_24(
		.A1(out_sel[4]),
		.A2(I4[24]),
		.B1(out_sel[5]),
		.B2(I5[24]),
		.Z(O2[24])
	);
	AO_CELL inst_3_24(
		.A1(out_sel[6]),
		.A2(I6[24]),
		.B1(out_sel[7]),
		.B2(I7[24]),
		.Z(O3[24])
	);
	AO_CELL inst_4_24(
		.A1(out_sel[8]),
		.A2(I8[24]),
		.B1(out_sel[9]),
		.B2(I9[24]),
		.Z(O4[24])
	);
	AO_CELL inst_5_24(
		.A1(out_sel[10]),
		.A2(I10[24]),
		.B1(out_sel[11]),
		.B2(I11[24]),
		.Z(O5[24])
	);
	AN_CELL inst_and_24(
		.A1(out_sel[12]),
		.A2(I12[24]),
		.Z(O6[24])
	);
	AO_CELL inst_0_25(
		.A1(out_sel[0]),
		.A2(I0[25]),
		.B1(out_sel[1]),
		.B2(I1[25]),
		.Z(O0[25])
	);
	AO_CELL inst_1_25(
		.A1(out_sel[2]),
		.A2(I2[25]),
		.B1(out_sel[3]),
		.B2(I3[25]),
		.Z(O1[25])
	);
	AO_CELL inst_2_25(
		.A1(out_sel[4]),
		.A2(I4[25]),
		.B1(out_sel[5]),
		.B2(I5[25]),
		.Z(O2[25])
	);
	AO_CELL inst_3_25(
		.A1(out_sel[6]),
		.A2(I6[25]),
		.B1(out_sel[7]),
		.B2(I7[25]),
		.Z(O3[25])
	);
	AO_CELL inst_4_25(
		.A1(out_sel[8]),
		.A2(I8[25]),
		.B1(out_sel[9]),
		.B2(I9[25]),
		.Z(O4[25])
	);
	AO_CELL inst_5_25(
		.A1(out_sel[10]),
		.A2(I10[25]),
		.B1(out_sel[11]),
		.B2(I11[25]),
		.Z(O5[25])
	);
	AN_CELL inst_and_25(
		.A1(out_sel[12]),
		.A2(I12[25]),
		.Z(O6[25])
	);
	AO_CELL inst_0_26(
		.A1(out_sel[0]),
		.A2(I0[26]),
		.B1(out_sel[1]),
		.B2(I1[26]),
		.Z(O0[26])
	);
	AO_CELL inst_1_26(
		.A1(out_sel[2]),
		.A2(I2[26]),
		.B1(out_sel[3]),
		.B2(I3[26]),
		.Z(O1[26])
	);
	AO_CELL inst_2_26(
		.A1(out_sel[4]),
		.A2(I4[26]),
		.B1(out_sel[5]),
		.B2(I5[26]),
		.Z(O2[26])
	);
	AO_CELL inst_3_26(
		.A1(out_sel[6]),
		.A2(I6[26]),
		.B1(out_sel[7]),
		.B2(I7[26]),
		.Z(O3[26])
	);
	AO_CELL inst_4_26(
		.A1(out_sel[8]),
		.A2(I8[26]),
		.B1(out_sel[9]),
		.B2(I9[26]),
		.Z(O4[26])
	);
	AO_CELL inst_5_26(
		.A1(out_sel[10]),
		.A2(I10[26]),
		.B1(out_sel[11]),
		.B2(I11[26]),
		.Z(O5[26])
	);
	AN_CELL inst_and_26(
		.A1(out_sel[12]),
		.A2(I12[26]),
		.Z(O6[26])
	);
	AO_CELL inst_0_27(
		.A1(out_sel[0]),
		.A2(I0[27]),
		.B1(out_sel[1]),
		.B2(I1[27]),
		.Z(O0[27])
	);
	AO_CELL inst_1_27(
		.A1(out_sel[2]),
		.A2(I2[27]),
		.B1(out_sel[3]),
		.B2(I3[27]),
		.Z(O1[27])
	);
	AO_CELL inst_2_27(
		.A1(out_sel[4]),
		.A2(I4[27]),
		.B1(out_sel[5]),
		.B2(I5[27]),
		.Z(O2[27])
	);
	AO_CELL inst_3_27(
		.A1(out_sel[6]),
		.A2(I6[27]),
		.B1(out_sel[7]),
		.B2(I7[27]),
		.Z(O3[27])
	);
	AO_CELL inst_4_27(
		.A1(out_sel[8]),
		.A2(I8[27]),
		.B1(out_sel[9]),
		.B2(I9[27]),
		.Z(O4[27])
	);
	AO_CELL inst_5_27(
		.A1(out_sel[10]),
		.A2(I10[27]),
		.B1(out_sel[11]),
		.B2(I11[27]),
		.Z(O5[27])
	);
	AN_CELL inst_and_27(
		.A1(out_sel[12]),
		.A2(I12[27]),
		.Z(O6[27])
	);
	AO_CELL inst_0_28(
		.A1(out_sel[0]),
		.A2(I0[28]),
		.B1(out_sel[1]),
		.B2(I1[28]),
		.Z(O0[28])
	);
	AO_CELL inst_1_28(
		.A1(out_sel[2]),
		.A2(I2[28]),
		.B1(out_sel[3]),
		.B2(I3[28]),
		.Z(O1[28])
	);
	AO_CELL inst_2_28(
		.A1(out_sel[4]),
		.A2(I4[28]),
		.B1(out_sel[5]),
		.B2(I5[28]),
		.Z(O2[28])
	);
	AO_CELL inst_3_28(
		.A1(out_sel[6]),
		.A2(I6[28]),
		.B1(out_sel[7]),
		.B2(I7[28]),
		.Z(O3[28])
	);
	AO_CELL inst_4_28(
		.A1(out_sel[8]),
		.A2(I8[28]),
		.B1(out_sel[9]),
		.B2(I9[28]),
		.Z(O4[28])
	);
	AO_CELL inst_5_28(
		.A1(out_sel[10]),
		.A2(I10[28]),
		.B1(out_sel[11]),
		.B2(I11[28]),
		.Z(O5[28])
	);
	AN_CELL inst_and_28(
		.A1(out_sel[12]),
		.A2(I12[28]),
		.Z(O6[28])
	);
	AO_CELL inst_0_29(
		.A1(out_sel[0]),
		.A2(I0[29]),
		.B1(out_sel[1]),
		.B2(I1[29]),
		.Z(O0[29])
	);
	AO_CELL inst_1_29(
		.A1(out_sel[2]),
		.A2(I2[29]),
		.B1(out_sel[3]),
		.B2(I3[29]),
		.Z(O1[29])
	);
	AO_CELL inst_2_29(
		.A1(out_sel[4]),
		.A2(I4[29]),
		.B1(out_sel[5]),
		.B2(I5[29]),
		.Z(O2[29])
	);
	AO_CELL inst_3_29(
		.A1(out_sel[6]),
		.A2(I6[29]),
		.B1(out_sel[7]),
		.B2(I7[29]),
		.Z(O3[29])
	);
	AO_CELL inst_4_29(
		.A1(out_sel[8]),
		.A2(I8[29]),
		.B1(out_sel[9]),
		.B2(I9[29]),
		.Z(O4[29])
	);
	AO_CELL inst_5_29(
		.A1(out_sel[10]),
		.A2(I10[29]),
		.B1(out_sel[11]),
		.B2(I11[29]),
		.Z(O5[29])
	);
	AN_CELL inst_and_29(
		.A1(out_sel[12]),
		.A2(I12[29]),
		.Z(O6[29])
	);
	AO_CELL inst_0_30(
		.A1(out_sel[0]),
		.A2(I0[30]),
		.B1(out_sel[1]),
		.B2(I1[30]),
		.Z(O0[30])
	);
	AO_CELL inst_1_30(
		.A1(out_sel[2]),
		.A2(I2[30]),
		.B1(out_sel[3]),
		.B2(I3[30]),
		.Z(O1[30])
	);
	AO_CELL inst_2_30(
		.A1(out_sel[4]),
		.A2(I4[30]),
		.B1(out_sel[5]),
		.B2(I5[30]),
		.Z(O2[30])
	);
	AO_CELL inst_3_30(
		.A1(out_sel[6]),
		.A2(I6[30]),
		.B1(out_sel[7]),
		.B2(I7[30]),
		.Z(O3[30])
	);
	AO_CELL inst_4_30(
		.A1(out_sel[8]),
		.A2(I8[30]),
		.B1(out_sel[9]),
		.B2(I9[30]),
		.Z(O4[30])
	);
	AO_CELL inst_5_30(
		.A1(out_sel[10]),
		.A2(I10[30]),
		.B1(out_sel[11]),
		.B2(I11[30]),
		.Z(O5[30])
	);
	AN_CELL inst_and_30(
		.A1(out_sel[12]),
		.A2(I12[30]),
		.Z(O6[30])
	);
	AO_CELL inst_0_31(
		.A1(out_sel[0]),
		.A2(I0[31]),
		.B1(out_sel[1]),
		.B2(I1[31]),
		.Z(O0[31])
	);
	AO_CELL inst_1_31(
		.A1(out_sel[2]),
		.A2(I2[31]),
		.B1(out_sel[3]),
		.B2(I3[31]),
		.Z(O1[31])
	);
	AO_CELL inst_2_31(
		.A1(out_sel[4]),
		.A2(I4[31]),
		.B1(out_sel[5]),
		.B2(I5[31]),
		.Z(O2[31])
	);
	AO_CELL inst_3_31(
		.A1(out_sel[6]),
		.A2(I6[31]),
		.B1(out_sel[7]),
		.B2(I7[31]),
		.Z(O3[31])
	);
	AO_CELL inst_4_31(
		.A1(out_sel[8]),
		.A2(I8[31]),
		.B1(out_sel[9]),
		.B2(I9[31]),
		.Z(O4[31])
	);
	AO_CELL inst_5_31(
		.A1(out_sel[10]),
		.A2(I10[31]),
		.B1(out_sel[11]),
		.B2(I11[31]),
		.Z(O5[31])
	);
	AN_CELL inst_and_31(
		.A1(out_sel[12]),
		.A2(I12[31]),
		.Z(O6[31])
	);
endmodule
module mantle_wire__typeBitIn32 (
	in,
	out
);
	output wire [31:0] in;
	input [31:0] out;
	assign in = out;
endmodule
module mantle_wire__typeBitIn17 (
	in,
	out
);
	output wire [16:0] in;
	input [16:0] out;
	assign in = out;
endmodule
module mantle_wire__typeBit8 (
	in,
	out
);
	input [7:0] in;
	output wire [7:0] out;
	assign out = in;
endmodule
module mantle_wire__typeBit4 (
	in,
	out
);
	input [3:0] in;
	output wire [3:0] out;
	assign out = in;
endmodule
module mantle_wire__typeBit32 (
	in,
	out
);
	input [31:0] in;
	output wire [31:0] out;
	assign out = in;
endmodule
module mantle_wire__typeBit17 (
	in,
	out
);
	input [16:0] in;
	output wire [16:0] out;
	assign out = in;
endmodule
module regCE_arst (
	in,
	ce,
	out,
	clk,
	arst
);
	parameter width = 1;
	parameter init = 1;
	input [width - 1:0] in;
	input ce;
	output wire [width - 1:0] out;
	input clk;
	input arst;
	reg [width - 1:0] value;
	always @(posedge clk or posedge arst)
		if (arst)
			value <= init;
		else if (ce)
			value <= in;
	assign out = value;
endmodule
module io_core (
	clk,
	clk_en,
	f2io_1,
	f2io_17,
	f2io_17_valid,
	f2io_1_valid,
	flush,
	glb2io_1,
	glb2io_17,
	glb2io_17_valid,
	glb2io_1_valid,
	io2f_17_ready,
	io2f_1_ready,
	io2glb_17_ready,
	io2glb_1_ready,
	rst_n,
	tile_en,
	f2io_17_ready,
	f2io_1_ready,
	glb2io_17_ready,
	glb2io_1_ready,
	io2f_1,
	io2f_17,
	io2f_17_valid,
	io2f_1_valid,
	io2glb_1,
	io2glb_17,
	io2glb_17_valid,
	io2glb_1_valid
);
	input wire clk;
	input wire clk_en;
	input wire f2io_1;
	input wire [16:0] f2io_17;
	input wire f2io_17_valid;
	input wire f2io_1_valid;
	input wire flush;
	input wire glb2io_1;
	input wire [16:0] glb2io_17;
	input wire glb2io_17_valid;
	input wire glb2io_1_valid;
	input wire io2f_17_ready;
	input wire io2f_1_ready;
	input wire io2glb_17_ready;
	input wire io2glb_1_ready;
	input wire rst_n;
	input wire tile_en;
	output wire f2io_17_ready;
	output wire f2io_1_ready;
	output wire glb2io_17_ready;
	output wire glb2io_1_ready;
	output wire io2f_1;
	output wire [16:0] io2f_17;
	output wire io2f_17_valid;
	output wire io2f_1_valid;
	output wire io2glb_1;
	output wire [16:0] io2glb_17;
	output wire io2glb_17_valid;
	output wire io2glb_1_valid;
	wire [16:0] f2io_2_io2glb_17_data_out;
	wire f2io_2_io2glb_17_empty;
	wire f2io_2_io2glb_17_full;
	wire [0:0] f2io_2_io2glb_1_data_out;
	wire f2io_2_io2glb_1_empty;
	wire f2io_2_io2glb_1_full;
	wire gclk;
	wire glb2io_2_io2f_17_empty;
	wire glb2io_2_io2f_17_full;
	wire glb2io_2_io2f_1_empty;
	wire glb2io_2_io2f_1_full;
	assign gclk = clk & tile_en;
	assign io2glb_1 = f2io_2_io2glb_1_data_out;
	assign f2io_1_ready = ~f2io_2_io2glb_1_full;
	assign io2glb_1_valid = ~f2io_2_io2glb_1_empty;
	assign glb2io_1_ready = ~glb2io_2_io2f_1_full;
	assign io2f_1_valid = ~glb2io_2_io2f_1_empty;
	assign io2glb_17 = f2io_2_io2glb_17_data_out[16-:17];
	assign f2io_17_ready = ~f2io_2_io2glb_17_full;
	assign io2glb_17_valid = ~f2io_2_io2glb_17_empty;
	assign glb2io_17_ready = ~glb2io_2_io2f_17_full;
	assign io2f_17_valid = ~glb2io_2_io2f_17_empty;
	reg_fifo_depth_2_w_1_afd_1_iocore_nof f2io_2_io2glb_1(
		.clk(clk),
		.clk_en(clk_en),
		.data_in(f2io_1),
		.flush(flush),
		.pop(io2glb_1_ready),
		.push(f2io_1_valid),
		.rst_n(rst_n),
		.data_out(f2io_2_io2glb_1_data_out),
		.empty(f2io_2_io2glb_1_empty),
		.full(f2io_2_io2glb_1_full)
	);
	reg_fifo_depth_2_w_1_afd_1_iocore_nof glb2io_2_io2f_1(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(glb2io_1),
		.flush(flush),
		.pop(io2f_1_ready),
		.push(glb2io_1_valid),
		.rst_n(rst_n),
		.data_out(io2f_1),
		.empty(glb2io_2_io2f_1_empty),
		.full(glb2io_2_io2f_1_full)
	);
	reg_fifo_depth_2_w_17_afd_1_iocore_nof f2io_2_io2glb_17(
		.clk(clk),
		.clk_en(clk_en),
		.data_in(f2io_17),
		.flush(flush),
		.pop(io2glb_17_ready),
		.push(f2io_17_valid),
		.rst_n(rst_n),
		.data_out(f2io_2_io2glb_17_data_out),
		.empty(f2io_2_io2glb_17_empty),
		.full(f2io_2_io2glb_17_full)
	);
	reg_fifo_depth_2_w_17_afd_1_iocore_nof glb2io_2_io2f_17(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(glb2io_17),
		.flush(flush),
		.pop(io2f_17_ready),
		.push(glb2io_17_valid),
		.rst_n(rst_n),
		.data_out(io2f_17),
		.empty(glb2io_2_io2f_17_empty),
		.full(glb2io_2_io2f_17_full)
	);
endmodule
module io_core_W (
	clk,
	clk_en,
	f2io_1,
	f2io_17,
	f2io_17_valid,
	f2io_1_valid,
	flush,
	glb2io_1,
	glb2io_17,
	glb2io_17_valid,
	glb2io_1_valid,
	io2f_17_ready,
	io2f_1_ready,
	io2glb_17_ready,
	io2glb_1_ready,
	rst_n,
	tile_en,
	f2io_17_ready,
	f2io_1_ready,
	glb2io_17_ready,
	glb2io_1_ready,
	io2f_1,
	io2f_17,
	io2f_17_valid,
	io2f_1_valid,
	io2glb_1,
	io2glb_17,
	io2glb_17_valid,
	io2glb_1_valid
);
	input wire clk;
	input wire clk_en;
	input wire f2io_1;
	input wire [16:0] f2io_17;
	input wire f2io_17_valid;
	input wire f2io_1_valid;
	input wire flush;
	input wire glb2io_1;
	input wire [16:0] glb2io_17;
	input wire glb2io_17_valid;
	input wire glb2io_1_valid;
	input wire io2f_17_ready;
	input wire io2f_1_ready;
	input wire io2glb_17_ready;
	input wire io2glb_1_ready;
	input wire rst_n;
	input wire tile_en;
	output wire f2io_17_ready;
	output wire f2io_1_ready;
	output wire glb2io_17_ready;
	output wire glb2io_1_ready;
	output wire io2f_1;
	output wire [16:0] io2f_17;
	output wire io2f_17_valid;
	output wire io2f_1_valid;
	output wire io2glb_1;
	output wire [16:0] io2glb_17;
	output wire io2glb_17_valid;
	output wire io2glb_1_valid;
	io_core io_core(
		.clk(clk),
		.clk_en(clk_en),
		.f2io_1(f2io_1),
		.f2io_17(f2io_17),
		.f2io_17_valid(f2io_17_valid),
		.f2io_1_valid(f2io_1_valid),
		.flush(flush),
		.glb2io_1(glb2io_1),
		.glb2io_17(glb2io_17),
		.glb2io_17_valid(glb2io_17_valid),
		.glb2io_1_valid(glb2io_1_valid),
		.io2f_17_ready(io2f_17_ready),
		.io2f_1_ready(io2f_1_ready),
		.io2glb_17_ready(io2glb_17_ready),
		.io2glb_1_ready(io2glb_1_ready),
		.rst_n(rst_n),
		.tile_en(tile_en),
		.f2io_17_ready(f2io_17_ready),
		.f2io_1_ready(f2io_1_ready),
		.glb2io_17_ready(glb2io_17_ready),
		.glb2io_1_ready(glb2io_1_ready),
		.io2f_1(io2f_1),
		.io2f_17(io2f_17),
		.io2f_17_valid(io2f_17_valid),
		.io2f_1_valid(io2f_1_valid),
		.io2glb_1(io2glb_1),
		.io2glb_17(io2glb_17),
		.io2glb_17_valid(io2glb_17_valid),
		.io2glb_1_valid(io2glb_1_valid)
	);
endmodule
module reg_fifo_depth_2_w_17_afd_1_iocore_nof (
	clk,
	clk_en,
	data_in,
	flush,
	pop,
	push,
	rst_n,
	almost_full,
	data_out,
	empty,
	full,
	valid
);
	input wire clk;
	input wire clk_en;
	input wire [16:0] data_in;
	input wire flush;
	input wire pop;
	input wire push;
	input wire rst_n;
	output wire almost_full;
	output reg [16:0] data_out;
	output wire empty;
	output wire full;
	output reg valid;
	reg [1:0] num_items;
	wire passthru;
	reg rd_ptr;
	wire read;
	reg [33:0] reg_array;
	reg wr_ptr;
	wire write;
	assign full = num_items == 2'h2;
	assign almost_full = num_items >= 2'h1;
	assign empty = num_items == 2'h0;
	assign read = (pop & ~passthru) & ~empty;
	assign passthru = 1'h0;
	assign write = (push & ~passthru) & ~full;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			num_items <= 2'h0;
		else if (flush)
			num_items <= 2'h0;
		else if (clk_en) begin
			if (write & ~read)
				num_items <= num_items + 2'h1;
			else if (~write & read)
				num_items <= num_items - 2'h1;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			reg_array <= 34'h000000000;
		else if (flush)
			reg_array <= 34'h000000000;
		else if (clk_en) begin
			if (write)
				reg_array[17 * wr_ptr+:17] <= data_in;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			wr_ptr <= 1'h0;
		else if (flush)
			wr_ptr <= 1'h0;
		else if (clk_en) begin
			if (write) begin
				if (wr_ptr == 1'h1)
					wr_ptr <= 1'h0;
				else
					wr_ptr <= wr_ptr + 1'h1;
			end
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			rd_ptr <= 1'h0;
		else if (flush)
			rd_ptr <= 1'h0;
		else if (clk_en) begin
			if (read)
				rd_ptr <= rd_ptr + 1'h1;
		end
	always @(*)
		if (passthru)
			data_out = data_in;
		else
			data_out = reg_array[17 * rd_ptr+:17];
	always @(*) valid = ~empty | passthru;
endmodule
module reg_fifo_depth_2_w_1_afd_1_iocore_nof (
	clk,
	clk_en,
	data_in,
	flush,
	pop,
	push,
	rst_n,
	almost_full,
	data_out,
	empty,
	full,
	valid
);
	input wire clk;
	input wire clk_en;
	input wire [0:0] data_in;
	input wire flush;
	input wire pop;
	input wire push;
	input wire rst_n;
	output wire almost_full;
	output reg [0:0] data_out;
	output wire empty;
	output wire full;
	output reg valid;
	reg [1:0] num_items;
	wire passthru;
	reg rd_ptr;
	wire read;
	reg [1:0] reg_array;
	reg wr_ptr;
	wire write;
	assign full = num_items == 2'h2;
	assign almost_full = num_items >= 2'h1;
	assign empty = num_items == 2'h0;
	assign read = (pop & ~passthru) & ~empty;
	assign passthru = 1'h0;
	assign write = (push & ~passthru) & ~full;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			num_items <= 2'h0;
		else if (flush)
			num_items <= 2'h0;
		else if (clk_en) begin
			if (write & ~read)
				num_items <= num_items + 2'h1;
			else if (~write & read)
				num_items <= num_items - 2'h1;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			reg_array <= 2'h0;
		else if (flush)
			reg_array <= 2'h0;
		else if (clk_en) begin
			if (write)
				reg_array[wr_ptr+:1] <= data_in;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			wr_ptr <= 1'h0;
		else if (flush)
			wr_ptr <= 1'h0;
		else if (clk_en) begin
			if (write) begin
				if (wr_ptr == 1'h1)
					wr_ptr <= 1'h0;
				else
					wr_ptr <= wr_ptr + 1'h1;
			end
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			rd_ptr <= 1'h0;
		else if (flush)
			rd_ptr <= 1'h0;
		else if (clk_en) begin
			if (read)
				rd_ptr <= rd_ptr + 1'h1;
		end
	always @(*)
		if (passthru)
			data_out = data_in;
		else
			data_out = reg_array[rd_ptr+:1];
	always @(*) valid = ~empty | passthru;
endmodule
module IN12LP_S1DB_W04096B064M08S2_HB (
	A,
	BW,
	CEN,
	CLK,
	D,
	MA_SAWL0,
	MA_SAWL1,
	MA_STABAS0,
	MA_STABAS1,
	MA_VD0,
	MA_VD1,
	MA_WL0,
	MA_WL1,
	MA_WRAS0,
	MA_WRAS1,
	MA_WRT,
	RDWEN,
	T_LOGIC,
	T_Q_RST,
	Q
);
	input wire [11:0] A;
	input wire [63:0] BW;
	input wire CEN;
	input wire CLK;
	input wire [63:0] D;
	input wire MA_SAWL0;
	input wire MA_SAWL1;
	input wire MA_STABAS0;
	input wire MA_STABAS1;
	input wire MA_VD0;
	input wire MA_VD1;
	input wire MA_WL0;
	input wire MA_WL1;
	input wire MA_WRAS0;
	input wire MA_WRAS1;
	input wire MA_WRT;
	input wire RDWEN;
	input wire T_LOGIC;
	input wire T_Q_RST;
	output reg [63:0] Q;
	reg [63:0] data_array [4095:0];
	function automatic [5:0] sv2v_cast_6;
		input reg [5:0] inp;
		sv2v_cast_6 = inp;
	endfunction
	always @(posedge CLK)
		if (CEN == 1'h0) begin
			Q <= data_array[A];
			if (RDWEN == 1'h0) begin : sv2v_autoblock_1
				reg [31:0] i;
				for (i = 0; i < 64; i = i + 1)
					if (BW[sv2v_cast_6(i)])
						data_array[A][sv2v_cast_6(i)] <= D[sv2v_cast_6(i)];
			end
		end
endmodule
module SC7P5T_CKGPRELATNX1_SSC14R (
	CLK,
	E,
	TE,
	Z
);
	input wire CLK;
	input wire E;
	input wire TE;
	output wire Z;
	reg enable_latch;
	always @(*)
		if (~CLK)
			enable_latch = E;
	assign Z = CLK & enable_latch;
endmodule
module clk_gate (
	clk,
	enable,
	gclk
);
	input wire clk;
	input wire enable;
	output wire gclk;
	SC7P5T_CKGPRELATNX1_SSC14R CG_CELL(
		.CLK(clk),
		.E(enable),
		.TE(1'h0),
		.Z(gclk)
	);
endmodule
module glb_addr_gen_7 (
	clk,
	clk_en,
	mux_sel,
	reset,
	restart,
	start_addr,
	step,
	strides,
	addr_out
);
	parameter addr_width = 32'h00000010;
	parameter loop_level = 32'h00000007;
	input wire clk;
	input wire clk_en;
	input wire [2:0] mux_sel;
	input wire reset;
	input wire restart;
	input wire [addr_width - 1:0] start_addr;
	input wire step;
	input wire [(loop_level * addr_width) - 1:0] strides;
	output wire [addr_width - 1:0] addr_out;
	reg [addr_width - 1:0] current_addr;
	assign addr_out = start_addr + current_addr;
	always @(posedge clk or posedge reset)
		if (reset)
			current_addr <= 16'h0000;
		else if (clk_en) begin
			if (restart)
				current_addr <= 16'h0000;
			else if (step)
				current_addr <= current_addr + strides[mux_sel * addr_width+:addr_width];
		end
endmodule
module glb_addr_gen_8 (
	clk,
	clk_en,
	mux_sel,
	reset,
	restart,
	start_addr,
	step,
	strides,
	addr_out
);
	parameter addr_width = 32'h00000010;
	parameter loop_level = 32'h00000008;
	input wire clk;
	input wire clk_en;
	input wire [2:0] mux_sel;
	input wire reset;
	input wire restart;
	input wire [addr_width - 1:0] start_addr;
	input wire step;
	input wire [(loop_level * addr_width) - 1:0] strides;
	output wire [addr_width - 1:0] addr_out;
	reg [addr_width - 1:0] current_addr;
	assign addr_out = start_addr + current_addr;
	always @(posedge clk or posedge reset)
		if (reset)
			current_addr <= 16'h0000;
		else if (clk_en) begin
			if (restart)
				current_addr <= 16'h0000;
			else if (step)
				current_addr <= current_addr + strides[mux_sel * addr_width+:addr_width];
		end
endmodule
module glb_bank (
	clk,
	rdrq_packet,
	reset,
	wr_packet,
	rdrs_packet
);
	input wire clk;
	input wire [17:0] rdrq_packet;
	input wire reset;
	input wire [89:0] wr_packet;
	output reg [64:0] rdrs_packet;
	reg [16:0] mem_addr;
	reg [63:0] mem_data_in;
	reg [63:0] mem_data_in_bit_sel;
	wire [63:0] mem_data_out;
	reg mem_rd_en;
	reg mem_wr_en;
	reg [63:0] packet_rd_data_r;
	wire packet_rd_en_d;
	wire [63:0] wr_data_bit_sel;
	assign wr_data_bit_sel[0] = wr_packet[81];
	assign wr_data_bit_sel[1] = wr_packet[81];
	assign wr_data_bit_sel[2] = wr_packet[81];
	assign wr_data_bit_sel[3] = wr_packet[81];
	assign wr_data_bit_sel[4] = wr_packet[81];
	assign wr_data_bit_sel[5] = wr_packet[81];
	assign wr_data_bit_sel[6] = wr_packet[81];
	assign wr_data_bit_sel[7] = wr_packet[81];
	assign wr_data_bit_sel[8] = wr_packet[82];
	assign wr_data_bit_sel[9] = wr_packet[82];
	assign wr_data_bit_sel[10] = wr_packet[82];
	assign wr_data_bit_sel[11] = wr_packet[82];
	assign wr_data_bit_sel[12] = wr_packet[82];
	assign wr_data_bit_sel[13] = wr_packet[82];
	assign wr_data_bit_sel[14] = wr_packet[82];
	assign wr_data_bit_sel[15] = wr_packet[82];
	assign wr_data_bit_sel[16] = wr_packet[83];
	assign wr_data_bit_sel[17] = wr_packet[83];
	assign wr_data_bit_sel[18] = wr_packet[83];
	assign wr_data_bit_sel[19] = wr_packet[83];
	assign wr_data_bit_sel[20] = wr_packet[83];
	assign wr_data_bit_sel[21] = wr_packet[83];
	assign wr_data_bit_sel[22] = wr_packet[83];
	assign wr_data_bit_sel[23] = wr_packet[83];
	assign wr_data_bit_sel[24] = wr_packet[84];
	assign wr_data_bit_sel[25] = wr_packet[84];
	assign wr_data_bit_sel[26] = wr_packet[84];
	assign wr_data_bit_sel[27] = wr_packet[84];
	assign wr_data_bit_sel[28] = wr_packet[84];
	assign wr_data_bit_sel[29] = wr_packet[84];
	assign wr_data_bit_sel[30] = wr_packet[84];
	assign wr_data_bit_sel[31] = wr_packet[84];
	assign wr_data_bit_sel[32] = wr_packet[85];
	assign wr_data_bit_sel[33] = wr_packet[85];
	assign wr_data_bit_sel[34] = wr_packet[85];
	assign wr_data_bit_sel[35] = wr_packet[85];
	assign wr_data_bit_sel[36] = wr_packet[85];
	assign wr_data_bit_sel[37] = wr_packet[85];
	assign wr_data_bit_sel[38] = wr_packet[85];
	assign wr_data_bit_sel[39] = wr_packet[85];
	assign wr_data_bit_sel[40] = wr_packet[86];
	assign wr_data_bit_sel[41] = wr_packet[86];
	assign wr_data_bit_sel[42] = wr_packet[86];
	assign wr_data_bit_sel[43] = wr_packet[86];
	assign wr_data_bit_sel[44] = wr_packet[86];
	assign wr_data_bit_sel[45] = wr_packet[86];
	assign wr_data_bit_sel[46] = wr_packet[86];
	assign wr_data_bit_sel[47] = wr_packet[86];
	assign wr_data_bit_sel[48] = wr_packet[87];
	assign wr_data_bit_sel[49] = wr_packet[87];
	assign wr_data_bit_sel[50] = wr_packet[87];
	assign wr_data_bit_sel[51] = wr_packet[87];
	assign wr_data_bit_sel[52] = wr_packet[87];
	assign wr_data_bit_sel[53] = wr_packet[87];
	assign wr_data_bit_sel[54] = wr_packet[87];
	assign wr_data_bit_sel[55] = wr_packet[87];
	assign wr_data_bit_sel[56] = wr_packet[88];
	assign wr_data_bit_sel[57] = wr_packet[88];
	assign wr_data_bit_sel[58] = wr_packet[88];
	assign wr_data_bit_sel[59] = wr_packet[88];
	assign wr_data_bit_sel[60] = wr_packet[88];
	assign wr_data_bit_sel[61] = wr_packet[88];
	assign wr_data_bit_sel[62] = wr_packet[88];
	assign wr_data_bit_sel[63] = wr_packet[88];
	always @(*)
		if (wr_packet[89]) begin
			mem_wr_en = 1'h1;
			mem_rd_en = 1'h0;
			mem_addr = wr_packet[80-:17];
			mem_data_in = wr_packet[63-:64];
			mem_data_in_bit_sel = wr_data_bit_sel;
		end
		else if (rdrq_packet[17]) begin
			mem_wr_en = 1'h0;
			mem_rd_en = 1'h1;
			mem_addr = rdrq_packet[16-:17];
			mem_data_in = 64'h0000000000000000;
			mem_data_in_bit_sel = 64'h0000000000000000;
		end
		else begin
			mem_wr_en = 1'h0;
			mem_rd_en = 1'h0;
			mem_addr = 17'h00000;
			mem_data_in = 64'h0000000000000000;
			mem_data_in_bit_sel = 64'h0000000000000000;
		end
	always @(posedge clk or posedge reset)
		if (reset)
			packet_rd_data_r <= 64'h0000000000000000;
		else
			packet_rd_data_r <= rdrs_packet[64-:64];
	always @(*) begin
		if (packet_rd_en_d)
			rdrs_packet[64-:64] = mem_data_out;
		else
			rdrs_packet[64-:64] = packet_rd_data_r;
		rdrs_packet[0] = packet_rd_en_d;
	end
	glb_bank_memory glb_bank_memory(
		.addr(mem_addr),
		.clk(clk),
		.data_in(mem_data_in),
		.data_in_bit_sel(mem_data_in_bit_sel),
		.ren(mem_rd_en),
		.reset(reset),
		.wen(mem_wr_en),
		.data_out(mem_data_out)
	);
	pipeline_w_1_d_1 packet_rdrq_pipeline(
		.clk(clk),
		.clk_en(1'h1),
		.in_(rdrq_packet[17]),
		.reset(reset),
		.out_(packet_rd_en_d)
	);
endmodule
module glb_bank_memory (
	addr,
	clk,
	data_in,
	data_in_bit_sel,
	ren,
	reset,
	wen,
	data_out
);
	input wire [16:0] addr;
	input wire clk;
	input wire [63:0] data_in;
	input wire [63:0] data_in_bit_sel;
	input wire ren;
	input wire reset;
	input wire wen;
	output reg [63:0] data_out;
	wire glb_bank_sram_gen_CEB;
	wire glb_bank_sram_gen_WEB;
	reg [13:0] sram_addr;
	wire [13:0] sram_addr_d;
	reg sram_cen;
	wire sram_cen_d;
	reg [63:0] sram_data_in;
	reg [63:0] sram_data_in_bit_sel;
	wire [63:0] sram_data_in_bit_sel_d;
	wire [63:0] sram_data_in_d;
	wire [63:0] sram_data_out;
	wire [143:0] sram_signals_pipeline_in_;
	wire [143:0] sram_signals_pipeline_out_;
	reg sram_wen;
	wire sram_wen_d;
	assign sram_signals_pipeline_in_ = {sram_wen, sram_cen, sram_addr, sram_data_in, sram_data_in_bit_sel};
	assign {sram_wen_d, sram_cen_d, sram_addr_d, sram_data_in_d, sram_data_in_bit_sel_d} = sram_signals_pipeline_out_;
	assign glb_bank_sram_gen_CEB = ~sram_cen_d;
	assign glb_bank_sram_gen_WEB = ~sram_wen_d;
	always @(*) begin
		sram_wen = wen;
		sram_cen = wen | ren;
		sram_addr = addr[16:3];
		sram_data_in = data_in;
		sram_data_in_bit_sel = data_in_bit_sel;
		data_out = sram_data_out;
	end
	pipeline_w_144_d_0 sram_signals_pipeline(
		.clk(clk),
		.clk_en(1'h1),
		.in_(sram_signals_pipeline_in_),
		.reset(reset),
		.out_(sram_signals_pipeline_out_)
	);
	glb_bank_sram_gen_14 glb_bank_sram_gen(
		.A(sram_addr_d),
		.BW(sram_data_in_bit_sel_d),
		.CEB(glb_bank_sram_gen_CEB),
		.CLK(clk),
		.D(sram_data_in_d),
		.RESET(reset),
		.WEB(glb_bank_sram_gen_WEB),
		.Q(sram_data_out)
	);
endmodule
module glb_bank_mux (
	cfg_pcfg_tile_connected_next,
	cfg_pcfg_tile_connected_prev,
	cfg_tile_connected_next,
	cfg_tile_connected_prev,
	clk,
	glb_tile_id,
	rdrq_packet_dma2bank,
	rdrq_packet_pcfgdma2bank,
	rdrq_packet_pcfgring2bank,
	rdrq_packet_procsw2bank,
	rdrq_packet_ring2bank,
	rdrs_packet_bankarr2sw,
	reset,
	wr_packet_dma2bank,
	wr_packet_procsw2bank,
	wr_packet_ring2bank,
	rdrq_packet_sw2bankarr,
	rdrs_packet_bank2dma,
	rdrs_packet_bank2pcfgdma,
	rdrs_packet_bank2pcfgring,
	rdrs_packet_bank2procsw,
	rdrs_packet_bank2ring,
	wr_packet_sw2bankarr
);
	input wire cfg_pcfg_tile_connected_next;
	input wire cfg_pcfg_tile_connected_prev;
	input wire cfg_tile_connected_next;
	input wire cfg_tile_connected_prev;
	input wire clk;
	input wire glb_tile_id;
	input wire [19:0] rdrq_packet_dma2bank;
	input wire [19:0] rdrq_packet_pcfgdma2bank;
	input wire [19:0] rdrq_packet_pcfgring2bank;
	input wire [19:0] rdrq_packet_procsw2bank;
	input wire [19:0] rdrq_packet_ring2bank;
	input wire [129:0] rdrs_packet_bankarr2sw;
	input wire reset;
	input wire [91:0] wr_packet_dma2bank;
	input wire [91:0] wr_packet_procsw2bank;
	input wire [91:0] wr_packet_ring2bank;
	output wire [35:0] rdrq_packet_sw2bankarr;
	output reg [64:0] rdrs_packet_bank2dma;
	output reg [64:0] rdrs_packet_bank2pcfgdma;
	output reg [64:0] rdrs_packet_bank2pcfgring;
	output reg [64:0] rdrs_packet_bank2procsw;
	output reg [64:0] rdrs_packet_bank2ring;
	output wire [179:0] wr_packet_sw2bankarr;
	reg [1:0] rd_type_0;
	reg [1:0] rd_type_1;
	wire [1:0] rd_type_d_0;
	wire [1:0] rd_type_d_1;
	wire [3:0] rd_type_pipeline_1_in_;
	wire [3:0] rd_type_pipeline_1_out_;
	reg [35:0] rdrq_packet_sw2bankarr_w;
	wire [17:0] rdrq_sw2bank_pipeline_0_out_;
	wire [17:0] rdrq_sw2bank_pipeline_1_out_;
	wire [64:0] rdrs_bank2sw_pipeline_0_out_;
	wire [64:0] rdrs_bank2sw_pipeline_1_out_;
	wire [129:0] rdrs_packet_bankarr2sw_d;
	reg [179:0] wr_packet_sw2bankarr_w;
	wire [89:0] wr_sw2bank_pipeline_0_out_;
	wire [89:0] wr_sw2bank_pipeline_1_out_;
	assign wr_packet_sw2bankarr[0+:90] = wr_sw2bank_pipeline_0_out_;
	assign wr_packet_sw2bankarr[90+:90] = wr_sw2bank_pipeline_1_out_;
	assign rdrq_packet_sw2bankarr[0+:18] = rdrq_sw2bank_pipeline_0_out_;
	assign rdrq_packet_sw2bankarr[18+:18] = rdrq_sw2bank_pipeline_1_out_;
	assign rd_type_pipeline_1_in_ = {rd_type_0, rd_type_1};
	assign {rd_type_d_0, rd_type_d_1} = rd_type_pipeline_1_out_;
	assign rdrs_packet_bankarr2sw_d[0+:65] = rdrs_bank2sw_pipeline_0_out_;
	assign rdrs_packet_bankarr2sw_d[65+:65] = rdrs_bank2sw_pipeline_1_out_;
	always @(*)
		if (((wr_packet_procsw2bank[91] == 1'h1) & (wr_packet_procsw2bank[82] == glb_tile_id)) & (wr_packet_procsw2bank[81] == 1'h0)) begin
			wr_packet_sw2bankarr_w[89] = wr_packet_procsw2bank[91];
			wr_packet_sw2bankarr_w[80-:17] = wr_packet_procsw2bank[80:64];
			wr_packet_sw2bankarr_w[88-:8] = wr_packet_procsw2bank[90-:8];
			wr_packet_sw2bankarr_w[63-:64] = wr_packet_procsw2bank[63-:64];
		end
		else if (((((wr_packet_dma2bank[91] == 1'h1) & ~cfg_tile_connected_prev) & ~cfg_tile_connected_next) & (wr_packet_dma2bank[82] == glb_tile_id)) & (wr_packet_dma2bank[81] == 1'h0)) begin
			wr_packet_sw2bankarr_w[89] = wr_packet_dma2bank[91];
			wr_packet_sw2bankarr_w[80-:17] = wr_packet_dma2bank[80:64];
			wr_packet_sw2bankarr_w[88-:8] = wr_packet_dma2bank[90-:8];
			wr_packet_sw2bankarr_w[63-:64] = wr_packet_dma2bank[63-:64];
		end
		else if (((wr_packet_ring2bank[91] == 1'h1) & (wr_packet_ring2bank[82] == glb_tile_id)) & (wr_packet_ring2bank[81] == 1'h0)) begin
			wr_packet_sw2bankarr_w[89] = wr_packet_ring2bank[91];
			wr_packet_sw2bankarr_w[80-:17] = wr_packet_ring2bank[80:64];
			wr_packet_sw2bankarr_w[88-:8] = wr_packet_ring2bank[90-:8];
			wr_packet_sw2bankarr_w[63-:64] = wr_packet_ring2bank[63-:64];
		end
		else
			wr_packet_sw2bankarr_w[0+:90] = 90'h00000000000000000000000;
	always @(*)
		if (((wr_packet_procsw2bank[91] == 1'h1) & (wr_packet_procsw2bank[82] == glb_tile_id)) & (wr_packet_procsw2bank[81] == 1'h1)) begin
			wr_packet_sw2bankarr_w[179] = wr_packet_procsw2bank[91];
			wr_packet_sw2bankarr_w[170-:17] = wr_packet_procsw2bank[80:64];
			wr_packet_sw2bankarr_w[178-:8] = wr_packet_procsw2bank[90-:8];
			wr_packet_sw2bankarr_w[153-:64] = wr_packet_procsw2bank[63-:64];
		end
		else if (((((wr_packet_dma2bank[91] == 1'h1) & ~cfg_tile_connected_prev) & ~cfg_tile_connected_next) & (wr_packet_dma2bank[82] == glb_tile_id)) & (wr_packet_dma2bank[81] == 1'h1)) begin
			wr_packet_sw2bankarr_w[179] = wr_packet_dma2bank[91];
			wr_packet_sw2bankarr_w[170-:17] = wr_packet_dma2bank[80:64];
			wr_packet_sw2bankarr_w[178-:8] = wr_packet_dma2bank[90-:8];
			wr_packet_sw2bankarr_w[153-:64] = wr_packet_dma2bank[63-:64];
		end
		else if (((wr_packet_ring2bank[91] == 1'h1) & (wr_packet_ring2bank[82] == glb_tile_id)) & (wr_packet_ring2bank[81] == 1'h1)) begin
			wr_packet_sw2bankarr_w[179] = wr_packet_ring2bank[91];
			wr_packet_sw2bankarr_w[170-:17] = wr_packet_ring2bank[80:64];
			wr_packet_sw2bankarr_w[178-:8] = wr_packet_ring2bank[90-:8];
			wr_packet_sw2bankarr_w[153-:64] = wr_packet_ring2bank[63-:64];
		end
		else
			wr_packet_sw2bankarr_w[90+:90] = 90'h00000000000000000000000;
	always @(*)
		if (((rdrq_packet_procsw2bank[19] == 1'h1) & (rdrq_packet_procsw2bank[18] == glb_tile_id)) & (rdrq_packet_procsw2bank[17] == 1'h0)) begin
			rdrq_packet_sw2bankarr_w[17] = rdrq_packet_procsw2bank[19];
			rdrq_packet_sw2bankarr_w[16-:17] = rdrq_packet_procsw2bank[16:0];
			rd_type_0 = 2'h1;
		end
		else if (((((rdrq_packet_pcfgdma2bank[19] == 1'h1) & ~cfg_pcfg_tile_connected_prev) & ~cfg_pcfg_tile_connected_next) & (rdrq_packet_pcfgdma2bank[18] == glb_tile_id)) & (rdrq_packet_pcfgdma2bank[17] == 1'h0)) begin
			rdrq_packet_sw2bankarr_w[17] = rdrq_packet_pcfgdma2bank[19];
			rdrq_packet_sw2bankarr_w[16-:17] = rdrq_packet_pcfgdma2bank[16:0];
			rd_type_0 = 2'h3;
		end
		else if (((rdrq_packet_pcfgring2bank[19] == 1'h1) & (rdrq_packet_pcfgring2bank[18] == glb_tile_id)) & (rdrq_packet_pcfgring2bank[17] == 1'h0)) begin
			rdrq_packet_sw2bankarr_w[17] = rdrq_packet_pcfgring2bank[19];
			rdrq_packet_sw2bankarr_w[16-:17] = rdrq_packet_pcfgring2bank[16:0];
			rd_type_0 = 2'h3;
		end
		else if (((((rdrq_packet_dma2bank[19] == 1'h1) & ~cfg_tile_connected_prev) & ~cfg_tile_connected_next) & (rdrq_packet_dma2bank[18] == glb_tile_id)) & (rdrq_packet_dma2bank[17] == 1'h0)) begin
			rdrq_packet_sw2bankarr_w[17] = rdrq_packet_dma2bank[19];
			rdrq_packet_sw2bankarr_w[16-:17] = rdrq_packet_dma2bank[16:0];
			rd_type_0 = 2'h2;
		end
		else if (((rdrq_packet_ring2bank[19] == 1'h1) & (rdrq_packet_ring2bank[18] == glb_tile_id)) & (rdrq_packet_ring2bank[17] == 1'h0)) begin
			rdrq_packet_sw2bankarr_w[17] = rdrq_packet_ring2bank[19];
			rdrq_packet_sw2bankarr_w[16-:17] = rdrq_packet_ring2bank[16:0];
			rd_type_0 = 2'h2;
		end
		else begin
			rdrq_packet_sw2bankarr_w[0+:18] = 18'h00000;
			rd_type_0 = 2'h0;
		end
	always @(*)
		if (((rdrq_packet_procsw2bank[19] == 1'h1) & (rdrq_packet_procsw2bank[18] == glb_tile_id)) & (rdrq_packet_procsw2bank[17] == 1'h1)) begin
			rdrq_packet_sw2bankarr_w[35] = rdrq_packet_procsw2bank[19];
			rdrq_packet_sw2bankarr_w[34-:17] = rdrq_packet_procsw2bank[16:0];
			rd_type_1 = 2'h1;
		end
		else if (((((rdrq_packet_pcfgdma2bank[19] == 1'h1) & ~cfg_pcfg_tile_connected_prev) & ~cfg_pcfg_tile_connected_next) & (rdrq_packet_pcfgdma2bank[18] == glb_tile_id)) & (rdrq_packet_pcfgdma2bank[17] == 1'h1)) begin
			rdrq_packet_sw2bankarr_w[35] = rdrq_packet_pcfgdma2bank[19];
			rdrq_packet_sw2bankarr_w[34-:17] = rdrq_packet_pcfgdma2bank[16:0];
			rd_type_1 = 2'h3;
		end
		else if (((rdrq_packet_pcfgring2bank[19] == 1'h1) & (rdrq_packet_pcfgring2bank[18] == glb_tile_id)) & (rdrq_packet_pcfgring2bank[17] == 1'h1)) begin
			rdrq_packet_sw2bankarr_w[35] = rdrq_packet_pcfgring2bank[19];
			rdrq_packet_sw2bankarr_w[34-:17] = rdrq_packet_pcfgring2bank[16:0];
			rd_type_1 = 2'h3;
		end
		else if (((((rdrq_packet_dma2bank[19] == 1'h1) & ~cfg_tile_connected_prev) & ~cfg_tile_connected_next) & (rdrq_packet_dma2bank[18] == glb_tile_id)) & (rdrq_packet_dma2bank[17] == 1'h1)) begin
			rdrq_packet_sw2bankarr_w[35] = rdrq_packet_dma2bank[19];
			rdrq_packet_sw2bankarr_w[34-:17] = rdrq_packet_dma2bank[16:0];
			rd_type_1 = 2'h2;
		end
		else if (((rdrq_packet_ring2bank[19] == 1'h1) & (rdrq_packet_ring2bank[18] == glb_tile_id)) & (rdrq_packet_ring2bank[17] == 1'h1)) begin
			rdrq_packet_sw2bankarr_w[35] = rdrq_packet_ring2bank[19];
			rdrq_packet_sw2bankarr_w[34-:17] = rdrq_packet_ring2bank[16:0];
			rd_type_1 = 2'h2;
		end
		else begin
			rdrq_packet_sw2bankarr_w[18+:18] = 18'h00000;
			rd_type_1 = 2'h0;
		end
	always @(*) begin
		rdrs_packet_bank2dma = 65'h00000000000000000;
		if (~cfg_tile_connected_next & ~cfg_tile_connected_prev) begin
			if (rd_type_d_0 == 2'h2)
				rdrs_packet_bank2dma = rdrs_packet_bankarr2sw_d[0+:65];
			if (rd_type_d_1 == 2'h2)
				rdrs_packet_bank2dma = rdrs_packet_bankarr2sw_d[65+:65];
		end
	end
	always @(*) begin
		rdrs_packet_bank2ring = 65'h00000000000000000;
		if (cfg_tile_connected_next | cfg_tile_connected_prev) begin
			if (rd_type_d_0 == 2'h2)
				rdrs_packet_bank2ring = rdrs_packet_bankarr2sw_d[0+:65];
			if (rd_type_d_1 == 2'h2)
				rdrs_packet_bank2ring = rdrs_packet_bankarr2sw_d[65+:65];
		end
	end
	always @(*) begin
		rdrs_packet_bank2procsw = 65'h00000000000000000;
		if (rd_type_d_0 == 2'h1)
			rdrs_packet_bank2procsw = rdrs_packet_bankarr2sw_d[0+:65];
		if (rd_type_d_1 == 2'h1)
			rdrs_packet_bank2procsw = rdrs_packet_bankarr2sw_d[65+:65];
	end
	always @(*) begin
		rdrs_packet_bank2pcfgdma = 65'h00000000000000000;
		if (~cfg_pcfg_tile_connected_next & ~cfg_pcfg_tile_connected_prev) begin
			if (rd_type_d_0 == 2'h3)
				rdrs_packet_bank2pcfgdma = rdrs_packet_bankarr2sw_d[0+:65];
			if (rd_type_d_1 == 2'h3)
				rdrs_packet_bank2pcfgdma = rdrs_packet_bankarr2sw_d[65+:65];
		end
	end
	always @(*) begin
		rdrs_packet_bank2pcfgring = 65'h00000000000000000;
		if (cfg_pcfg_tile_connected_next | cfg_pcfg_tile_connected_prev) begin
			if (rd_type_d_0 == 2'h3)
				rdrs_packet_bank2pcfgring = rdrs_packet_bankarr2sw_d[0+:65];
			if (rd_type_d_1 == 2'h3)
				rdrs_packet_bank2pcfgring = rdrs_packet_bankarr2sw_d[65+:65];
		end
	end
	pipeline_w_90_d_0 wr_sw2bank_pipeline_0(
		.clk(clk),
		.clk_en(1'h1),
		.in_(wr_packet_sw2bankarr_w[0+:90]),
		.reset(reset),
		.out_(wr_sw2bank_pipeline_0_out_)
	);
	pipeline_w_90_d_0 wr_sw2bank_pipeline_1(
		.clk(clk),
		.clk_en(1'h1),
		.in_(wr_packet_sw2bankarr_w[90+:90]),
		.reset(reset),
		.out_(wr_sw2bank_pipeline_1_out_)
	);
	pipeline_w_18_d_0 rdrq_sw2bank_pipeline_0(
		.clk(clk),
		.clk_en(1'h1),
		.in_(rdrq_packet_sw2bankarr_w[0+:18]),
		.reset(reset),
		.out_(rdrq_sw2bank_pipeline_0_out_)
	);
	pipeline_w_18_d_0 rdrq_sw2bank_pipeline_1(
		.clk(clk),
		.clk_en(1'h1),
		.in_(rdrq_packet_sw2bankarr_w[18+:18]),
		.reset(reset),
		.out_(rdrq_sw2bank_pipeline_1_out_)
	);
	pipeline_w_4_d_2 rd_type_pipeline_1(
		.clk(clk),
		.clk_en(1'h1),
		.in_(rd_type_pipeline_1_in_),
		.reset(reset),
		.out_(rd_type_pipeline_1_out_)
	);
	pipeline_w_65_d_1 rdrs_bank2sw_pipeline_0(
		.clk(clk),
		.clk_en(1'h1),
		.in_(rdrs_packet_bankarr2sw[0+:65]),
		.reset(reset),
		.out_(rdrs_bank2sw_pipeline_0_out_)
	);
	pipeline_w_65_d_1 rdrs_bank2sw_pipeline_1(
		.clk(clk),
		.clk_en(1'h1),
		.in_(rdrs_packet_bankarr2sw[65+:65]),
		.reset(reset),
		.out_(rdrs_bank2sw_pipeline_1_out_)
	);
endmodule
module glb_bank_sram_gen_14 (
	A,
	BW,
	CEB,
	CLK,
	D,
	RESET,
	WEB,
	Q
);
	input wire [13:0] A;
	input wire [63:0] BW;
	input wire CEB;
	input wire CLK;
	input wire [63:0] D;
	input wire RESET;
	input wire WEB;
	output wire [63:0] Q;
	wire [11:0] A_SRAM;
	wire [11:0] A_SRAM_d;
	wire [63:0] BW_d;
	reg [3:0] CEB_DEMUX;
	wire [3:0] CEB_DEMUX_d;
	wire CEB_d;
	wire [63:0] D_d;
	reg [1:0] Q_SEL;
	wire [63:0] Q_SRAM2MUX [3:0];
	wire [63:0] Q_w;
	wire [1:0] SRAM_SEL;
	wire [1:0] SRAM_SEL_d;
	reg [3:0] WEB_DEMUX;
	wire [3:0] WEB_DEMUX_d;
	wire WEB_d;
	wire [63:0] sram_array_0_Q;
	wire [63:0] sram_array_1_Q;
	wire [63:0] sram_array_2_Q;
	wire [63:0] sram_array_3_Q;
	wire [77:0] sram_signals_pipeline_in_;
	wire [77:0] sram_signals_pipeline_out_;
	wire [73:0] sram_signals_reset_high_pipeline_in_;
	wire [73:0] sram_signals_reset_high_pipeline_out_;
	assign SRAM_SEL = A[13:12];
	assign A_SRAM = A[11:0];
	assign sram_signals_reset_high_pipeline_in_ = {WEB, CEB, WEB_DEMUX, CEB_DEMUX, BW};
	assign {WEB_d, CEB_d, WEB_DEMUX_d, CEB_DEMUX_d, BW_d} = sram_signals_reset_high_pipeline_out_;
	assign sram_signals_pipeline_in_ = {A_SRAM, SRAM_SEL, D};
	assign {A_SRAM_d, SRAM_SEL_d, D_d} = sram_signals_pipeline_out_;
	always @(posedge CLK or posedge RESET)
		if (RESET)
			Q_SEL <= 2'h0;
		else if ((CEB_d == 1'h0) & (WEB_d == 1'h1))
			Q_SEL <= SRAM_SEL_d;
	function automatic [3:0] sv2v_cast_4;
		input reg [3:0] inp;
		sv2v_cast_4 = inp;
	endfunction
	always @(*) begin
		if (~WEB)
			WEB_DEMUX = ~(4'h1 << sv2v_cast_4(SRAM_SEL));
		else
			WEB_DEMUX = 4'hf;
		if (~CEB)
			CEB_DEMUX = ~(4'h1 << sv2v_cast_4(SRAM_SEL));
		else
			CEB_DEMUX = 4'hf;
	end
	assign Q_SRAM2MUX[0] = sram_array_0_Q;
	assign Q_SRAM2MUX[1] = sram_array_1_Q;
	assign Q_SRAM2MUX[2] = sram_array_2_Q;
	assign Q_SRAM2MUX[3] = sram_array_3_Q;
	assign Q_w = Q_SRAM2MUX[Q_SEL];
	pipeline_w_74_d_0_reset_high sram_signals_reset_high_pipeline(
		.clk(CLK),
		.clk_en(1'h1),
		.in_(sram_signals_reset_high_pipeline_in_),
		.reset(RESET),
		.out_(sram_signals_reset_high_pipeline_out_)
	);
	pipeline_w_78_d_0 sram_signals_pipeline(
		.clk(CLK),
		.clk_en(1'h1),
		.in_(sram_signals_pipeline_in_),
		.reset(RESET),
		.out_(sram_signals_pipeline_out_)
	);
	pipeline_w_64_d_0 sram_signals_output_pipeline(
		.clk(CLK),
		.clk_en(1'h1),
		.in_(Q_w),
		.reset(RESET),
		.out_(Q)
	);
	IN12LP_S1DB_W04096B064M08S2_HB sram_array_0(
		.A(A_SRAM_d),
		.BW(BW_d),
		.CEN(CEB_DEMUX_d[0]),
		.CLK(CLK),
		.D(D_d),
		.MA_SAWL0(1'h0),
		.MA_SAWL1(1'h0),
		.MA_STABAS0(1'h0),
		.MA_STABAS1(1'h0),
		.MA_VD0(1'h0),
		.MA_VD1(1'h0),
		.MA_WL0(1'h0),
		.MA_WL1(1'h0),
		.MA_WRAS0(1'h0),
		.MA_WRAS1(1'h0),
		.MA_WRT(1'h0),
		.RDWEN(WEB_DEMUX_d[0]),
		.T_LOGIC(1'h0),
		.T_Q_RST(1'h0),
		.Q(sram_array_0_Q)
	);
	IN12LP_S1DB_W04096B064M08S2_HB sram_array_1(
		.A(A_SRAM_d),
		.BW(BW_d),
		.CEN(CEB_DEMUX_d[1]),
		.CLK(CLK),
		.D(D_d),
		.MA_SAWL0(1'h0),
		.MA_SAWL1(1'h0),
		.MA_STABAS0(1'h0),
		.MA_STABAS1(1'h0),
		.MA_VD0(1'h0),
		.MA_VD1(1'h0),
		.MA_WL0(1'h0),
		.MA_WL1(1'h0),
		.MA_WRAS0(1'h0),
		.MA_WRAS1(1'h0),
		.MA_WRT(1'h0),
		.RDWEN(WEB_DEMUX_d[1]),
		.T_LOGIC(1'h0),
		.T_Q_RST(1'h0),
		.Q(sram_array_1_Q)
	);
	IN12LP_S1DB_W04096B064M08S2_HB sram_array_2(
		.A(A_SRAM_d),
		.BW(BW_d),
		.CEN(CEB_DEMUX_d[2]),
		.CLK(CLK),
		.D(D_d),
		.MA_SAWL0(1'h0),
		.MA_SAWL1(1'h0),
		.MA_STABAS0(1'h0),
		.MA_STABAS1(1'h0),
		.MA_VD0(1'h0),
		.MA_VD1(1'h0),
		.MA_WL0(1'h0),
		.MA_WL1(1'h0),
		.MA_WRAS0(1'h0),
		.MA_WRAS1(1'h0),
		.MA_WRT(1'h0),
		.RDWEN(WEB_DEMUX_d[2]),
		.T_LOGIC(1'h0),
		.T_Q_RST(1'h0),
		.Q(sram_array_2_Q)
	);
	IN12LP_S1DB_W04096B064M08S2_HB sram_array_3(
		.A(A_SRAM_d),
		.BW(BW_d),
		.CEN(CEB_DEMUX_d[3]),
		.CLK(CLK),
		.D(D_d),
		.MA_SAWL0(1'h0),
		.MA_SAWL1(1'h0),
		.MA_STABAS0(1'h0),
		.MA_STABAS1(1'h0),
		.MA_VD0(1'h0),
		.MA_VD1(1'h0),
		.MA_WL0(1'h0),
		.MA_WL1(1'h0),
		.MA_WRAS0(1'h0),
		.MA_WRAS1(1'h0),
		.MA_WRT(1'h0),
		.RDWEN(WEB_DEMUX_d[3]),
		.T_LOGIC(1'h0),
		.T_Q_RST(1'h0),
		.Q(sram_array_3_Q)
	);
endmodule
module glb_clk_en_gen_11 (
	clk,
	enable,
	reset,
	clk_en
);
	parameter cnt = 32'h0000000b;
	input wire clk;
	input wire enable;
	input wire reset;
	output wire clk_en;
	reg [31:0] clk_en_cnt;
	always @(posedge clk or posedge reset)
		if (reset)
			clk_en_cnt <= 32'h00000000;
		else if (enable)
			clk_en_cnt <= cnt - 32'h00000001;
		else if (clk_en_cnt > 32'h00000000)
			clk_en_cnt <= clk_en_cnt - 32'h00000001;
	assign clk_en = enable | (clk_en_cnt > 32'h00000000);
endmodule
module glb_clk_en_gen_4 (
	clk,
	enable,
	reset,
	clk_en
);
	parameter cnt = 32'h00000004;
	input wire clk;
	input wire enable;
	input wire reset;
	output wire clk_en;
	reg [31:0] clk_en_cnt;
	always @(posedge clk or posedge reset)
		if (reset)
			clk_en_cnt <= 32'h00000000;
		else if (enable)
			clk_en_cnt <= cnt - 32'h00000001;
		else if (clk_en_cnt > 32'h00000000)
			clk_en_cnt <= clk_en_cnt - 32'h00000001;
	assign clk_en = enable | (clk_en_cnt > 32'h00000000);
endmodule
module glb_clk_en_gen_5 (
	clk,
	enable,
	reset,
	clk_en
);
	parameter cnt = 32'h00000005;
	input wire clk;
	input wire enable;
	input wire reset;
	output wire clk_en;
	reg [31:0] clk_en_cnt;
	always @(posedge clk or posedge reset)
		if (reset)
			clk_en_cnt <= 32'h00000000;
		else if (enable)
			clk_en_cnt <= cnt - 32'h00000001;
		else if (clk_en_cnt > 32'h00000000)
			clk_en_cnt <= clk_en_cnt - 32'h00000001;
	assign clk_en = enable | (clk_en_cnt > 32'h00000000);
endmodule
module glb_clk_en_gen_6 (
	clk,
	enable,
	reset,
	clk_en
);
	parameter cnt = 32'h00000006;
	input wire clk;
	input wire enable;
	input wire reset;
	output wire clk_en;
	reg [31:0] clk_en_cnt;
	always @(posedge clk or posedge reset)
		if (reset)
			clk_en_cnt <= 32'h00000000;
		else if (enable)
			clk_en_cnt <= cnt - 32'h00000001;
		else if (clk_en_cnt > 32'h00000000)
			clk_en_cnt <= clk_en_cnt - 32'h00000001;
	assign clk_en = enable | (clk_en_cnt > 32'h00000000);
endmodule
module glb_crossbar_I_2_O_1_W_1 (
	in_,
	sel_,
	out_
);
	input wire [1:0] in_;
	input wire sel_;
	output reg out_;
	always @(*) out_ = in_[sel_];
endmodule
module glb_load_dma (
	cfg_data_network_g2f_mux,
	cfg_data_network_latency,
	cfg_ld_dma_ctrl_flush_mode,
	cfg_ld_dma_ctrl_mode,
	cfg_ld_dma_ctrl_valid_mode,
	cfg_ld_dma_header,
	cfg_ld_dma_num_repeat,
	cfg_tile_connected_next,
	cfg_tile_connected_prev,
	clk,
	data_g2f_rdy,
	glb_tile_id,
	ld_dma_start_pulse,
	rdrs_packet_bank2dma,
	rdrs_packet_ring2dma,
	reset,
	clk_en_dma2bank,
	ctrl_g2f,
	data_flush,
	data_g2f,
	data_g2f_vld,
	ld_dma_done_interrupt,
	rdrq_packet_dma2bank,
	rdrq_packet_dma2ring
);
	input wire [1:0] cfg_data_network_g2f_mux;
	input wire [5:0] cfg_data_network_latency;
	input wire cfg_ld_dma_ctrl_flush_mode;
	input wire [1:0] cfg_ld_dma_ctrl_mode;
	input wire [1:0] cfg_ld_dma_ctrl_valid_mode;
	input wire [582:0] cfg_ld_dma_header;
	input wire cfg_ld_dma_num_repeat;
	input wire cfg_tile_connected_next;
	input wire cfg_tile_connected_prev;
	input wire clk;
	input wire [1:0] data_g2f_rdy;
	input wire glb_tile_id;
	input wire ld_dma_start_pulse;
	input wire [64:0] rdrs_packet_bank2dma;
	input wire [64:0] rdrs_packet_ring2dma;
	input wire reset;
	output wire clk_en_dma2bank;
	output wire [1:0] ctrl_g2f;
	output wire data_flush;
	output wire [31:0] data_g2f;
	output wire [1:0] data_g2f_vld;
	output reg ld_dma_done_interrupt;
	output reg [19:0] rdrq_packet_dma2bank;
	output reg [19:0] rdrq_packet_dma2ring;
	reg all_skid_empty;
	reg [18:0] bank_rdrq_rd_addr;
	reg bank_rdrq_rd_en;
	reg [63:0] bank_rdrs_data_cache_r;
	reg [1:0] ctrl_g2f_w;
	wire [582:0] current_dma_header;
	reg [15:0] cycle_count;
	wire cycle_counter_en;
	wire [15:0] cycle_current_addr;
	wire [127:0] cycle_stride_addr_gen_strides;
	wire cycle_valid;
	wire [19:0] data_current_addr;
	wire [15:0] data_dma2fifo;
	wire [15:0] data_fifo2cgra;
	reg data_flush_w;
	reg [1:0] data_g2f_rdy_muxed;
	wire [15:0] data_g2f_skid_0_data_out;
	wire data_g2f_skid_0_empty;
	wire data_g2f_skid_0_full;
	wire [15:0] data_g2f_skid_1_data_out;
	wire data_g2f_skid_1_empty;
	wire data_g2f_skid_1_full;
	wire [19:0] data_stride_addr_gen_start_addr;
	wire [159:0] data_stride_addr_gen_strides;
	wire dma2bank_clk_en;
	wire [1:0] fifo2skid_rdy;
	reg fifo2skid_rdy_muxed;
	reg [1:0] fifo2skid_vld;
	wire fifo2skid_vld_muxed;
	wire fifo_almost_full;
	reg [4:0] fifo_almost_full_diff;
	wire fifo_empty;
	wire fifo_full;
	wire fifo_pop;
	wire fifo_push;
	wire fifo_push_ready;
	reg is_cached;
	reg is_first;
	reg iter_step_valid;
	reg [18:0] last_strm_rd_addr_r;
	reg ld_dma_done_pulse;
	reg ld_dma_done_pulse_anded;
	wire [23:0] ld_dma_done_pulse_d_arr;
	wire ld_dma_done_pulse_last;
	reg ld_dma_done_pulse_latch;
	wire ld_dma_done_pulse_pipeline_out;
	reg ld_dma_done_pulse_w;
	reg ld_dma_start_pulse_next;
	reg ld_dma_start_pulse_r;
	wire loop_done;
	wire [255:0] loop_iter_ranges;
	wire [2:0] loop_mux_sel;
	wire [1:0] pipeline_ctrl_in;
	wire [1:0] pipeline_ctrl_out;
	reg [19:0] rdrq_packet_dma2bank_w;
	reg [19:0] rdrq_packet_dma2ring_w;
	reg [64:0] rdrs_packet;
	reg repeat_cnt;
	wire [1:0] skid_empty;
	wire [1:0] skid_full;
	reg [31:0] skid_in;
	wire [31:0] skid_out;
	wire [1:0] skid_pop;
	wire [1:0] skid_push;
	reg strm_ctrl_muxed;
	reg [15:0] strm_data;
	wire [43:0] strm_data_sel_arr;
	wire [1:0] strm_data_sel_w;
	wire strm_data_start_pulse;
	wire [21:0] strm_data_start_pulse_d_arr;
	wire strm_data_valid;
	reg [18:0] strm_rd_addr_w;
	wire [21:0] strm_rd_en_d_arr;
	reg strm_rd_en_w;
	reg strm_run;
	assign fifo_push_ready = ~fifo_almost_full;
	assign data_dma2fifo = strm_data;
	assign fifo_push = ~fifo_full & strm_data_valid;
	assign fifo2skid_vld_muxed = ~fifo_empty;
	assign fifo_pop = fifo2skid_vld_muxed & fifo2skid_rdy_muxed;
	function automatic [4:0] sv2v_cast_5;
		input reg [4:0] inp;
		sv2v_cast_5 = inp;
	endfunction
	always @(*) fifo_almost_full_diff = sv2v_cast_5(6'h05 + cfg_data_network_latency);
	assign skid_out[0+:16] = data_g2f_skid_0_data_out;
	assign skid_full[0] = data_g2f_skid_0_full;
	assign skid_empty[0] = data_g2f_skid_0_empty;
	assign data_g2f[0+:16] = skid_out[0+:16];
	assign fifo2skid_rdy[0] = ~skid_full[0];
	assign skid_push[0] = fifo2skid_rdy[0] & fifo2skid_vld[0];
	assign data_g2f_vld[0] = ~skid_empty[0];
	assign skid_pop[0] = ~skid_empty[0] & data_g2f_rdy_muxed[0];
	assign skid_out[16+:16] = data_g2f_skid_1_data_out;
	assign skid_full[1] = data_g2f_skid_1_full;
	assign skid_empty[1] = data_g2f_skid_1_empty;
	assign data_g2f[16+:16] = skid_out[16+:16];
	assign fifo2skid_rdy[1] = ~skid_full[1];
	assign skid_push[1] = fifo2skid_rdy[1] & fifo2skid_vld[1];
	assign data_g2f_vld[1] = ~skid_empty[1];
	assign skid_pop[1] = ~skid_empty[1] & data_g2f_rdy_muxed[1];
	always @(*) begin
		fifo2skid_rdy_muxed = 1'h0;
		if (cfg_data_network_g2f_mux[0] == 1'h1) begin
			fifo2skid_rdy_muxed = fifo2skid_rdy[0];
			fifo2skid_vld[0] = fifo2skid_vld_muxed;
			skid_in[0+:16] = data_fifo2cgra;
		end
		else begin
			fifo2skid_rdy_muxed = fifo2skid_rdy_muxed;
			fifo2skid_vld[0] = 1'h0;
			skid_in[0+:16] = 16'h0000;
		end
		if (cfg_data_network_g2f_mux[1] == 1'h1) begin
			fifo2skid_rdy_muxed = fifo2skid_rdy[1];
			fifo2skid_vld[1] = fifo2skid_vld_muxed;
			skid_in[16+:16] = data_fifo2cgra;
		end
		else begin
			fifo2skid_rdy_muxed = fifo2skid_rdy_muxed;
			fifo2skid_vld[1] = 1'h0;
			skid_in[16+:16] = 16'h0000;
		end
	end
	always @(*) begin
		if (cfg_ld_dma_ctrl_valid_mode == 2'h2)
			data_g2f_rdy_muxed[0] = data_g2f_rdy[0];
		else
			data_g2f_rdy_muxed[0] = 1'h1;
		if (cfg_ld_dma_ctrl_valid_mode == 2'h2)
			data_g2f_rdy_muxed[1] = data_g2f_rdy[1];
		else
			data_g2f_rdy_muxed[1] = 1'h1;
	end
	always @(*) begin
		all_skid_empty = 1'h1;
		if (cfg_data_network_g2f_mux[0])
			all_skid_empty = all_skid_empty & skid_empty[0];
		else
			all_skid_empty = all_skid_empty;
		if (cfg_data_network_g2f_mux[1])
			all_skid_empty = all_skid_empty & skid_empty[1];
		else
			all_skid_empty = all_skid_empty;
	end
	assign current_dma_header = cfg_ld_dma_header;
	always @(*)
		if (cycle_counter_en)
			iter_step_valid = cycle_valid;
		else
			iter_step_valid = strm_run & fifo_push_ready;
	always @(posedge clk or posedge reset)
		if (reset)
			repeat_cnt <= 1'h0;
		else if (cfg_ld_dma_ctrl_mode == 2'h2) begin
			if (ld_dma_done_pulse) begin
				if ((repeat_cnt + 1'h1) < cfg_ld_dma_num_repeat)
					repeat_cnt <= repeat_cnt + 1'h1;
			end
		end
		else if (cfg_ld_dma_ctrl_mode == 2'h3) begin
			if (ld_dma_done_pulse) begin
				if (((repeat_cnt + 1'h1) < cfg_ld_dma_num_repeat) & ((repeat_cnt + 1'h1) < 1'h1))
					repeat_cnt <= repeat_cnt + 1'h1;
			end
		end
	always @(posedge clk or posedge reset)
		if (reset)
			cycle_count <= 16'h0000;
		else if (ld_dma_start_pulse_r)
			cycle_count <= 16'h0000;
		else if (loop_done)
			cycle_count <= 16'h0000;
		else if (cycle_counter_en & strm_run)
			cycle_count <= cycle_count + 16'h0001;
	always @(posedge clk or posedge reset)
		if (reset)
			is_first <= 1'h0;
		else if (ld_dma_start_pulse_r)
			is_first <= 1'h1;
		else if (bank_rdrq_rd_en)
			is_first <= 1'h0;
	always @(posedge clk or posedge reset)
		if (reset)
			strm_run <= 1'h0;
		else if (ld_dma_start_pulse_r)
			strm_run <= 1'h1;
		else if (loop_done)
			strm_run <= 1'h0;
	assign strm_data_start_pulse = strm_data_start_pulse_d_arr[sv2v_cast_5(cfg_data_network_latency) + 5'h03];
	assign strm_data_valid = strm_rd_en_d_arr[sv2v_cast_5(cfg_data_network_latency) + 5'h03];
	assign strm_data_sel_w = strm_rd_addr_w[2:1];
	always @(*)
		if (cfg_ld_dma_ctrl_mode == 2'h0)
			ld_dma_start_pulse_next = 1'h0;
		else if (cfg_ld_dma_ctrl_mode == 2'h1)
			ld_dma_start_pulse_next = ~strm_run & ld_dma_start_pulse;
		else if ((cfg_ld_dma_ctrl_mode == 2'h2) | (cfg_ld_dma_ctrl_mode == 2'h3))
			ld_dma_start_pulse_next = (~strm_run & ld_dma_start_pulse) | (ld_dma_done_pulse & ((repeat_cnt + 1'h1) < cfg_ld_dma_num_repeat));
		else
			ld_dma_start_pulse_next = 1'h0;
	always @(posedge clk or posedge reset)
		if (reset)
			ld_dma_start_pulse_r <= 1'h0;
		else if (ld_dma_start_pulse_r)
			ld_dma_start_pulse_r <= 1'h0;
		else
			ld_dma_start_pulse_r <= ld_dma_start_pulse_next;
	always @(*)
		if (cfg_ld_dma_ctrl_flush_mode == 1'h0) begin
			data_flush_w = strm_data_start_pulse;
			if (cfg_ld_dma_ctrl_valid_mode == 2'h1)
				strm_ctrl_muxed = strm_data_valid;
			else
				strm_ctrl_muxed = 1'h0;
		end
		else begin
			data_flush_w = 1'h0;
			if (cfg_ld_dma_ctrl_valid_mode == 2'h1)
				strm_ctrl_muxed = strm_data_valid;
			else
				strm_ctrl_muxed = strm_data_start_pulse;
		end
	always @(*) begin
		if (cfg_data_network_g2f_mux[0] == 1'h1) begin
			if (cfg_ld_dma_ctrl_valid_mode != 2'h2)
				ctrl_g2f_w[0] = strm_ctrl_muxed;
			else
				ctrl_g2f_w[0] = 1'h0;
		end
		else
			ctrl_g2f_w[0] = 1'h0;
		if (cfg_data_network_g2f_mux[1] == 1'h1) begin
			if (cfg_ld_dma_ctrl_valid_mode != 2'h2)
				ctrl_g2f_w[1] = strm_ctrl_muxed;
			else
				ctrl_g2f_w[1] = 1'h0;
		end
		else
			ctrl_g2f_w[1] = 1'h0;
	end
	always @(*) ld_dma_done_pulse_w = strm_run & loop_done;
	function automatic [18:0] sv2v_cast_19;
		input reg [18:0] inp;
		sv2v_cast_19 = inp;
	endfunction
	always @(*) begin
		strm_rd_en_w = iter_step_valid;
		strm_rd_addr_w = sv2v_cast_19(data_current_addr);
	end
	always @(posedge clk or posedge reset)
		if (reset)
			last_strm_rd_addr_r <= 19'h00000;
		else if (strm_rd_en_w)
			last_strm_rd_addr_r <= strm_rd_addr_w;
	always @(*)
		if (cfg_tile_connected_next | cfg_tile_connected_prev) begin
			rdrq_packet_dma2bank_w = 20'h00000;
			rdrq_packet_dma2ring_w[19] = bank_rdrq_rd_en;
			rdrq_packet_dma2ring_w[18-:19] = bank_rdrq_rd_addr;
		end
		else begin
			rdrq_packet_dma2bank_w[19] = bank_rdrq_rd_en;
			rdrq_packet_dma2bank_w[18-:19] = bank_rdrq_rd_addr;
			rdrq_packet_dma2ring_w = 20'h00000;
		end
	always @(posedge clk or posedge reset)
		if (reset) begin
			rdrq_packet_dma2bank <= 20'h00000;
			rdrq_packet_dma2ring <= 20'h00000;
		end
		else begin
			rdrq_packet_dma2bank <= rdrq_packet_dma2bank_w;
			rdrq_packet_dma2ring <= rdrq_packet_dma2ring_w;
		end
	always @(*) begin
		is_cached = strm_rd_addr_w[18:3] == last_strm_rd_addr_r[18:3];
		bank_rdrq_rd_en = strm_rd_en_w & (is_first | ~is_cached);
		bank_rdrq_rd_addr = strm_rd_addr_w;
	end
	always @(*)
		if (cfg_tile_connected_next | cfg_tile_connected_prev)
			rdrs_packet = rdrs_packet_ring2dma;
		else
			rdrs_packet = rdrs_packet_bank2dma;
	always @(posedge clk or posedge reset)
		if (reset)
			bank_rdrs_data_cache_r <= 64'h0000000000000000;
		else if (rdrs_packet[0])
			bank_rdrs_data_cache_r <= rdrs_packet[64-:64];
	always @(*)
		case (strm_data_sel_arr[(sv2v_cast_5(cfg_data_network_latency) + 5'h03) * 2+:2])
			2'h0: strm_data = bank_rdrs_data_cache_r[15:0];
			2'h1: strm_data = bank_rdrs_data_cache_r[31:16];
			2'h2: strm_data = bank_rdrs_data_cache_r[47:32];
			2'h3: strm_data = bank_rdrs_data_cache_r[63:48];
			default: strm_data = bank_rdrs_data_cache_r[15:0];
		endcase
	always @(posedge clk or posedge reset)
		if (reset)
			ld_dma_done_pulse_latch <= 1'h0;
		else if (ld_dma_done_pulse_pipeline_out)
			ld_dma_done_pulse_latch <= 1'h1;
		else if (ld_dma_done_pulse_latch & all_skid_empty)
			ld_dma_done_pulse_latch <= 1'h0;
	always @(*)
		if (cfg_ld_dma_ctrl_valid_mode != 2'h2)
			ld_dma_done_pulse = ld_dma_done_pulse_pipeline_out;
		else
			ld_dma_done_pulse = ld_dma_done_pulse_anded;
	always @(*) ld_dma_done_pulse_anded = ld_dma_done_pulse_latch & all_skid_empty;
	assign ld_dma_done_pulse_pipeline_out = ld_dma_done_pulse_d_arr[sv2v_cast_5(cfg_data_network_latency) + (5'h03 + 5'h02)];
	always @(posedge clk or posedge reset)
		if (reset)
			ld_dma_done_interrupt <= 1'h0;
		else if (ld_dma_done_pulse)
			ld_dma_done_interrupt <= 1'h1;
		else if (ld_dma_done_pulse_last)
			ld_dma_done_interrupt <= 1'h0;
	assign clk_en_dma2bank = dma2bank_clk_en;
	assign pipeline_ctrl_in[0] = ctrl_g2f_w[0];
	assign pipeline_ctrl_in[1] = ctrl_g2f_w[1];
	assign ctrl_g2f[0] = pipeline_ctrl_out[0];
	assign ctrl_g2f[1] = pipeline_ctrl_out[1];
	assign loop_iter_ranges[0+:32] = current_dma_header[543-:32];
	assign loop_iter_ranges[32+:32] = current_dma_header[475-:32];
	assign loop_iter_ranges[64+:32] = current_dma_header[407-:32];
	assign loop_iter_ranges[96+:32] = current_dma_header[339-:32];
	assign loop_iter_ranges[128+:32] = current_dma_header[271-:32];
	assign loop_iter_ranges[160+:32] = current_dma_header[203-:32];
	assign loop_iter_ranges[192+:32] = current_dma_header[135-:32];
	assign loop_iter_ranges[224+:32] = current_dma_header[67-:32];
	assign cycle_counter_en = cfg_ld_dma_ctrl_valid_mode != 2'h2;
	assign cycle_stride_addr_gen_strides[0+:16] = current_dma_header[491-:16];
	assign cycle_stride_addr_gen_strides[16+:16] = current_dma_header[423-:16];
	assign cycle_stride_addr_gen_strides[32+:16] = current_dma_header[355-:16];
	assign cycle_stride_addr_gen_strides[48+:16] = current_dma_header[287-:16];
	assign cycle_stride_addr_gen_strides[64+:16] = current_dma_header[219-:16];
	assign cycle_stride_addr_gen_strides[80+:16] = current_dma_header[151-:16];
	assign cycle_stride_addr_gen_strides[96+:16] = current_dma_header[83-:16];
	assign cycle_stride_addr_gen_strides[112+:16] = current_dma_header[15-:16];
	function automatic [19:0] sv2v_cast_20;
		input reg [19:0] inp;
		sv2v_cast_20 = inp;
	endfunction
	assign data_stride_addr_gen_start_addr = sv2v_cast_20(current_dma_header[582-:19]);
	assign data_stride_addr_gen_strides[0+:20] = current_dma_header[511-:20];
	assign data_stride_addr_gen_strides[20+:20] = current_dma_header[443-:20];
	assign data_stride_addr_gen_strides[40+:20] = current_dma_header[375-:20];
	assign data_stride_addr_gen_strides[60+:20] = current_dma_header[307-:20];
	assign data_stride_addr_gen_strides[80+:20] = current_dma_header[239-:20];
	assign data_stride_addr_gen_strides[100+:20] = current_dma_header[171-:20];
	assign data_stride_addr_gen_strides[120+:20] = current_dma_header[103-:20];
	assign data_stride_addr_gen_strides[140+:20] = current_dma_header[35-:20];
	reg_fifo_d_19_w_16 #(.data_width(16'h0010)) data_g2f_fifo(
		.almost_empty_diff(5'h02),
		.almost_full_diff(fifo_almost_full_diff),
		.clk(clk),
		.clk_en(1'h1),
		.data_in(data_dma2fifo),
		.flush(ld_dma_start_pulse_r),
		.pop(fifo_pop),
		.push(fifo_push),
		.reset(reset),
		.almost_full(fifo_almost_full),
		.data_out(data_fifo2cgra),
		.empty(fifo_empty),
		.full(fifo_full)
	);
	reg_fifo_d_2_w_16 #(.data_width(16'h0010)) data_g2f_skid_0(
		.almost_empty_diff(1'h0),
		.almost_full_diff(1'h0),
		.clk(clk),
		.clk_en(1'h1),
		.data_in(skid_in[0+:16]),
		.flush(ld_dma_start_pulse_r),
		.pop(skid_pop[0]),
		.push(skid_push[0]),
		.reset(reset),
		.data_out(data_g2f_skid_0_data_out),
		.empty(data_g2f_skid_0_empty),
		.full(data_g2f_skid_0_full)
	);
	reg_fifo_d_2_w_16 #(.data_width(16'h0010)) data_g2f_skid_1(
		.almost_empty_diff(1'h0),
		.almost_full_diff(1'h0),
		.clk(clk),
		.clk_en(1'h1),
		.data_in(skid_in[16+:16]),
		.flush(ld_dma_start_pulse_r),
		.pop(skid_pop[1]),
		.push(skid_push[1]),
		.reset(reset),
		.data_out(data_g2f_skid_1_data_out),
		.empty(data_g2f_skid_1_empty),
		.full(data_g2f_skid_1_full)
	);
	pipeline_w_1_d_22_array strm_dma_start_pulse_pipeline(
		.clk(clk),
		.clk_en(1'h1),
		.in_(ld_dma_start_pulse_r),
		.reset(reset),
		.out_(strm_data_start_pulse_d_arr)
	);
	pipeline_w_1_d_22_array strm_rd_en_pipeline(
		.clk(clk),
		.clk_en(1'h1),
		.in_(strm_rd_en_w),
		.reset(reset),
		.out_(strm_rd_en_d_arr)
	);
	pipeline_w_2_d_22_array strm_data_sel_pipeline(
		.clk(clk),
		.clk_en(1'h1),
		.in_(strm_data_sel_w),
		.reset(reset),
		.out_(strm_data_sel_arr)
	);
	pipeline_w_1_d_24_array ld_dma_done_pulse_pipeline(
		.clk(clk),
		.clk_en(1'h1),
		.in_(ld_dma_done_pulse_w),
		.reset(reset),
		.out_(ld_dma_done_pulse_d_arr)
	);
	pipeline_w_1_d_5 ld_dma_interrupt_pipeline(
		.clk(clk),
		.clk_en(1'h1),
		.in_(ld_dma_done_pulse),
		.reset(reset),
		.out_(ld_dma_done_pulse_last)
	);
	glb_clk_en_gen_6 #(.cnt(32'h00000006)) dma2bank_clk_en_gen(
		.clk(clk),
		.enable(rdrq_packet_dma2bank_w[19]),
		.reset(reset),
		.clk_en(dma2bank_clk_en)
	);
	pipeline_w_2_d_2 pipeline_ctrl(
		.clk(clk),
		.clk_en(1'h1),
		.in_(pipeline_ctrl_in),
		.reset(reset),
		.out_(pipeline_ctrl_out)
	);
	pipeline_w_1_d_0 pipeline_flush(
		.clk(clk),
		.clk_en(1'h1),
		.in_(data_flush_w),
		.reset(reset),
		.out_(data_flush)
	);
	glb_loop_iter_8 loop_iter(
		.clk(clk),
		.clk_en(1'h1),
		.dim(current_dma_header[547-:4]),
		.ranges(loop_iter_ranges),
		.reset(reset),
		.step(iter_step_valid),
		.mux_sel_out(loop_mux_sel),
		.restart(loop_done)
	);
	glb_sched_gen cycle_stride_sched_gen(
		.clk(clk),
		.clk_en(cycle_counter_en),
		.current_addr(cycle_current_addr),
		.cycle_count(cycle_count),
		.finished(loop_done),
		.reset(reset),
		.restart(ld_dma_start_pulse_r),
		.valid_output(cycle_valid)
	);
	glb_addr_gen_8 #(
		.addr_width(32'h00000010),
		.loop_level(32'h00000008)
	) cycle_stride_addr_gen(
		.clk(clk),
		.clk_en(cycle_counter_en),
		.mux_sel(loop_mux_sel),
		.reset(reset),
		.restart(ld_dma_start_pulse_r),
		.start_addr(current_dma_header[563-:16]),
		.step(iter_step_valid),
		.strides(cycle_stride_addr_gen_strides),
		.addr_out(cycle_current_addr)
	);
	glb_addr_gen_8 #(
		.addr_width(32'h00000014),
		.loop_level(32'h00000008)
	) data_stride_addr_gen(
		.clk(clk),
		.clk_en(1'h1),
		.mux_sel(loop_mux_sel),
		.reset(reset),
		.restart(ld_dma_start_pulse_r),
		.start_addr(data_stride_addr_gen_start_addr),
		.step(iter_step_valid),
		.strides(data_stride_addr_gen_strides),
		.addr_out(data_current_addr)
	);
endmodule
module glb_loop_iter_7 (
	clk,
	clk_en,
	dim,
	ranges,
	reset,
	step,
	mux_sel_out,
	restart
);
	input wire clk;
	input wire clk_en;
	input wire [3:0] dim;
	input wire [223:0] ranges;
	input wire reset;
	input wire step;
	output wire [2:0] mux_sel_out;
	output wire restart;
	reg [6:0] clear;
	reg [223:0] dim_counter;
	reg [6:0] inc;
	wire is_maxed;
	reg [6:0] max_value;
	reg [2:0] mux_sel;
	reg not_done;
	assign mux_sel_out = mux_sel;
	assign is_maxed = (dim_counter[mux_sel * 32+:32] == ranges[mux_sel * 32+:32]) & inc[mux_sel];
	function automatic [2:0] sv2v_cast_3;
		input reg [2:0] inp;
		sv2v_cast_3 = inp;
	endfunction
	function automatic [3:0] sv2v_cast_4;
		input reg [3:0] inp;
		sv2v_cast_4 = inp;
	endfunction
	always @(*) begin
		mux_sel = 3'h0;
		not_done = 1'h0;
		begin : sv2v_autoblock_1
			reg [31:0] i;
			for (i = 0; i < 7; i = i + 1)
				if (~not_done) begin
					if (~max_value[sv2v_cast_3(i)] & (sv2v_cast_4(i) < dim)) begin
						mux_sel = sv2v_cast_3(i);
						not_done = 1'h1;
					end
				end
		end
	end
	always @(*) begin
		clear[0] = 1'h0;
		if (((mux_sel > 3'h0) | ~not_done) & step)
			clear[0] = 1'h1;
	end
	always @(*) begin
		inc[0] = 1'h0;
		if ((1'd1 & step) & (dim > 4'h0))
			inc[0] = 1'h1;
		else if (((mux_sel == 3'h0) & step) & (dim > 4'h0))
			inc[0] = 1'h1;
	end
	always @(posedge clk or posedge reset)
		if (reset)
			dim_counter[0+:32] <= 32'h00000000;
		else if (clear[0])
			dim_counter[0+:32] <= 32'h00000000;
		else if (inc[0])
			dim_counter[0+:32] <= dim_counter[mux_sel * 32+:32] + 32'h00000001;
	always @(posedge clk or posedge reset)
		if (reset)
			max_value[0] <= 1'h0;
		else if (clk_en) begin
			if (clear[0])
				max_value[0] <= 1'h0;
			else if (inc[0])
				max_value[0] <= is_maxed;
		end
	always @(*) begin
		clear[1] = 1'h0;
		if (((mux_sel > 3'h1) | ~not_done) & step)
			clear[1] = 1'h1;
	end
	always @(*) begin
		inc[1] = 1'h0;
		if ((1'd0 & step) & (dim > 4'h1))
			inc[1] = 1'h1;
		else if (((mux_sel == 3'h1) & step) & (dim > 4'h1))
			inc[1] = 1'h1;
	end
	always @(posedge clk or posedge reset)
		if (reset)
			dim_counter[32+:32] <= 32'h00000000;
		else if (clear[1])
			dim_counter[32+:32] <= 32'h00000000;
		else if (inc[1])
			dim_counter[32+:32] <= dim_counter[mux_sel * 32+:32] + 32'h00000001;
	always @(posedge clk or posedge reset)
		if (reset)
			max_value[1] <= 1'h0;
		else if (clk_en) begin
			if (clear[1])
				max_value[1] <= 1'h0;
			else if (inc[1])
				max_value[1] <= is_maxed;
		end
	always @(*) begin
		clear[2] = 1'h0;
		if (((mux_sel > 3'h2) | ~not_done) & step)
			clear[2] = 1'h1;
	end
	always @(*) begin
		inc[2] = 1'h0;
		if ((1'd0 & step) & (dim > 4'h2))
			inc[2] = 1'h1;
		else if (((mux_sel == 3'h2) & step) & (dim > 4'h2))
			inc[2] = 1'h1;
	end
	always @(posedge clk or posedge reset)
		if (reset)
			dim_counter[64+:32] <= 32'h00000000;
		else if (clear[2])
			dim_counter[64+:32] <= 32'h00000000;
		else if (inc[2])
			dim_counter[64+:32] <= dim_counter[mux_sel * 32+:32] + 32'h00000001;
	always @(posedge clk or posedge reset)
		if (reset)
			max_value[2] <= 1'h0;
		else if (clk_en) begin
			if (clear[2])
				max_value[2] <= 1'h0;
			else if (inc[2])
				max_value[2] <= is_maxed;
		end
	always @(*) begin
		clear[3] = 1'h0;
		if (((mux_sel > 3'h3) | ~not_done) & step)
			clear[3] = 1'h1;
	end
	always @(*) begin
		inc[3] = 1'h0;
		if ((1'd0 & step) & (dim > 4'h3))
			inc[3] = 1'h1;
		else if (((mux_sel == 3'h3) & step) & (dim > 4'h3))
			inc[3] = 1'h1;
	end
	always @(posedge clk or posedge reset)
		if (reset)
			dim_counter[96+:32] <= 32'h00000000;
		else if (clear[3])
			dim_counter[96+:32] <= 32'h00000000;
		else if (inc[3])
			dim_counter[96+:32] <= dim_counter[mux_sel * 32+:32] + 32'h00000001;
	always @(posedge clk or posedge reset)
		if (reset)
			max_value[3] <= 1'h0;
		else if (clk_en) begin
			if (clear[3])
				max_value[3] <= 1'h0;
			else if (inc[3])
				max_value[3] <= is_maxed;
		end
	always @(*) begin
		clear[4] = 1'h0;
		if (((mux_sel > 3'h4) | ~not_done) & step)
			clear[4] = 1'h1;
	end
	always @(*) begin
		inc[4] = 1'h0;
		if ((1'd0 & step) & (dim > 4'h4))
			inc[4] = 1'h1;
		else if (((mux_sel == 3'h4) & step) & (dim > 4'h4))
			inc[4] = 1'h1;
	end
	always @(posedge clk or posedge reset)
		if (reset)
			dim_counter[128+:32] <= 32'h00000000;
		else if (clear[4])
			dim_counter[128+:32] <= 32'h00000000;
		else if (inc[4])
			dim_counter[128+:32] <= dim_counter[mux_sel * 32+:32] + 32'h00000001;
	always @(posedge clk or posedge reset)
		if (reset)
			max_value[4] <= 1'h0;
		else if (clk_en) begin
			if (clear[4])
				max_value[4] <= 1'h0;
			else if (inc[4])
				max_value[4] <= is_maxed;
		end
	always @(*) begin
		clear[5] = 1'h0;
		if (((mux_sel > 3'h5) | ~not_done) & step)
			clear[5] = 1'h1;
	end
	always @(*) begin
		inc[5] = 1'h0;
		if ((1'd0 & step) & (dim > 4'h5))
			inc[5] = 1'h1;
		else if (((mux_sel == 3'h5) & step) & (dim > 4'h5))
			inc[5] = 1'h1;
	end
	always @(posedge clk or posedge reset)
		if (reset)
			dim_counter[160+:32] <= 32'h00000000;
		else if (clear[5])
			dim_counter[160+:32] <= 32'h00000000;
		else if (inc[5])
			dim_counter[160+:32] <= dim_counter[mux_sel * 32+:32] + 32'h00000001;
	always @(posedge clk or posedge reset)
		if (reset)
			max_value[5] <= 1'h0;
		else if (clk_en) begin
			if (clear[5])
				max_value[5] <= 1'h0;
			else if (inc[5])
				max_value[5] <= is_maxed;
		end
	always @(*) begin
		clear[6] = 1'h0;
		if (((mux_sel > 3'h6) | ~not_done) & step)
			clear[6] = 1'h1;
	end
	always @(*) begin
		inc[6] = 1'h0;
		if ((1'd0 & step) & (dim > 4'h6))
			inc[6] = 1'h1;
		else if (((mux_sel == 3'h6) & step) & (dim > 4'h6))
			inc[6] = 1'h1;
	end
	always @(posedge clk or posedge reset)
		if (reset)
			dim_counter[192+:32] <= 32'h00000000;
		else if (clear[6])
			dim_counter[192+:32] <= 32'h00000000;
		else if (inc[6])
			dim_counter[192+:32] <= dim_counter[mux_sel * 32+:32] + 32'h00000001;
	always @(posedge clk or posedge reset)
		if (reset)
			max_value[6] <= 1'h0;
		else if (clk_en) begin
			if (clear[6])
				max_value[6] <= 1'h0;
			else if (inc[6])
				max_value[6] <= is_maxed;
		end
	assign restart = step & ~not_done;
endmodule
module glb_loop_iter_8 (
	clk,
	clk_en,
	dim,
	ranges,
	reset,
	step,
	mux_sel_out,
	restart
);
	input wire clk;
	input wire clk_en;
	input wire [3:0] dim;
	input wire [255:0] ranges;
	input wire reset;
	input wire step;
	output wire [2:0] mux_sel_out;
	output wire restart;
	reg [7:0] clear;
	reg [255:0] dim_counter;
	reg [7:0] inc;
	wire is_maxed;
	reg [7:0] max_value;
	reg [2:0] mux_sel;
	reg not_done;
	assign mux_sel_out = mux_sel;
	assign is_maxed = (dim_counter[mux_sel * 32+:32] == ranges[mux_sel * 32+:32]) & inc[mux_sel];
	function automatic [2:0] sv2v_cast_3;
		input reg [2:0] inp;
		sv2v_cast_3 = inp;
	endfunction
	function automatic [3:0] sv2v_cast_4;
		input reg [3:0] inp;
		sv2v_cast_4 = inp;
	endfunction
	always @(*) begin
		mux_sel = 3'h0;
		not_done = 1'h0;
		begin : sv2v_autoblock_1
			reg [31:0] i;
			for (i = 0; i < 8; i = i + 1)
				if (~not_done) begin
					if (~max_value[sv2v_cast_3(i)] & (sv2v_cast_4(i) < dim)) begin
						mux_sel = sv2v_cast_3(i);
						not_done = 1'h1;
					end
				end
		end
	end
	always @(*) begin
		clear[0] = 1'h0;
		if (((mux_sel > 3'h0) | ~not_done) & step)
			clear[0] = 1'h1;
	end
	always @(*) begin
		inc[0] = 1'h0;
		if ((1'd1 & step) & (dim > 4'h0))
			inc[0] = 1'h1;
		else if (((mux_sel == 3'h0) & step) & (dim > 4'h0))
			inc[0] = 1'h1;
	end
	always @(posedge clk or posedge reset)
		if (reset)
			dim_counter[0+:32] <= 32'h00000000;
		else if (clear[0])
			dim_counter[0+:32] <= 32'h00000000;
		else if (inc[0])
			dim_counter[0+:32] <= dim_counter[mux_sel * 32+:32] + 32'h00000001;
	always @(posedge clk or posedge reset)
		if (reset)
			max_value[0] <= 1'h0;
		else if (clk_en) begin
			if (clear[0])
				max_value[0] <= 1'h0;
			else if (inc[0])
				max_value[0] <= is_maxed;
		end
	always @(*) begin
		clear[1] = 1'h0;
		if (((mux_sel > 3'h1) | ~not_done) & step)
			clear[1] = 1'h1;
	end
	always @(*) begin
		inc[1] = 1'h0;
		if ((1'd0 & step) & (dim > 4'h1))
			inc[1] = 1'h1;
		else if (((mux_sel == 3'h1) & step) & (dim > 4'h1))
			inc[1] = 1'h1;
	end
	always @(posedge clk or posedge reset)
		if (reset)
			dim_counter[32+:32] <= 32'h00000000;
		else if (clear[1])
			dim_counter[32+:32] <= 32'h00000000;
		else if (inc[1])
			dim_counter[32+:32] <= dim_counter[mux_sel * 32+:32] + 32'h00000001;
	always @(posedge clk or posedge reset)
		if (reset)
			max_value[1] <= 1'h0;
		else if (clk_en) begin
			if (clear[1])
				max_value[1] <= 1'h0;
			else if (inc[1])
				max_value[1] <= is_maxed;
		end
	always @(*) begin
		clear[2] = 1'h0;
		if (((mux_sel > 3'h2) | ~not_done) & step)
			clear[2] = 1'h1;
	end
	always @(*) begin
		inc[2] = 1'h0;
		if ((1'd0 & step) & (dim > 4'h2))
			inc[2] = 1'h1;
		else if (((mux_sel == 3'h2) & step) & (dim > 4'h2))
			inc[2] = 1'h1;
	end
	always @(posedge clk or posedge reset)
		if (reset)
			dim_counter[64+:32] <= 32'h00000000;
		else if (clear[2])
			dim_counter[64+:32] <= 32'h00000000;
		else if (inc[2])
			dim_counter[64+:32] <= dim_counter[mux_sel * 32+:32] + 32'h00000001;
	always @(posedge clk or posedge reset)
		if (reset)
			max_value[2] <= 1'h0;
		else if (clk_en) begin
			if (clear[2])
				max_value[2] <= 1'h0;
			else if (inc[2])
				max_value[2] <= is_maxed;
		end
	always @(*) begin
		clear[3] = 1'h0;
		if (((mux_sel > 3'h3) | ~not_done) & step)
			clear[3] = 1'h1;
	end
	always @(*) begin
		inc[3] = 1'h0;
		if ((1'd0 & step) & (dim > 4'h3))
			inc[3] = 1'h1;
		else if (((mux_sel == 3'h3) & step) & (dim > 4'h3))
			inc[3] = 1'h1;
	end
	always @(posedge clk or posedge reset)
		if (reset)
			dim_counter[96+:32] <= 32'h00000000;
		else if (clear[3])
			dim_counter[96+:32] <= 32'h00000000;
		else if (inc[3])
			dim_counter[96+:32] <= dim_counter[mux_sel * 32+:32] + 32'h00000001;
	always @(posedge clk or posedge reset)
		if (reset)
			max_value[3] <= 1'h0;
		else if (clk_en) begin
			if (clear[3])
				max_value[3] <= 1'h0;
			else if (inc[3])
				max_value[3] <= is_maxed;
		end
	always @(*) begin
		clear[4] = 1'h0;
		if (((mux_sel > 3'h4) | ~not_done) & step)
			clear[4] = 1'h1;
	end
	always @(*) begin
		inc[4] = 1'h0;
		if ((1'd0 & step) & (dim > 4'h4))
			inc[4] = 1'h1;
		else if (((mux_sel == 3'h4) & step) & (dim > 4'h4))
			inc[4] = 1'h1;
	end
	always @(posedge clk or posedge reset)
		if (reset)
			dim_counter[128+:32] <= 32'h00000000;
		else if (clear[4])
			dim_counter[128+:32] <= 32'h00000000;
		else if (inc[4])
			dim_counter[128+:32] <= dim_counter[mux_sel * 32+:32] + 32'h00000001;
	always @(posedge clk or posedge reset)
		if (reset)
			max_value[4] <= 1'h0;
		else if (clk_en) begin
			if (clear[4])
				max_value[4] <= 1'h0;
			else if (inc[4])
				max_value[4] <= is_maxed;
		end
	always @(*) begin
		clear[5] = 1'h0;
		if (((mux_sel > 3'h5) | ~not_done) & step)
			clear[5] = 1'h1;
	end
	always @(*) begin
		inc[5] = 1'h0;
		if ((1'd0 & step) & (dim > 4'h5))
			inc[5] = 1'h1;
		else if (((mux_sel == 3'h5) & step) & (dim > 4'h5))
			inc[5] = 1'h1;
	end
	always @(posedge clk or posedge reset)
		if (reset)
			dim_counter[160+:32] <= 32'h00000000;
		else if (clear[5])
			dim_counter[160+:32] <= 32'h00000000;
		else if (inc[5])
			dim_counter[160+:32] <= dim_counter[mux_sel * 32+:32] + 32'h00000001;
	always @(posedge clk or posedge reset)
		if (reset)
			max_value[5] <= 1'h0;
		else if (clk_en) begin
			if (clear[5])
				max_value[5] <= 1'h0;
			else if (inc[5])
				max_value[5] <= is_maxed;
		end
	always @(*) begin
		clear[6] = 1'h0;
		if (((mux_sel > 3'h6) | ~not_done) & step)
			clear[6] = 1'h1;
	end
	always @(*) begin
		inc[6] = 1'h0;
		if ((1'd0 & step) & (dim > 4'h6))
			inc[6] = 1'h1;
		else if (((mux_sel == 3'h6) & step) & (dim > 4'h6))
			inc[6] = 1'h1;
	end
	always @(posedge clk or posedge reset)
		if (reset)
			dim_counter[192+:32] <= 32'h00000000;
		else if (clear[6])
			dim_counter[192+:32] <= 32'h00000000;
		else if (inc[6])
			dim_counter[192+:32] <= dim_counter[mux_sel * 32+:32] + 32'h00000001;
	always @(posedge clk or posedge reset)
		if (reset)
			max_value[6] <= 1'h0;
		else if (clk_en) begin
			if (clear[6])
				max_value[6] <= 1'h0;
			else if (inc[6])
				max_value[6] <= is_maxed;
		end
	always @(*) begin
		clear[7] = 1'h0;
		if (((mux_sel > 3'h7) | ~not_done) & step)
			clear[7] = 1'h1;
	end
	always @(*) begin
		inc[7] = 1'h0;
		if ((1'd0 & step) & (dim > 4'h7))
			inc[7] = 1'h1;
		else if (((mux_sel == 3'h7) & step) & (dim > 4'h7))
			inc[7] = 1'h1;
	end
	always @(posedge clk or posedge reset)
		if (reset)
			dim_counter[224+:32] <= 32'h00000000;
		else if (clear[7])
			dim_counter[224+:32] <= 32'h00000000;
		else if (inc[7])
			dim_counter[224+:32] <= dim_counter[mux_sel * 32+:32] + 32'h00000001;
	always @(posedge clk or posedge reset)
		if (reset)
			max_value[7] <= 1'h0;
		else if (clk_en) begin
			if (clear[7])
				max_value[7] <= 1'h0;
			else if (inc[7])
				max_value[7] <= is_maxed;
		end
	assign restart = step & ~not_done;
endmodule
module glb_pcfg_broadcast (
	cfg_pcfg_broadcast_mux,
	cgra_cfg_dma2mux,
	cgra_cfg_jtag_addr_bypass_wsti,
	cgra_cfg_jtag_rd_en_bypass_wsti,
	cgra_cfg_jtag_wsti,
	cgra_cfg_pcfg_esti,
	cgra_cfg_pcfg_wsti,
	clk,
	reset,
	cgra_cfg_g2f,
	cgra_cfg_jtag_addr_bypass_esto,
	cgra_cfg_jtag_esto,
	cgra_cfg_jtag_rd_en_bypass_esto,
	cgra_cfg_pcfg_esto,
	cgra_cfg_pcfg_wsto
);
	input wire [5:0] cfg_pcfg_broadcast_mux;
	input wire [65:0] cgra_cfg_dma2mux;
	input wire [31:0] cgra_cfg_jtag_addr_bypass_wsti;
	input wire cgra_cfg_jtag_rd_en_bypass_wsti;
	input wire [65:0] cgra_cfg_jtag_wsti;
	input wire [65:0] cgra_cfg_pcfg_esti;
	input wire [65:0] cgra_cfg_pcfg_wsti;
	input wire clk;
	input wire reset;
	output reg [131:0] cgra_cfg_g2f;
	output reg [31:0] cgra_cfg_jtag_addr_bypass_esto;
	output reg [65:0] cgra_cfg_jtag_esto;
	output reg cgra_cfg_jtag_rd_en_bypass_esto;
	output reg [65:0] cgra_cfg_pcfg_esto;
	output reg [65:0] cgra_cfg_pcfg_wsto;
	reg [131:0] cgra_cfg_g2f_w;
	reg [65:0] pcfg_east_muxed;
	reg [65:0] pcfg_south_muxed;
	reg [65:0] pcfg_west_muxed;
	always @(*) begin
		cgra_cfg_jtag_rd_en_bypass_esto = cgra_cfg_jtag_rd_en_bypass_wsti;
		cgra_cfg_jtag_addr_bypass_esto = cgra_cfg_jtag_addr_bypass_wsti;
	end
	always @(*)
		if (cfg_pcfg_broadcast_mux[1-:2] == 2'h0)
			pcfg_south_muxed = 66'h00000000000000000;
		else if (cfg_pcfg_broadcast_mux[1-:2] == 2'h1)
			pcfg_south_muxed = cgra_cfg_dma2mux;
		else if (cfg_pcfg_broadcast_mux[1-:2] == 2'h2)
			pcfg_south_muxed = cgra_cfg_pcfg_wsti;
		else if (cfg_pcfg_broadcast_mux[1-:2] == 2'h3)
			pcfg_south_muxed = cgra_cfg_pcfg_esti;
		else
			pcfg_south_muxed = 66'h00000000000000000;
	always @(*)
		if (cfg_pcfg_broadcast_mux[5-:2] == 2'h0)
			pcfg_west_muxed = 66'h00000000000000000;
		else if (cfg_pcfg_broadcast_mux[5-:2] == 2'h1)
			pcfg_west_muxed = cgra_cfg_dma2mux;
		else if (cfg_pcfg_broadcast_mux[5-:2] == 2'h2)
			pcfg_west_muxed = cgra_cfg_pcfg_esti;
		else
			pcfg_west_muxed = 66'h00000000000000000;
	always @(*)
		if (cfg_pcfg_broadcast_mux[3-:2] == 2'h0)
			pcfg_east_muxed = 66'h00000000000000000;
		else if (cfg_pcfg_broadcast_mux[3-:2] == 2'h1)
			pcfg_east_muxed = cgra_cfg_dma2mux;
		else if (cfg_pcfg_broadcast_mux[3-:2] == 2'h2)
			pcfg_east_muxed = cgra_cfg_pcfg_wsti;
		else
			pcfg_east_muxed = 66'h00000000000000000;
	always @(posedge clk or posedge reset)
		if (reset)
			cgra_cfg_jtag_esto <= 66'h00000000000000000;
		else
			cgra_cfg_jtag_esto <= cgra_cfg_jtag_wsti;
	always @(posedge clk or posedge reset)
		if (reset) begin
			cgra_cfg_pcfg_esto <= 66'h00000000000000000;
			cgra_cfg_pcfg_wsto <= 66'h00000000000000000;
		end
		else begin
			cgra_cfg_pcfg_esto <= pcfg_east_muxed;
			cgra_cfg_pcfg_wsto <= pcfg_west_muxed;
		end
	always @(*)
		if (cgra_cfg_jtag_rd_en_bypass_esto) begin
			cgra_cfg_g2f_w[64] = 1'h0;
			cgra_cfg_g2f_w[65] = 1'h1;
			cgra_cfg_g2f_w[63-:32] = cgra_cfg_jtag_addr_bypass_esto;
			cgra_cfg_g2f_w[31-:32] = 32'h00000000;
		end
		else
			cgra_cfg_g2f_w[0+:66] = cgra_cfg_jtag_wsti | pcfg_south_muxed;
	always @(*)
		if (cgra_cfg_jtag_rd_en_bypass_esto) begin
			cgra_cfg_g2f_w[130] = 1'h0;
			cgra_cfg_g2f_w[131] = 1'h1;
			cgra_cfg_g2f_w[129-:32] = cgra_cfg_jtag_addr_bypass_esto;
			cgra_cfg_g2f_w[97-:32] = 32'h00000000;
		end
		else
			cgra_cfg_g2f_w[66+:66] = cgra_cfg_jtag_wsti | pcfg_south_muxed;
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	always @(posedge clk or posedge reset)
		if (reset) begin : sv2v_autoblock_1
			reg [31:0] i;
			for (i = 0; i < 2; i = i + 1)
				cgra_cfg_g2f[sv2v_cast_1(i) * 66+:66] <= 66'h00000000000000000;
		end
		else begin : sv2v_autoblock_2
			reg [31:0] i;
			for (i = 0; i < 2; i = i + 1)
				cgra_cfg_g2f[sv2v_cast_1(i) * 66+:66] <= cgra_cfg_g2f_w[sv2v_cast_1(i) * 66+:66];
		end
endmodule
module glb_pcfg_dma (
	cfg_pcfg_dma_ctrl_mode,
	cfg_pcfg_dma_ctrl_relocation_is_msb,
	cfg_pcfg_dma_ctrl_relocation_value,
	cfg_pcfg_dma_header,
	cfg_pcfg_network_latency,
	cfg_pcfg_tile_connected_next,
	cfg_pcfg_tile_connected_prev,
	clk,
	glb_tile_id,
	pcfg_dma_start_pulse,
	rdrs_packet_bank2dma,
	rdrs_packet_ring2dma,
	reset,
	cgra_cfg_pcfg,
	clk_en_dma2bank,
	pcfg_dma_done_interrupt,
	rdrq_packet_dma2bank,
	rdrq_packet_dma2ring
);
	input wire cfg_pcfg_dma_ctrl_mode;
	input wire cfg_pcfg_dma_ctrl_relocation_is_msb;
	input wire [15:0] cfg_pcfg_dma_ctrl_relocation_value;
	input wire [34:0] cfg_pcfg_dma_header;
	input wire [5:0] cfg_pcfg_network_latency;
	input wire cfg_pcfg_tile_connected_next;
	input wire cfg_pcfg_tile_connected_prev;
	input wire clk;
	input wire glb_tile_id;
	input wire pcfg_dma_start_pulse;
	input wire [64:0] rdrs_packet_bank2dma;
	input wire [64:0] rdrs_packet_ring2dma;
	input wire reset;
	output reg [65:0] cgra_cfg_pcfg;
	output wire clk_en_dma2bank;
	output reg pcfg_dma_done_interrupt;
	output reg [19:0] rdrq_packet_dma2bank;
	output reg [19:0] rdrq_packet_dma2ring;
	reg [18:0] addr_next;
	reg [18:0] addr_r;
	wire dma2bank_clk_en;
	wire [11:0] done_pulse_d_arr;
	reg done_pulse_r;
	reg is_running_r;
	reg [15:0] num_cfg_cnt_next;
	reg [15:0] num_cfg_cnt_r;
	wire pcfg_done_pulse;
	wire pcfg_done_pulse_last;
	reg [19:0] rdrq_packet_dma2bank_w;
	reg [19:0] rdrq_packet_dma2ring_w;
	reg [18:0] rdrq_packet_rd_addr_next;
	reg rdrq_packet_rd_en_next;
	reg [64:0] rdrs_packet;
	reg [63:0] rdrs_packet_rd_data_r;
	reg rdrs_packet_rd_data_valid_r;
	reg start_pulse_r;
	always @(posedge clk or posedge reset)
		if (reset)
			start_pulse_r <= 1'h0;
		else if (((cfg_pcfg_dma_ctrl_mode == 1'h1) & ~is_running_r) & pcfg_dma_start_pulse)
			start_pulse_r <= 1'h1;
		else
			start_pulse_r <= 1'h0;
	always @(posedge clk or posedge reset)
		if (reset)
			done_pulse_r <= 1'h0;
		else if (is_running_r & (num_cfg_cnt_r == 16'h0000))
			done_pulse_r <= 1'h1;
		else
			done_pulse_r <= 1'h0;
	always @(posedge clk or posedge reset)
		if (reset)
			is_running_r <= 1'h0;
		else if (start_pulse_r)
			is_running_r <= 1'h1;
		else if ((is_running_r == 1'h1) & (num_cfg_cnt_r == 16'h0000))
			is_running_r <= 1'h0;
	always @(*)
		if (start_pulse_r) begin
			num_cfg_cnt_next = cfg_pcfg_dma_header[15-:16];
			addr_next = cfg_pcfg_dma_header[34-:19];
		end
		else if ((is_running_r == 1'h1) & (num_cfg_cnt_r > 16'h0000)) begin
			num_cfg_cnt_next = num_cfg_cnt_r - 16'h0001;
			addr_next = addr_r + 19'h00008;
		end
		else begin
			num_cfg_cnt_next = 16'h0000;
			addr_next = 19'h00000;
		end
	always @(posedge clk or posedge reset)
		if (reset) begin
			num_cfg_cnt_r <= 16'h0000;
			addr_r <= 19'h00000;
		end
		else begin
			num_cfg_cnt_r <= num_cfg_cnt_next;
			addr_r <= addr_next;
		end
	always @(*)
		if (is_running_r & (num_cfg_cnt_r > 16'h0000)) begin
			rdrq_packet_rd_en_next = 1'h1;
			rdrq_packet_rd_addr_next = addr_r;
		end
		else begin
			rdrq_packet_rd_en_next = 1'h0;
			rdrq_packet_rd_addr_next = 19'h00000;
		end
	always @(posedge clk or posedge reset)
		if (reset) begin
			rdrq_packet_dma2ring <= 20'h00000;
			rdrq_packet_dma2bank <= 20'h00000;
		end
		else begin
			rdrq_packet_dma2ring <= rdrq_packet_dma2ring_w;
			rdrq_packet_dma2bank <= rdrq_packet_dma2bank_w;
		end
	always @(posedge clk or posedge reset)
		if (reset) begin
			rdrs_packet_rd_data_r <= 64'h0000000000000000;
			rdrs_packet_rd_data_valid_r <= 1'h0;
		end
		else if (rdrs_packet[0]) begin
			rdrs_packet_rd_data_r <= rdrs_packet[64-:64];
			rdrs_packet_rd_data_valid_r <= 1'h1;
		end
		else begin
			rdrs_packet_rd_data_r <= 64'h0000000000000000;
			rdrs_packet_rd_data_valid_r <= 1'h0;
		end
	always @(*)
		if (cfg_pcfg_tile_connected_next | cfg_pcfg_tile_connected_prev) begin
			rdrq_packet_dma2ring_w[19] = rdrq_packet_rd_en_next;
			rdrq_packet_dma2ring_w[18-:19] = rdrq_packet_rd_addr_next;
			rdrq_packet_dma2bank_w[19] = 1'h0;
			rdrq_packet_dma2bank_w[18-:19] = 19'h00000;
		end
		else begin
			rdrq_packet_dma2ring_w[19] = 1'h0;
			rdrq_packet_dma2ring_w[18-:19] = 19'h00000;
			rdrq_packet_dma2bank_w[19] = rdrq_packet_rd_en_next;
			rdrq_packet_dma2bank_w[18-:19] = rdrq_packet_rd_addr_next;
		end
	always @(*)
		if (cfg_pcfg_tile_connected_next | cfg_pcfg_tile_connected_prev)
			rdrs_packet = rdrs_packet_ring2dma;
		else
			rdrs_packet = rdrs_packet_bank2dma;
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	always @(*) begin
		cgra_cfg_pcfg[65] = 1'h0;
		cgra_cfg_pcfg[64] = rdrs_packet_rd_data_valid_r;
		cgra_cfg_pcfg[31-:32] = rdrs_packet_rd_data_r[31:0];
		if (cfg_pcfg_dma_ctrl_relocation_is_msb)
			cgra_cfg_pcfg[63-:32] = rdrs_packet_rd_data_r[63:32] + sv2v_cast_32(cfg_pcfg_dma_ctrl_relocation_value << 16'h0010);
		else
			cgra_cfg_pcfg[63-:32] = rdrs_packet_rd_data_r[63:32] + sv2v_cast_32(cfg_pcfg_dma_ctrl_relocation_value);
	end
	function automatic [3:0] sv2v_cast_4;
		input reg [3:0] inp;
		sv2v_cast_4 = inp;
	endfunction
	assign pcfg_done_pulse = done_pulse_d_arr[sv2v_cast_4(cfg_pcfg_network_latency) + (4'h3 + 4'h2)];
	always @(posedge clk or posedge reset)
		if (reset)
			pcfg_dma_done_interrupt <= 1'h0;
		else if (pcfg_done_pulse)
			pcfg_dma_done_interrupt <= 1'h1;
		else if (pcfg_done_pulse_last)
			pcfg_dma_done_interrupt <= 1'h0;
	assign clk_en_dma2bank = dma2bank_clk_en;
	pipeline_w_1_d_12_array done_pulse_pipeline(
		.clk(clk),
		.clk_en(1'h1),
		.in_(done_pulse_r),
		.reset(reset),
		.out_(done_pulse_d_arr)
	);
	pipeline_w_1_d_5 pcfg_dma_interrupt_pipeline(
		.clk(clk),
		.clk_en(1'h1),
		.in_(pcfg_done_pulse),
		.reset(reset),
		.out_(pcfg_done_pulse_last)
	);
	glb_clk_en_gen_6 #(.cnt(32'h00000006)) dma2bank_clk_en_gen(
		.clk(clk),
		.enable(rdrq_packet_dma2bank_w[19]),
		.reset(reset),
		.clk_en(dma2bank_clk_en)
	);
endmodule
module glb_ring_switch_RD (
	cfg_ld_dma_on,
	cfg_tile_connected_next,
	cfg_tile_connected_prev,
	clk,
	glb_tile_id,
	rdrq_packet_dma2ring,
	rdrq_packet_e2w_esti,
	rdrq_packet_w2e_wsti,
	rdrs_packet_bank2ring,
	rdrs_packet_e2w_esti,
	rdrs_packet_w2e_wsti,
	reset,
	clk_en_ring2bank,
	rdrq_packet_e2w_wsto,
	rdrq_packet_ring2bank,
	rdrq_packet_w2e_esto,
	rdrs_packet_e2w_wsto,
	rdrs_packet_ring2dma,
	rdrs_packet_w2e_esto
);
	input wire cfg_ld_dma_on;
	input wire cfg_tile_connected_next;
	input wire cfg_tile_connected_prev;
	input wire clk;
	input wire glb_tile_id;
	input wire [19:0] rdrq_packet_dma2ring;
	input wire [19:0] rdrq_packet_e2w_esti;
	input wire [19:0] rdrq_packet_w2e_wsti;
	input wire [64:0] rdrs_packet_bank2ring;
	input wire [64:0] rdrs_packet_e2w_esti;
	input wire [64:0] rdrs_packet_w2e_wsti;
	input wire reset;
	output wire clk_en_ring2bank;
	output reg [19:0] rdrq_packet_e2w_wsto;
	output reg [19:0] rdrq_packet_ring2bank;
	output reg [19:0] rdrq_packet_w2e_esto;
	output reg [64:0] rdrs_packet_e2w_wsto;
	output reg [64:0] rdrs_packet_ring2dma;
	output reg [64:0] rdrs_packet_w2e_esto;
	reg [19:0] rdrq_packet_e2w_esti_muxed;
	reg [19:0] rdrq_packet_e2w_wsto_w;
	reg [19:0] rdrq_packet_ring2bank_w;
	reg [19:0] rdrq_packet_w2e_esto_w;
	reg [19:0] rdrq_packet_w2e_wsti_muxed;
	reg [64:0] rdrs_packet_e2w_esti_muxed;
	reg [64:0] rdrs_packet_e2w_wsto_w;
	reg [64:0] rdrs_packet_ring2dma_w;
	reg [64:0] rdrs_packet_w2e_esto_w;
	reg [64:0] rdrs_packet_w2e_wsti_muxed;
	wire ring2bank_rd_clk_en;
	always @(*)
		if (cfg_tile_connected_prev) begin
			rdrq_packet_w2e_wsti_muxed = rdrq_packet_w2e_wsti;
			rdrs_packet_w2e_wsti_muxed = rdrs_packet_w2e_wsti;
		end
		else begin
			rdrq_packet_w2e_wsti_muxed = rdrq_packet_e2w_wsto;
			rdrs_packet_w2e_wsti_muxed = rdrs_packet_e2w_wsto;
		end
	always @(*)
		if (cfg_tile_connected_next) begin
			rdrq_packet_e2w_esti_muxed = rdrq_packet_e2w_esti;
			rdrs_packet_e2w_esti_muxed = rdrs_packet_e2w_esti;
		end
		else begin
			rdrq_packet_e2w_esti_muxed = rdrq_packet_w2e_esto;
			rdrs_packet_e2w_esti_muxed = rdrs_packet_w2e_esto;
		end
	always @(*) begin
		if (rdrq_packet_dma2ring[19] == 1'h1) begin
			if (rdrq_packet_dma2ring[18] == glb_tile_id) begin
				rdrq_packet_ring2bank_w = rdrq_packet_dma2ring;
				rdrq_packet_w2e_esto_w = 20'h00000;
			end
			else begin
				rdrq_packet_ring2bank_w = 20'h00000;
				rdrq_packet_w2e_esto_w = rdrq_packet_dma2ring;
			end
		end
		else if (rdrq_packet_w2e_wsti_muxed[19] == 1'h1) begin
			if (rdrq_packet_w2e_wsti_muxed[18] == glb_tile_id) begin
				rdrq_packet_ring2bank_w = rdrq_packet_w2e_wsti_muxed;
				rdrq_packet_w2e_esto_w = 20'h00000;
			end
			else begin
				rdrq_packet_ring2bank_w = 20'h00000;
				rdrq_packet_w2e_esto_w = rdrq_packet_w2e_wsti_muxed;
			end
		end
		else begin
			rdrq_packet_ring2bank_w = 20'h00000;
			rdrq_packet_w2e_esto_w = 20'h00000;
		end
		rdrq_packet_e2w_wsto_w = rdrq_packet_e2w_esti_muxed;
	end
	always @(*) begin
		if (rdrs_packet_bank2ring[0] == 1'h1)
			rdrs_packet_w2e_esto_w = rdrs_packet_bank2ring;
		else if (rdrs_packet_w2e_wsti_muxed[0] & cfg_ld_dma_on)
			rdrs_packet_w2e_esto_w = 65'h00000000000000000;
		else
			rdrs_packet_w2e_esto_w = rdrs_packet_w2e_wsti_muxed;
		if (rdrs_packet_w2e_wsti_muxed[0] & cfg_ld_dma_on)
			rdrs_packet_ring2dma_w = rdrs_packet_w2e_wsti_muxed;
		else
			rdrs_packet_ring2dma_w = 65'h00000000000000000;
		rdrs_packet_e2w_wsto_w = rdrs_packet_e2w_esti_muxed;
	end
	always @(posedge clk or posedge reset)
		if (reset) begin
			rdrq_packet_w2e_esto <= 20'h00000;
			rdrq_packet_e2w_wsto <= 20'h00000;
			rdrq_packet_ring2bank <= 20'h00000;
			rdrs_packet_w2e_esto <= 65'h00000000000000000;
			rdrs_packet_e2w_wsto <= 65'h00000000000000000;
		end
		else begin
			rdrq_packet_w2e_esto <= rdrq_packet_w2e_esto_w;
			rdrq_packet_e2w_wsto <= rdrq_packet_e2w_wsto_w;
			rdrq_packet_ring2bank <= rdrq_packet_ring2bank_w;
			rdrs_packet_w2e_esto <= rdrs_packet_w2e_esto_w;
			rdrs_packet_e2w_wsto <= rdrs_packet_e2w_wsto_w;
		end
	always @(*) rdrs_packet_ring2dma = rdrs_packet_ring2dma_w;
	assign clk_en_ring2bank = ring2bank_rd_clk_en;
	glb_clk_en_gen_6 #(.cnt(32'h00000006)) ring2bank_rd_clk_en_gen(
		.clk(clk),
		.enable(rdrq_packet_ring2bank_w[19]),
		.reset(reset),
		.clk_en(ring2bank_rd_clk_en)
	);
endmodule
module glb_ring_switch_WR_RD (
	cfg_ld_dma_on,
	cfg_tile_connected_next,
	cfg_tile_connected_prev,
	clk,
	glb_tile_id,
	rdrq_packet_dma2ring,
	rdrq_packet_e2w_esti,
	rdrq_packet_w2e_wsti,
	rdrs_packet_bank2ring,
	rdrs_packet_e2w_esti,
	rdrs_packet_w2e_wsti,
	reset,
	wr_packet_dma2ring,
	wr_packet_e2w_esti,
	wr_packet_w2e_wsti,
	clk_en_ring2bank,
	rdrq_packet_e2w_wsto,
	rdrq_packet_ring2bank,
	rdrq_packet_w2e_esto,
	rdrs_packet_e2w_wsto,
	rdrs_packet_ring2dma,
	rdrs_packet_w2e_esto,
	wr_packet_e2w_wsto,
	wr_packet_ring2bank,
	wr_packet_w2e_esto
);
	input wire cfg_ld_dma_on;
	input wire cfg_tile_connected_next;
	input wire cfg_tile_connected_prev;
	input wire clk;
	input wire glb_tile_id;
	input wire [19:0] rdrq_packet_dma2ring;
	input wire [19:0] rdrq_packet_e2w_esti;
	input wire [19:0] rdrq_packet_w2e_wsti;
	input wire [64:0] rdrs_packet_bank2ring;
	input wire [64:0] rdrs_packet_e2w_esti;
	input wire [64:0] rdrs_packet_w2e_wsti;
	input wire reset;
	input wire [91:0] wr_packet_dma2ring;
	input wire [91:0] wr_packet_e2w_esti;
	input wire [91:0] wr_packet_w2e_wsti;
	output wire clk_en_ring2bank;
	output reg [19:0] rdrq_packet_e2w_wsto;
	output reg [19:0] rdrq_packet_ring2bank;
	output reg [19:0] rdrq_packet_w2e_esto;
	output reg [64:0] rdrs_packet_e2w_wsto;
	output reg [64:0] rdrs_packet_ring2dma;
	output reg [64:0] rdrs_packet_w2e_esto;
	output reg [91:0] wr_packet_e2w_wsto;
	output reg [91:0] wr_packet_ring2bank;
	output reg [91:0] wr_packet_w2e_esto;
	reg [19:0] rdrq_packet_e2w_esti_muxed;
	reg [19:0] rdrq_packet_e2w_wsto_w;
	reg [19:0] rdrq_packet_ring2bank_w;
	reg [19:0] rdrq_packet_w2e_esto_w;
	reg [19:0] rdrq_packet_w2e_wsti_muxed;
	reg [64:0] rdrs_packet_e2w_esti_muxed;
	reg [64:0] rdrs_packet_e2w_wsto_w;
	reg [64:0] rdrs_packet_ring2dma_w;
	reg [64:0] rdrs_packet_w2e_esto_w;
	reg [64:0] rdrs_packet_w2e_wsti_muxed;
	wire ring2bank_rd_clk_en;
	wire ring2bank_wr_clk_en;
	reg [91:0] wr_packet_e2w_esti_muxed;
	reg [91:0] wr_packet_e2w_wsto_w;
	reg [91:0] wr_packet_ring2bank_w;
	reg [91:0] wr_packet_w2e_esto_w;
	reg [91:0] wr_packet_w2e_wsti_muxed;
	always @(*)
		if (cfg_tile_connected_prev) begin
			wr_packet_w2e_wsti_muxed = wr_packet_w2e_wsti;
			rdrq_packet_w2e_wsti_muxed = rdrq_packet_w2e_wsti;
			rdrs_packet_w2e_wsti_muxed = rdrs_packet_w2e_wsti;
		end
		else begin
			wr_packet_w2e_wsti_muxed = wr_packet_e2w_wsto;
			rdrq_packet_w2e_wsti_muxed = rdrq_packet_e2w_wsto;
			rdrs_packet_w2e_wsti_muxed = rdrs_packet_e2w_wsto;
		end
	always @(*)
		if (cfg_tile_connected_next) begin
			wr_packet_e2w_esti_muxed = wr_packet_e2w_esti;
			rdrq_packet_e2w_esti_muxed = rdrq_packet_e2w_esti;
			rdrs_packet_e2w_esti_muxed = rdrs_packet_e2w_esti;
		end
		else begin
			wr_packet_e2w_esti_muxed = wr_packet_w2e_esto;
			rdrq_packet_e2w_esti_muxed = rdrq_packet_w2e_esto;
			rdrs_packet_e2w_esti_muxed = rdrs_packet_w2e_esto;
		end
	always @(*) begin
		if (wr_packet_dma2ring[91] == 1'h1) begin
			if (wr_packet_dma2ring[82] == glb_tile_id) begin
				wr_packet_ring2bank_w = wr_packet_dma2ring;
				wr_packet_w2e_esto_w = 92'h00000000000000000000000;
			end
			else begin
				wr_packet_ring2bank_w = 92'h00000000000000000000000;
				wr_packet_w2e_esto_w = wr_packet_dma2ring;
			end
		end
		else if (wr_packet_w2e_wsti_muxed[91] == 1'h1) begin
			if (wr_packet_w2e_wsti_muxed[82] == glb_tile_id) begin
				wr_packet_ring2bank_w = wr_packet_w2e_wsti_muxed;
				wr_packet_w2e_esto_w = 92'h00000000000000000000000;
			end
			else begin
				wr_packet_ring2bank_w = 92'h00000000000000000000000;
				wr_packet_w2e_esto_w = wr_packet_w2e_wsti_muxed;
			end
		end
		else begin
			wr_packet_ring2bank_w = 92'h00000000000000000000000;
			wr_packet_w2e_esto_w = 92'h00000000000000000000000;
		end
		wr_packet_e2w_wsto_w = wr_packet_e2w_esti_muxed;
	end
	always @(*) begin
		if (rdrq_packet_dma2ring[19] == 1'h1) begin
			if (rdrq_packet_dma2ring[18] == glb_tile_id) begin
				rdrq_packet_ring2bank_w = rdrq_packet_dma2ring;
				rdrq_packet_w2e_esto_w = 20'h00000;
			end
			else begin
				rdrq_packet_ring2bank_w = 20'h00000;
				rdrq_packet_w2e_esto_w = rdrq_packet_dma2ring;
			end
		end
		else if (rdrq_packet_w2e_wsti_muxed[19] == 1'h1) begin
			if (rdrq_packet_w2e_wsti_muxed[18] == glb_tile_id) begin
				rdrq_packet_ring2bank_w = rdrq_packet_w2e_wsti_muxed;
				rdrq_packet_w2e_esto_w = 20'h00000;
			end
			else begin
				rdrq_packet_ring2bank_w = 20'h00000;
				rdrq_packet_w2e_esto_w = rdrq_packet_w2e_wsti_muxed;
			end
		end
		else begin
			rdrq_packet_ring2bank_w = 20'h00000;
			rdrq_packet_w2e_esto_w = 20'h00000;
		end
		rdrq_packet_e2w_wsto_w = rdrq_packet_e2w_esti_muxed;
	end
	always @(*) begin
		if (rdrs_packet_bank2ring[0] == 1'h1)
			rdrs_packet_w2e_esto_w = rdrs_packet_bank2ring;
		else if (rdrs_packet_w2e_wsti_muxed[0] & cfg_ld_dma_on)
			rdrs_packet_w2e_esto_w = 65'h00000000000000000;
		else
			rdrs_packet_w2e_esto_w = rdrs_packet_w2e_wsti_muxed;
		if (rdrs_packet_w2e_wsti_muxed[0] & cfg_ld_dma_on)
			rdrs_packet_ring2dma_w = rdrs_packet_w2e_wsti_muxed;
		else
			rdrs_packet_ring2dma_w = 65'h00000000000000000;
		rdrs_packet_e2w_wsto_w = rdrs_packet_e2w_esti_muxed;
	end
	always @(posedge clk or posedge reset)
		if (reset) begin
			wr_packet_w2e_esto <= 92'h00000000000000000000000;
			wr_packet_e2w_wsto <= 92'h00000000000000000000000;
			wr_packet_ring2bank <= 92'h00000000000000000000000;
			rdrq_packet_w2e_esto <= 20'h00000;
			rdrq_packet_e2w_wsto <= 20'h00000;
			rdrq_packet_ring2bank <= 20'h00000;
			rdrs_packet_w2e_esto <= 65'h00000000000000000;
			rdrs_packet_e2w_wsto <= 65'h00000000000000000;
		end
		else begin
			wr_packet_w2e_esto <= wr_packet_w2e_esto_w;
			wr_packet_e2w_wsto <= wr_packet_e2w_wsto_w;
			wr_packet_ring2bank <= wr_packet_ring2bank_w;
			rdrq_packet_w2e_esto <= rdrq_packet_w2e_esto_w;
			rdrq_packet_e2w_wsto <= rdrq_packet_e2w_wsto_w;
			rdrq_packet_ring2bank <= rdrq_packet_ring2bank_w;
			rdrs_packet_w2e_esto <= rdrs_packet_w2e_esto_w;
			rdrs_packet_e2w_wsto <= rdrs_packet_e2w_wsto_w;
		end
	always @(*) rdrs_packet_ring2dma = rdrs_packet_ring2dma_w;
	assign clk_en_ring2bank = ring2bank_wr_clk_en | ring2bank_rd_clk_en;
	glb_clk_en_gen_4 #(.cnt(32'h00000004)) ring2bank_wr_clk_en_gen(
		.clk(clk),
		.enable(wr_packet_ring2bank_w[91]),
		.reset(reset),
		.clk_en(ring2bank_wr_clk_en)
	);
	glb_clk_en_gen_6 #(.cnt(32'h00000006)) ring2bank_rd_clk_en_gen(
		.clk(clk),
		.enable(rdrq_packet_ring2bank_w[19]),
		.reset(reset),
		.clk_en(ring2bank_rd_clk_en)
	);
endmodule
module glb_sched_gen (
	clk,
	clk_en,
	current_addr,
	cycle_count,
	finished,
	reset,
	restart,
	valid_output
);
	input wire clk;
	input wire clk_en;
	input wire [15:0] current_addr;
	input wire [15:0] cycle_count;
	input wire finished;
	input wire reset;
	input wire restart;
	output reg valid_output;
	reg valid_gate;
	always @(posedge clk or posedge reset)
		if (reset)
			valid_gate <= 1'h1;
		else if (clk_en) begin
			if (restart)
				valid_gate <= 1'h0;
			else if (finished)
				valid_gate <= 1'h1;
		end
	always @(*) valid_output = (cycle_count == current_addr) & ~valid_gate;
endmodule
module glb_store_dma (
	cfg_data_network_f2g_mux,
	cfg_data_network_latency,
	cfg_st_dma_ctrl_mode,
	cfg_st_dma_ctrl_valid_mode,
	cfg_st_dma_header,
	cfg_st_dma_num_blocks,
	cfg_st_dma_num_repeat,
	cfg_tile_connected_next,
	cfg_tile_connected_prev,
	clk,
	ctrl_f2g,
	data_f2g,
	data_f2g_vld,
	reset,
	st_dma_start_pulse,
	clk_en_dma2bank,
	data_f2g_rdy,
	st_dma_done_interrupt,
	wr_packet_dma2bank,
	wr_packet_dma2ring
);
	input wire [1:0] cfg_data_network_f2g_mux;
	input wire [5:0] cfg_data_network_latency;
	input wire [1:0] cfg_st_dma_ctrl_mode;
	input wire [1:0] cfg_st_dma_ctrl_valid_mode;
	input wire [514:0] cfg_st_dma_header;
	input wire [31:0] cfg_st_dma_num_blocks;
	input wire cfg_st_dma_num_repeat;
	input wire cfg_tile_connected_next;
	input wire cfg_tile_connected_prev;
	input wire clk;
	input wire [1:0] ctrl_f2g;
	input wire [31:0] data_f2g;
	input wire [1:0] data_f2g_vld;
	input wire reset;
	input wire st_dma_start_pulse;
	output wire clk_en_dma2bank;
	output reg [1:0] data_f2g_rdy;
	output reg st_dma_done_interrupt;
	output reg [91:0] wr_packet_dma2bank;
	output reg [91:0] wr_packet_dma2ring;
	reg bank_addr_match;
	reg [18:0] bank_wr_addr;
	reg [63:0] bank_wr_data_cache_r;
	reg [63:0] bank_wr_data_cache_w;
	reg bank_wr_en;
	reg [7:0] bank_wr_strb_cache_r;
	reg [7:0] bank_wr_strb_cache_w;
	reg block_done;
	reg [1:0] ctrl_f2g_r;
	wire [514:0] current_dma_header;
	reg [15:0] cycle_count;
	wire cycle_counter_en;
	wire [15:0] cycle_current_addr;
	wire [111:0] cycle_stride_addr_gen_strides;
	wire cycle_valid;
	wire [15:0] data_cgra2fifo;
	wire [19:0] data_current_addr;
	reg [31:0] data_f2g_r;
	reg [1:0] data_f2g_vld_r;
	wire [15:0] data_fifo2dma;
	reg data_ready_g2f_w;
	wire [19:0] data_stride_addr_gen_start_addr;
	wire [139:0] data_stride_addr_gen_strides;
	wire dma2bank_clk_en;
	wire [19:0] done_pulse_d_arr;
	reg done_pulse_w;
	wire fifo2cgra_ready;
	wire fifo_almost_full;
	wire fifo_empty;
	wire fifo_full;
	wire fifo_pop;
	wire fifo_pop_ready;
	wire fifo_push;
	reg is_first;
	reg is_last;
	reg is_last_block;
	reg iter_step_valid;
	reg [18:0] last_strm_wr_addr_r;
	wire loop_done;
	reg loop_done_muxed;
	wire [223:0] loop_iter_ranges;
	wire [2:0] loop_mux_sel;
	reg repeat_cnt;
	reg rv_is_metadata;
	wire rv_mode_on;
	reg [31:0] rv_num_blocks_cnt;
	reg [15:0] rv_num_data_cnt;
	wire st_dma_done_pulse;
	wire st_dma_done_pulse_last;
	reg st_dma_start_pulse_next;
	reg st_dma_start_pulse_r;
	reg [15:0] strm_data;
	reg [1:0] strm_data_sel;
	reg strm_data_valid;
	reg strm_run;
	reg [18:0] strm_wr_addr_w;
	reg [15:0] strm_wr_data_w;
	reg strm_wr_en_w;
	reg [91:0] wr_packet_dma2bank_w;
	reg [91:0] wr_packet_dma2ring_w;
	assign current_dma_header = cfg_st_dma_header;
	always @(posedge clk or posedge reset)
		if (reset)
			repeat_cnt <= 1'h0;
		else if (cfg_st_dma_ctrl_mode == 2'h2) begin
			if (st_dma_done_pulse) begin
				if ((repeat_cnt + 1'h1) < cfg_st_dma_num_repeat)
					repeat_cnt <= repeat_cnt + 1'h1;
			end
		end
		else if (cfg_st_dma_ctrl_mode == 2'h3) begin
			if (st_dma_done_pulse) begin
				if (((repeat_cnt + 1'h1) < cfg_st_dma_num_repeat) & ((repeat_cnt + 1'h1) < 1'h1))
					repeat_cnt <= repeat_cnt + 1'h1;
			end
		end
	always @(posedge clk or posedge reset)
		if (reset)
			is_first <= 1'h0;
		else if (st_dma_start_pulse_r)
			is_first <= 1'h1;
		else if (strm_wr_en_w)
			is_first <= 1'h0;
	always @(posedge clk or posedge reset)
		if (reset)
			is_last <= 1'h0;
		else if (loop_done_muxed)
			is_last <= 1'h1;
		else if (bank_wr_en)
			is_last <= 1'h0;
	always @(posedge clk or posedge reset)
		if (reset)
			strm_run <= 1'h0;
		else if (st_dma_start_pulse_r)
			strm_run <= 1'h1;
		else if (loop_done_muxed)
			strm_run <= 1'h0;
	always @(*)
		if (cfg_st_dma_ctrl_mode == 2'h0)
			st_dma_start_pulse_next = 1'h0;
		else if (cfg_st_dma_ctrl_mode == 2'h1)
			st_dma_start_pulse_next = ~strm_run & st_dma_start_pulse;
		else if ((cfg_st_dma_ctrl_mode == 2'h2) | (cfg_st_dma_ctrl_mode == 2'h3))
			st_dma_start_pulse_next = (~strm_run & st_dma_start_pulse) | (st_dma_done_pulse & ((repeat_cnt + 1'h1) < cfg_st_dma_num_repeat));
		else
			st_dma_start_pulse_next = 1'h0;
	always @(posedge clk or posedge reset)
		if (reset)
			st_dma_start_pulse_r <= 1'h0;
		else if (st_dma_start_pulse_r)
			st_dma_start_pulse_r <= 1'h0;
		else
			st_dma_start_pulse_r <= st_dma_start_pulse_next;
	always @(posedge clk or posedge reset)
		if (reset)
			cycle_count <= 16'h0000;
		else if (st_dma_start_pulse_r)
			cycle_count <= 16'h0000;
		else if (loop_done_muxed)
			cycle_count <= 16'h0000;
		else if (cycle_counter_en & strm_run)
			cycle_count <= cycle_count + 16'h0001;
	always @(posedge clk or posedge reset)
		if (reset) begin
			data_f2g_r <= 32'h00000000;
			data_f2g_vld_r <= 2'h0;
			ctrl_f2g_r <= 2'h0;
		end
		else begin
			data_f2g_r[0+:16] <= data_f2g[0+:16];
			data_f2g_r[16+:16] <= data_f2g[16+:16];
			data_f2g_vld_r <= data_f2g_vld;
			ctrl_f2g_r <= ctrl_f2g;
		end
	always @(*) begin
		strm_data = 16'h0000;
		strm_data_valid = 1'h0;
		if (cfg_data_network_f2g_mux[0] == 1'h1) begin
			strm_data = data_f2g_r[0+:16];
			data_f2g_rdy[0] = data_ready_g2f_w;
			if (rv_mode_on)
				strm_data_valid = data_f2g_vld_r[0];
			else
				strm_data_valid = ctrl_f2g_r[0];
		end
		else begin
			strm_data = strm_data;
			strm_data_valid = strm_data_valid;
			data_f2g_rdy[0] = 1'h0;
		end
		if (cfg_data_network_f2g_mux[1] == 1'h1) begin
			strm_data = data_f2g_r[16+:16];
			data_f2g_rdy[1] = data_ready_g2f_w;
			if (rv_mode_on)
				strm_data_valid = data_f2g_vld_r[1];
			else
				strm_data_valid = ctrl_f2g_r[1];
		end
		else begin
			strm_data = strm_data;
			strm_data_valid = strm_data_valid;
			data_f2g_rdy[1] = 1'h0;
		end
	end
	always @(*)
		if (cycle_counter_en)
			iter_step_valid = cycle_valid;
		else if (rv_mode_on)
			iter_step_valid = strm_run & fifo_pop_ready;
		else
			iter_step_valid = strm_data_valid;
	function automatic [18:0] sv2v_cast_19;
		input reg [18:0] inp;
		sv2v_cast_19 = inp;
	endfunction
	always @(*) begin
		strm_wr_en_w = iter_step_valid;
		if (rv_mode_on) begin
			strm_wr_addr_w = sv2v_cast_19(data_current_addr);
			strm_wr_data_w = data_fifo2dma;
		end
		else begin
			strm_wr_addr_w = sv2v_cast_19(data_current_addr);
			strm_wr_data_w = strm_data;
		end
	end
	always @(posedge clk or posedge reset)
		if (reset)
			last_strm_wr_addr_r <= 19'h00000;
		else if (strm_wr_en_w)
			last_strm_wr_addr_r <= strm_wr_addr_w;
	always @(*) strm_data_sel = strm_wr_addr_w[2:1];
	always @(*) begin
		bank_wr_strb_cache_w = bank_wr_strb_cache_r;
		bank_wr_data_cache_w = bank_wr_data_cache_r;
		if (bank_wr_en) begin
			bank_wr_strb_cache_w = 8'h00;
			bank_wr_data_cache_w = 64'h0000000000000000;
		end
		if (strm_wr_en_w) begin
			if (strm_data_sel == 2'h0) begin
				bank_wr_strb_cache_w[1:0] = 2'h3;
				bank_wr_data_cache_w[15:0] = strm_wr_data_w;
			end
			else if (strm_data_sel == 2'h1) begin
				bank_wr_strb_cache_w[3:2] = 2'h3;
				bank_wr_data_cache_w[31:16] = strm_wr_data_w;
			end
			else if (strm_data_sel == 2'h2) begin
				bank_wr_strb_cache_w[5:4] = 2'h3;
				bank_wr_data_cache_w[47:32] = strm_wr_data_w;
			end
			else if (strm_data_sel == 2'h3) begin
				bank_wr_strb_cache_w[7:6] = 2'h3;
				bank_wr_data_cache_w[63:48] = strm_wr_data_w;
			end
			else begin
				bank_wr_strb_cache_w = bank_wr_strb_cache_r;
				bank_wr_data_cache_w = bank_wr_data_cache_r;
			end
		end
	end
	always @(posedge clk or posedge reset)
		if (reset) begin
			bank_wr_strb_cache_r <= 8'h00;
			bank_wr_data_cache_r <= 64'h0000000000000000;
		end
		else begin
			bank_wr_strb_cache_r <= bank_wr_strb_cache_w;
			bank_wr_data_cache_r <= bank_wr_data_cache_w;
		end
	always @(*) begin
		bank_addr_match = strm_wr_addr_w[18:3] == last_strm_wr_addr_r[18:3];
		bank_wr_en = ((strm_wr_en_w & ~bank_addr_match) & ~is_first) | is_last;
		bank_wr_addr = last_strm_wr_addr_r;
	end
	always @(posedge clk or posedge reset)
		if (reset) begin
			wr_packet_dma2bank <= 92'h00000000000000000000000;
			wr_packet_dma2ring <= 92'h00000000000000000000000;
		end
		else begin
			wr_packet_dma2bank <= wr_packet_dma2bank_w;
			wr_packet_dma2ring <= wr_packet_dma2ring_w;
		end
	always @(*)
		if (cfg_tile_connected_next | cfg_tile_connected_prev) begin
			wr_packet_dma2bank_w = 92'h00000000000000000000000;
			wr_packet_dma2ring_w[91] = bank_wr_en;
			wr_packet_dma2ring_w[90-:8] = bank_wr_strb_cache_r;
			wr_packet_dma2ring_w[63-:64] = bank_wr_data_cache_r;
			wr_packet_dma2ring_w[82-:19] = bank_wr_addr;
		end
		else begin
			wr_packet_dma2bank_w[91] = bank_wr_en;
			wr_packet_dma2bank_w[90-:8] = bank_wr_strb_cache_r;
			wr_packet_dma2bank_w[63-:64] = bank_wr_data_cache_r;
			wr_packet_dma2bank_w[82-:19] = bank_wr_addr;
			wr_packet_dma2ring_w = 92'h00000000000000000000000;
		end
	assign clk_en_dma2bank = dma2bank_clk_en;
	always @(*) done_pulse_w = loop_done_muxed & strm_run;
	function automatic [4:0] sv2v_cast_5;
		input reg [4:0] inp;
		sv2v_cast_5 = inp;
	endfunction
	assign st_dma_done_pulse = done_pulse_d_arr[sv2v_cast_5(cfg_data_network_latency) + 5'h01];
	always @(posedge clk or posedge reset)
		if (reset)
			st_dma_done_interrupt <= 1'h0;
		else if (st_dma_done_pulse)
			st_dma_done_interrupt <= 1'h1;
		else if (st_dma_done_pulse_last)
			st_dma_done_interrupt <= 1'h0;
	always @(*)
		if (rv_mode_on)
			block_done = (strm_run & ~rv_is_metadata) & (((rv_num_data_cnt == 16'h0001) & fifo_pop_ready) | (rv_num_data_cnt == 16'h0000));
		else
			block_done = 1'h0;
	always @(*)
		if (rv_mode_on)
			loop_done_muxed = block_done & is_last_block;
		else
			loop_done_muxed = loop_done;
	always @(posedge clk or posedge reset)
		if (reset)
			rv_num_blocks_cnt <= 32'h00000000;
		else if (rv_mode_on) begin
			if (st_dma_start_pulse_r)
				rv_num_blocks_cnt <= cfg_st_dma_num_blocks;
			else if (block_done & (rv_num_blocks_cnt > 32'h00000000))
				rv_num_blocks_cnt <= rv_num_blocks_cnt - 32'h00000001;
		end
	always @(*) is_last_block = rv_num_blocks_cnt == 32'h00000001;
	always @(posedge clk or posedge reset)
		if (reset)
			rv_is_metadata <= 1'h0;
		else if (rv_mode_on) begin
			if (st_dma_start_pulse_r)
				rv_is_metadata <= 1'h1;
			else if ((rv_mode_on & block_done) & ~is_last_block)
				rv_is_metadata <= 1'h1;
			else if (rv_is_metadata & fifo_pop_ready)
				rv_is_metadata <= 1'h0;
		end
	always @(posedge clk or posedge reset)
		if (reset)
			rv_num_data_cnt <= 16'h0000;
		else if (st_dma_start_pulse_r)
			rv_num_data_cnt <= 16'h0000;
		else if ((strm_run & rv_is_metadata) & fifo_pop_ready)
			rv_num_data_cnt <= data_fifo2dma;
		else if ((rv_num_data_cnt > 16'h0000) & fifo_pop_ready)
			rv_num_data_cnt <= rv_num_data_cnt - 16'h0001;
	always @(*)
		if (rv_mode_on)
			data_ready_g2f_w = fifo2cgra_ready;
		else
			data_ready_g2f_w = 1'h0;
	assign rv_mode_on = cfg_st_dma_ctrl_valid_mode == 2'h1;
	assign data_cgra2fifo = strm_data;
	assign fifo_pop_ready = ~fifo_empty;
	assign fifo_pop = ~fifo_empty & strm_run;
	assign fifo_push = ~fifo_full & strm_data_valid;
	assign fifo2cgra_ready = ~fifo_almost_full;
	assign loop_iter_ranges[0+:32] = current_dma_header[475-:32];
	assign loop_iter_ranges[32+:32] = current_dma_header[407-:32];
	assign loop_iter_ranges[64+:32] = current_dma_header[339-:32];
	assign loop_iter_ranges[96+:32] = current_dma_header[271-:32];
	assign loop_iter_ranges[128+:32] = current_dma_header[203-:32];
	assign loop_iter_ranges[160+:32] = current_dma_header[135-:32];
	assign loop_iter_ranges[192+:32] = current_dma_header[67-:32];
	assign cycle_counter_en = cfg_st_dma_ctrl_valid_mode == 2'h2;
	assign cycle_stride_addr_gen_strides[0+:16] = current_dma_header[423-:16];
	assign cycle_stride_addr_gen_strides[16+:16] = current_dma_header[355-:16];
	assign cycle_stride_addr_gen_strides[32+:16] = current_dma_header[287-:16];
	assign cycle_stride_addr_gen_strides[48+:16] = current_dma_header[219-:16];
	assign cycle_stride_addr_gen_strides[64+:16] = current_dma_header[151-:16];
	assign cycle_stride_addr_gen_strides[80+:16] = current_dma_header[83-:16];
	assign cycle_stride_addr_gen_strides[96+:16] = current_dma_header[15-:16];
	function automatic [19:0] sv2v_cast_20;
		input reg [19:0] inp;
		sv2v_cast_20 = inp;
	endfunction
	assign data_stride_addr_gen_start_addr = sv2v_cast_20(current_dma_header[514-:19]);
	assign data_stride_addr_gen_strides[0+:20] = current_dma_header[443-:20];
	assign data_stride_addr_gen_strides[20+:20] = current_dma_header[375-:20];
	assign data_stride_addr_gen_strides[40+:20] = current_dma_header[307-:20];
	assign data_stride_addr_gen_strides[60+:20] = current_dma_header[239-:20];
	assign data_stride_addr_gen_strides[80+:20] = current_dma_header[171-:20];
	assign data_stride_addr_gen_strides[100+:20] = current_dma_header[103-:20];
	assign data_stride_addr_gen_strides[120+:20] = current_dma_header[35-:20];
	glb_clk_en_gen_4 #(.cnt(32'h00000004)) dma2bank_clk_en_gen(
		.clk(clk),
		.enable(wr_packet_dma2bank_w[91]),
		.reset(reset),
		.clk_en(dma2bank_clk_en)
	);
	pipeline_w_1_d_20_array done_pulse_pipeline(
		.clk(clk),
		.clk_en(1'h1),
		.in_(done_pulse_w),
		.reset(reset),
		.out_(done_pulse_d_arr)
	);
	pipeline_w_1_d_5 st_dma_interrupt_pipeline(
		.clk(clk),
		.clk_en(1'h1),
		.in_(st_dma_done_pulse),
		.reset(reset),
		.out_(st_dma_done_pulse_last)
	);
	reg_fifo_d_4_w_16 #(.data_width(16'h0010)) data_f2g_fifo(
		.almost_empty_diff(2'h2),
		.almost_full_diff(2'h2),
		.clk(clk),
		.clk_en(rv_mode_on),
		.data_in(data_cgra2fifo),
		.flush(st_dma_start_pulse_r),
		.pop(fifo_pop),
		.push(fifo_push),
		.reset(reset),
		.almost_full(fifo_almost_full),
		.data_out(data_fifo2dma),
		.empty(fifo_empty),
		.full(fifo_full)
	);
	glb_loop_iter_7 loop_iter(
		.clk(clk),
		.clk_en(1'h1),
		.dim(current_dma_header[479-:4]),
		.ranges(loop_iter_ranges),
		.reset(reset),
		.step(iter_step_valid),
		.mux_sel_out(loop_mux_sel),
		.restart(loop_done)
	);
	glb_sched_gen cycle_stride_sched_gen(
		.clk(clk),
		.clk_en(cycle_counter_en),
		.current_addr(cycle_current_addr),
		.cycle_count(cycle_count),
		.finished(loop_done_muxed),
		.reset(reset),
		.restart(st_dma_start_pulse_r),
		.valid_output(cycle_valid)
	);
	glb_addr_gen_7 #(
		.addr_width(32'h00000010),
		.loop_level(32'h00000007)
	) cycle_stride_addr_gen(
		.clk(clk),
		.clk_en(cycle_counter_en),
		.mux_sel(loop_mux_sel),
		.reset(reset),
		.restart(st_dma_start_pulse_r),
		.start_addr(current_dma_header[495-:16]),
		.step(iter_step_valid),
		.strides(cycle_stride_addr_gen_strides),
		.addr_out(cycle_current_addr)
	);
	glb_addr_gen_7 #(
		.addr_width(32'h00000014),
		.loop_level(32'h00000007)
	) data_stride_addr_gen(
		.clk(clk),
		.clk_en(1'h1),
		.mux_sel(loop_mux_sel),
		.reset(reset),
		.restart(st_dma_start_pulse_r),
		.start_addr(data_stride_addr_gen_start_addr),
		.step(iter_step_valid),
		.strides(data_stride_addr_gen_strides),
		.addr_out(data_current_addr)
	);
endmodule
module glb_tile (
	cfg_pcfg_tile_connected_wsti,
	cfg_tile_connected_wsti,
	cgra_cfg_jtag_addr_bypass_wsti,
	cgra_cfg_jtag_addr_wsti,
	cgra_cfg_jtag_data_wsti,
	cgra_cfg_jtag_rd_en_bypass_wsti,
	cgra_cfg_jtag_rd_en_wsti,
	cgra_cfg_jtag_wr_en_wsti,
	cgra_cfg_pcfg_addr_e2w_esti,
	cgra_cfg_pcfg_addr_w2e_wsti,
	cgra_cfg_pcfg_data_e2w_esti,
	cgra_cfg_pcfg_data_w2e_wsti,
	cgra_cfg_pcfg_rd_en_e2w_esti,
	cgra_cfg_pcfg_rd_en_w2e_wsti,
	cgra_cfg_pcfg_wr_en_e2w_esti,
	cgra_cfg_pcfg_wr_en_w2e_wsti,
	clk,
	clk_en_bank_master,
	clk_en_master,
	clk_en_pcfg_broadcast,
	glb_tile_id,
	if_cfg_est_m_rd_data,
	if_cfg_est_m_rd_data_valid,
	if_cfg_wst_s_rd_addr,
	if_cfg_wst_s_rd_clk_en,
	if_cfg_wst_s_rd_en,
	if_cfg_wst_s_wr_addr,
	if_cfg_wst_s_wr_clk_en,
	if_cfg_wst_s_wr_data,
	if_cfg_wst_s_wr_en,
	if_proc_est_m_rd_data,
	if_proc_est_m_rd_data_valid,
	if_proc_wst_s_rd_addr,
	if_proc_wst_s_rd_clk_en,
	if_proc_wst_s_rd_en,
	if_proc_wst_s_wr_addr,
	if_proc_wst_s_wr_clk_en,
	if_proc_wst_s_wr_data,
	if_proc_wst_s_wr_en,
	if_proc_wst_s_wr_strb,
	pcfg_rd_addr_e2w_esti,
	pcfg_rd_addr_w2e_wsti,
	pcfg_rd_data_e2w_esti,
	pcfg_rd_data_valid_e2w_esti,
	pcfg_rd_data_valid_w2e_wsti,
	pcfg_rd_data_w2e_wsti,
	pcfg_rd_en_e2w_esti,
	pcfg_rd_en_w2e_wsti,
	pcfg_start_pulse,
	reset,
	strm_ctrl_f2g,
	strm_data_f2g,
	strm_data_f2g_vld,
	strm_data_g2f_rdy,
	strm_f2g_start_pulse,
	strm_g2f_start_pulse,
	strm_rd_addr_e2w_esti,
	strm_rd_addr_w2e_wsti,
	strm_rd_data_e2w_esti,
	strm_rd_data_valid_e2w_esti,
	strm_rd_data_valid_w2e_wsti,
	strm_rd_data_w2e_wsti,
	strm_rd_en_e2w_esti,
	strm_rd_en_w2e_wsti,
	strm_wr_addr_e2w_esti,
	strm_wr_addr_w2e_wsti,
	strm_wr_data_e2w_esti,
	strm_wr_data_w2e_wsti,
	strm_wr_en_e2w_esti,
	strm_wr_en_w2e_wsti,
	strm_wr_strb_e2w_esti,
	strm_wr_strb_w2e_wsti,
	cfg_pcfg_tile_connected_esto,
	cfg_tile_connected_esto,
	cgra_cfg_g2f_cfg_addr,
	cgra_cfg_g2f_cfg_data,
	cgra_cfg_g2f_cfg_rd_en,
	cgra_cfg_g2f_cfg_wr_en,
	cgra_cfg_jtag_addr_bypass_esto,
	cgra_cfg_jtag_addr_esto,
	cgra_cfg_jtag_data_esto,
	cgra_cfg_jtag_rd_en_bypass_esto,
	cgra_cfg_jtag_rd_en_esto,
	cgra_cfg_jtag_wr_en_esto,
	cgra_cfg_pcfg_addr_e2w_wsto,
	cgra_cfg_pcfg_addr_w2e_esto,
	cgra_cfg_pcfg_data_e2w_wsto,
	cgra_cfg_pcfg_data_w2e_esto,
	cgra_cfg_pcfg_rd_en_e2w_wsto,
	cgra_cfg_pcfg_rd_en_w2e_esto,
	cgra_cfg_pcfg_wr_en_e2w_wsto,
	cgra_cfg_pcfg_wr_en_w2e_esto,
	data_flush,
	if_cfg_est_m_rd_addr,
	if_cfg_est_m_rd_clk_en,
	if_cfg_est_m_rd_en,
	if_cfg_est_m_wr_addr,
	if_cfg_est_m_wr_clk_en,
	if_cfg_est_m_wr_data,
	if_cfg_est_m_wr_en,
	if_cfg_wst_s_rd_data,
	if_cfg_wst_s_rd_data_valid,
	if_proc_est_m_rd_addr,
	if_proc_est_m_rd_clk_en,
	if_proc_est_m_rd_en,
	if_proc_est_m_wr_addr,
	if_proc_est_m_wr_clk_en,
	if_proc_est_m_wr_data,
	if_proc_est_m_wr_en,
	if_proc_est_m_wr_strb,
	if_proc_wst_s_rd_data,
	if_proc_wst_s_rd_data_valid,
	pcfg_g2f_interrupt_pulse,
	pcfg_rd_addr_e2w_wsto,
	pcfg_rd_addr_w2e_esto,
	pcfg_rd_data_e2w_wsto,
	pcfg_rd_data_valid_e2w_wsto,
	pcfg_rd_data_valid_w2e_esto,
	pcfg_rd_data_w2e_esto,
	pcfg_rd_en_e2w_wsto,
	pcfg_rd_en_w2e_esto,
	strm_ctrl_g2f,
	strm_data_f2g_rdy,
	strm_data_g2f,
	strm_data_g2f_vld,
	strm_f2g_interrupt_pulse,
	strm_g2f_interrupt_pulse,
	strm_rd_addr_e2w_wsto,
	strm_rd_addr_w2e_esto,
	strm_rd_data_e2w_wsto,
	strm_rd_data_valid_e2w_wsto,
	strm_rd_data_valid_w2e_esto,
	strm_rd_data_w2e_esto,
	strm_rd_en_e2w_wsto,
	strm_rd_en_w2e_esto,
	strm_wr_addr_e2w_wsto,
	strm_wr_addr_w2e_esto,
	strm_wr_data_e2w_wsto,
	strm_wr_data_w2e_esto,
	strm_wr_en_e2w_wsto,
	strm_wr_en_w2e_esto,
	strm_wr_strb_e2w_wsto,
	strm_wr_strb_w2e_esto
);
	input wire cfg_pcfg_tile_connected_wsti;
	input wire cfg_tile_connected_wsti;
	input wire [31:0] cgra_cfg_jtag_addr_bypass_wsti;
	input wire [31:0] cgra_cfg_jtag_addr_wsti;
	input wire [31:0] cgra_cfg_jtag_data_wsti;
	input wire cgra_cfg_jtag_rd_en_bypass_wsti;
	input wire cgra_cfg_jtag_rd_en_wsti;
	input wire cgra_cfg_jtag_wr_en_wsti;
	input wire [31:0] cgra_cfg_pcfg_addr_e2w_esti;
	input wire [31:0] cgra_cfg_pcfg_addr_w2e_wsti;
	input wire [31:0] cgra_cfg_pcfg_data_e2w_esti;
	input wire [31:0] cgra_cfg_pcfg_data_w2e_wsti;
	input wire cgra_cfg_pcfg_rd_en_e2w_esti;
	input wire cgra_cfg_pcfg_rd_en_w2e_wsti;
	input wire cgra_cfg_pcfg_wr_en_e2w_esti;
	input wire cgra_cfg_pcfg_wr_en_w2e_wsti;
	input wire clk;
	input wire clk_en_bank_master;
	input wire clk_en_master;
	input wire clk_en_pcfg_broadcast;
	input wire glb_tile_id;
	input wire [31:0] if_cfg_est_m_rd_data;
	input wire if_cfg_est_m_rd_data_valid;
	input wire [11:0] if_cfg_wst_s_rd_addr;
	input wire if_cfg_wst_s_rd_clk_en;
	input wire if_cfg_wst_s_rd_en;
	input wire [11:0] if_cfg_wst_s_wr_addr;
	input wire if_cfg_wst_s_wr_clk_en;
	input wire [31:0] if_cfg_wst_s_wr_data;
	input wire if_cfg_wst_s_wr_en;
	input wire [63:0] if_proc_est_m_rd_data;
	input wire if_proc_est_m_rd_data_valid;
	input wire [18:0] if_proc_wst_s_rd_addr;
	input wire if_proc_wst_s_rd_clk_en;
	input wire if_proc_wst_s_rd_en;
	input wire [18:0] if_proc_wst_s_wr_addr;
	input wire if_proc_wst_s_wr_clk_en;
	input wire [63:0] if_proc_wst_s_wr_data;
	input wire if_proc_wst_s_wr_en;
	input wire [7:0] if_proc_wst_s_wr_strb;
	input wire [18:0] pcfg_rd_addr_e2w_esti;
	input wire [18:0] pcfg_rd_addr_w2e_wsti;
	input wire [63:0] pcfg_rd_data_e2w_esti;
	input wire pcfg_rd_data_valid_e2w_esti;
	input wire pcfg_rd_data_valid_w2e_wsti;
	input wire [63:0] pcfg_rd_data_w2e_wsti;
	input wire pcfg_rd_en_e2w_esti;
	input wire pcfg_rd_en_w2e_wsti;
	input wire pcfg_start_pulse;
	input wire reset;
	input wire [1:0] strm_ctrl_f2g;
	input wire [31:0] strm_data_f2g;
	input wire [1:0] strm_data_f2g_vld;
	input wire [1:0] strm_data_g2f_rdy;
	input wire strm_f2g_start_pulse;
	input wire strm_g2f_start_pulse;
	input wire [18:0] strm_rd_addr_e2w_esti;
	input wire [18:0] strm_rd_addr_w2e_wsti;
	input wire [63:0] strm_rd_data_e2w_esti;
	input wire strm_rd_data_valid_e2w_esti;
	input wire strm_rd_data_valid_w2e_wsti;
	input wire [63:0] strm_rd_data_w2e_wsti;
	input wire strm_rd_en_e2w_esti;
	input wire strm_rd_en_w2e_wsti;
	input wire [18:0] strm_wr_addr_e2w_esti;
	input wire [18:0] strm_wr_addr_w2e_wsti;
	input wire [63:0] strm_wr_data_e2w_esti;
	input wire [63:0] strm_wr_data_w2e_wsti;
	input wire strm_wr_en_e2w_esti;
	input wire strm_wr_en_w2e_wsti;
	input wire [7:0] strm_wr_strb_e2w_esti;
	input wire [7:0] strm_wr_strb_w2e_wsti;
	output wire cfg_pcfg_tile_connected_esto;
	output wire cfg_tile_connected_esto;
	output wire [63:0] cgra_cfg_g2f_cfg_addr;
	output wire [63:0] cgra_cfg_g2f_cfg_data;
	output wire [1:0] cgra_cfg_g2f_cfg_rd_en;
	output wire [1:0] cgra_cfg_g2f_cfg_wr_en;
	output wire [31:0] cgra_cfg_jtag_addr_bypass_esto;
	output wire [31:0] cgra_cfg_jtag_addr_esto;
	output wire [31:0] cgra_cfg_jtag_data_esto;
	output wire cgra_cfg_jtag_rd_en_bypass_esto;
	output wire cgra_cfg_jtag_rd_en_esto;
	output wire cgra_cfg_jtag_wr_en_esto;
	output wire [31:0] cgra_cfg_pcfg_addr_e2w_wsto;
	output wire [31:0] cgra_cfg_pcfg_addr_w2e_esto;
	output wire [31:0] cgra_cfg_pcfg_data_e2w_wsto;
	output wire [31:0] cgra_cfg_pcfg_data_w2e_esto;
	output wire cgra_cfg_pcfg_rd_en_e2w_wsto;
	output wire cgra_cfg_pcfg_rd_en_w2e_esto;
	output wire cgra_cfg_pcfg_wr_en_e2w_wsto;
	output wire cgra_cfg_pcfg_wr_en_w2e_esto;
	output wire data_flush;
	output wire [11:0] if_cfg_est_m_rd_addr;
	output wire if_cfg_est_m_rd_clk_en;
	output wire if_cfg_est_m_rd_en;
	output wire [11:0] if_cfg_est_m_wr_addr;
	output wire if_cfg_est_m_wr_clk_en;
	output wire [31:0] if_cfg_est_m_wr_data;
	output wire if_cfg_est_m_wr_en;
	output wire [31:0] if_cfg_wst_s_rd_data;
	output wire if_cfg_wst_s_rd_data_valid;
	output wire [18:0] if_proc_est_m_rd_addr;
	output wire if_proc_est_m_rd_clk_en;
	output wire if_proc_est_m_rd_en;
	output wire [18:0] if_proc_est_m_wr_addr;
	output wire if_proc_est_m_wr_clk_en;
	output wire [63:0] if_proc_est_m_wr_data;
	output wire if_proc_est_m_wr_en;
	output wire [7:0] if_proc_est_m_wr_strb;
	output wire [63:0] if_proc_wst_s_rd_data;
	output wire if_proc_wst_s_rd_data_valid;
	output wire pcfg_g2f_interrupt_pulse;
	output wire [18:0] pcfg_rd_addr_e2w_wsto;
	output wire [18:0] pcfg_rd_addr_w2e_esto;
	output wire [63:0] pcfg_rd_data_e2w_wsto;
	output wire pcfg_rd_data_valid_e2w_wsto;
	output wire pcfg_rd_data_valid_w2e_esto;
	output wire [63:0] pcfg_rd_data_w2e_esto;
	output wire pcfg_rd_en_e2w_wsto;
	output wire pcfg_rd_en_w2e_esto;
	output wire [1:0] strm_ctrl_g2f;
	output wire [1:0] strm_data_f2g_rdy;
	output wire [31:0] strm_data_g2f;
	output wire [1:0] strm_data_g2f_vld;
	output wire strm_f2g_interrupt_pulse;
	output wire strm_g2f_interrupt_pulse;
	output wire [18:0] strm_rd_addr_e2w_wsto;
	output wire [18:0] strm_rd_addr_w2e_esto;
	output wire [63:0] strm_rd_data_e2w_wsto;
	output wire strm_rd_data_valid_e2w_wsto;
	output wire strm_rd_data_valid_w2e_esto;
	output wire [63:0] strm_rd_data_w2e_esto;
	output wire strm_rd_en_e2w_wsto;
	output wire strm_rd_en_w2e_esto;
	output wire [18:0] strm_wr_addr_e2w_wsto;
	output wire [18:0] strm_wr_addr_w2e_esto;
	output wire [63:0] strm_wr_data_e2w_wsto;
	output wire [63:0] strm_wr_data_w2e_esto;
	output wire strm_wr_en_e2w_wsto;
	output wire strm_wr_en_w2e_esto;
	output wire [7:0] strm_wr_strb_e2w_wsto;
	output wire [7:0] strm_wr_strb_w2e_esto;
	wire [7:0] cfg_ld_dma_ctrl;
	wire [582:0] cfg_ld_dma_header;
	wire [5:0] cfg_pcfg_broadcast_mux;
	wire [17:0] cfg_pcfg_dma_ctrl;
	wire [34:0] cfg_pcfg_dma_header;
	wire cfg_pcfg_tile_connected_next;
	wire cfg_pcfg_tile_connected_prev;
	wire [6:0] cfg_st_dma_ctrl;
	wire [514:0] cfg_st_dma_header;
	wire [31:0] cfg_st_dma_num_blocks;
	wire cfg_tile_connected_next;
	wire cfg_tile_connected_prev;
	wire [131:0] cgra_cfg_g2f_cfg_w;
	wire [65:0] cgra_cfg_pcfgdma2mux;
	wire clk_en_bank;
	wire clk_en_cfg;
	wire clk_en_ld_dma;
	wire clk_en_lddma2bank;
	wire clk_en_pcfg_dma;
	wire clk_en_pcfg_switch;
	wire clk_en_pcfgdma2bank;
	wire clk_en_pcfgring2bank;
	wire clk_en_proc_switch;
	wire clk_en_procsw2bank;
	wire clk_en_ring2bank;
	wire clk_en_st_dma;
	wire clk_en_stdma2bank;
	wire clk_en_strm_switch;
	wire gclk_bank;
	wire gclk_cfg;
	wire gclk_ld_dma;
	wire gclk_pcfg_broadcast;
	wire gclk_pcfg_dma;
	wire gclk_pcfg_switch;
	wire gclk_proc_switch;
	wire gclk_st_dma;
	wire gclk_strm_switch;
	wire [64:0] glb_bank_0_rdrs_packet;
	wire [64:0] glb_bank_1_rdrs_packet;
	wire [6:0] glb_cfg_cfg_data_network;
	wire [6:0] glb_cfg_cfg_pcfg_network;
	wire glb_clk_gate_bank_enable;
	wire glb_clk_gate_cfg_enable;
	wire glb_clk_gate_ld_dma_enable;
	wire glb_clk_gate_pcfg_broadcast_enable;
	wire glb_clk_gate_pcfg_dma_enable;
	wire glb_clk_gate_pcfg_switch_enable;
	wire glb_clk_gate_proc_switch_enable;
	wire glb_clk_gate_st_dma_enable;
	wire glb_clk_gate_strm_switch_enable;
	wire [65:0] glb_pcfg_broadcast_cgra_cfg_jtag_esto;
	wire [65:0] glb_pcfg_broadcast_cgra_cfg_jtag_wsti;
	wire [65:0] glb_pcfg_broadcast_cgra_cfg_pcfg_esti;
	wire [65:0] glb_pcfg_broadcast_cgra_cfg_pcfg_esto;
	wire [65:0] glb_pcfg_broadcast_cgra_cfg_pcfg_wsti;
	wire [65:0] glb_pcfg_broadcast_cgra_cfg_pcfg_wsto;
	wire glb_pcfg_ring_switch_cfg_ld_dma_on;
	wire glb_strm_ring_switch_cfg_ld_dma_on;
	wire [19:0] pcfg_rdrq_packet_e2w_esti;
	wire [19:0] pcfg_rdrq_packet_e2w_wsto;
	wire [19:0] pcfg_rdrq_packet_w2e_esto;
	wire [19:0] pcfg_rdrq_packet_w2e_wsti;
	wire [64:0] pcfg_rdrs_packet_e2w_esti;
	wire [64:0] pcfg_rdrs_packet_e2w_wsto;
	wire [64:0] pcfg_rdrs_packet_w2e_esto;
	wire [64:0] pcfg_rdrs_packet_w2e_wsti;
	wire [19:0] rdrq_packet_dma2bank;
	wire [19:0] rdrq_packet_dma2ring;
	wire [19:0] rdrq_packet_pcfgdma2bank;
	wire [19:0] rdrq_packet_pcfgdma2ring;
	wire [19:0] rdrq_packet_pcfgring2bank;
	wire [19:0] rdrq_packet_procsw2bank;
	wire [19:0] rdrq_packet_ring2bank;
	wire [35:0] rdrq_packet_sw2bankarr;
	wire [64:0] rdrs_packet_bank2dma;
	wire [64:0] rdrs_packet_bank2pcfgdma;
	wire [64:0] rdrs_packet_bank2pcfgring;
	wire [64:0] rdrs_packet_bank2procsw;
	wire [64:0] rdrs_packet_bank2ring;
	wire [129:0] rdrs_packet_bankarr2sw;
	wire [64:0] rdrs_packet_pcfgring2dma;
	wire [64:0] rdrs_packet_ring2dma;
	wire [19:0] strm_rdrq_packet_e2w_esti;
	wire [19:0] strm_rdrq_packet_e2w_wsto;
	wire [19:0] strm_rdrq_packet_w2e_esto;
	wire [19:0] strm_rdrq_packet_w2e_wsti;
	wire [64:0] strm_rdrs_packet_e2w_esti;
	wire [64:0] strm_rdrs_packet_e2w_wsto;
	wire [64:0] strm_rdrs_packet_w2e_esto;
	wire [64:0] strm_rdrs_packet_w2e_wsti;
	wire [91:0] strm_wr_packet_e2w_esti;
	wire [91:0] strm_wr_packet_e2w_wsto;
	wire [91:0] strm_wr_packet_w2e_esto;
	wire [91:0] strm_wr_packet_w2e_wsti;
	wire [91:0] wr_packet_dma2bank;
	wire [91:0] wr_packet_dma2ring;
	wire [91:0] wr_packet_procsw2bank;
	wire [91:0] wr_packet_ring2bank;
	wire [179:0] wr_packet_sw2bankarr;
	generate
		if (1) begin : if_cfg_est_m
			reg [11:0] rd_addr;
			reg rd_clk_en;
			wire [31:0] rd_data;
			wire rd_data_valid;
			reg rd_en;
			reg [11:0] wr_addr;
			reg wr_clk_en;
			reg [31:0] wr_data;
			reg wr_en;
		end
		if (1) begin : if_cfg_wst_s
			wire [11:0] rd_addr;
			wire rd_clk_en;
			reg [31:0] rd_data;
			reg rd_data_valid;
			wire rd_en;
			wire [11:0] wr_addr;
			wire wr_clk_en;
			wire [31:0] wr_data;
			wire wr_en;
		end
		if (1) begin : if_proc_est_m
			reg [18:0] rd_addr;
			reg rd_clk_en;
			wire [63:0] rd_data;
			wire rd_data_valid;
			reg rd_en;
			reg [18:0] wr_addr;
			reg wr_clk_en;
			reg [63:0] wr_data;
			reg wr_en;
			reg [7:0] wr_strb;
		end
		if (1) begin : if_proc_wst_s
			wire [18:0] rd_addr;
			wire rd_clk_en;
			reg [63:0] rd_data;
			reg rd_data_valid;
			wire rd_en;
			wire [18:0] wr_addr;
			wire wr_clk_en;
			wire [63:0] wr_data;
			wire wr_en;
			wire [7:0] wr_strb;
		end
	endgenerate
	assign if_proc_est_m_wr_en = if_proc_est_m.wr_en;
	assign if_proc_wst_s.wr_en = if_proc_wst_s_wr_en;
	assign if_proc_est_m_wr_addr = if_proc_est_m.wr_addr;
	assign if_proc_wst_s.wr_addr = if_proc_wst_s_wr_addr;
	assign if_proc_est_m_wr_data = if_proc_est_m.wr_data;
	assign if_proc_wst_s.wr_data = if_proc_wst_s_wr_data;
	assign if_proc_est_m_rd_en = if_proc_est_m.rd_en;
	assign if_proc_wst_s.rd_en = if_proc_wst_s_rd_en;
	assign if_proc_est_m_rd_addr = if_proc_est_m.rd_addr;
	assign if_proc_wst_s.rd_addr = if_proc_wst_s_rd_addr;
	assign if_proc_est_m_wr_strb = if_proc_est_m.wr_strb;
	assign if_proc_wst_s.wr_strb = if_proc_wst_s_wr_strb;
	assign if_proc_est_m_wr_clk_en = if_proc_est_m.wr_clk_en;
	assign if_proc_wst_s.wr_clk_en = if_proc_wst_s_wr_clk_en;
	assign if_proc_est_m_rd_clk_en = if_proc_est_m.rd_clk_en;
	assign if_proc_wst_s.rd_clk_en = if_proc_wst_s_rd_clk_en;
	assign if_proc_est_m.rd_data = if_proc_est_m_rd_data;
	assign if_proc_wst_s_rd_data = if_proc_wst_s.rd_data;
	assign if_proc_est_m.rd_data_valid = if_proc_est_m_rd_data_valid;
	assign if_proc_wst_s_rd_data_valid = if_proc_wst_s.rd_data_valid;
	assign if_cfg_est_m_wr_en = if_cfg_est_m.wr_en;
	assign if_cfg_wst_s.wr_en = if_cfg_wst_s_wr_en;
	assign if_cfg_est_m_wr_addr = if_cfg_est_m.wr_addr;
	assign if_cfg_wst_s.wr_addr = if_cfg_wst_s_wr_addr;
	assign if_cfg_est_m_wr_data = if_cfg_est_m.wr_data;
	assign if_cfg_wst_s.wr_data = if_cfg_wst_s_wr_data;
	assign if_cfg_est_m_rd_en = if_cfg_est_m.rd_en;
	assign if_cfg_wst_s.rd_en = if_cfg_wst_s_rd_en;
	assign if_cfg_est_m_rd_addr = if_cfg_est_m.rd_addr;
	assign if_cfg_wst_s.rd_addr = if_cfg_wst_s_rd_addr;
	assign if_cfg_est_m_wr_clk_en = if_cfg_est_m.wr_clk_en;
	assign if_cfg_wst_s.wr_clk_en = if_cfg_wst_s_wr_clk_en;
	assign if_cfg_est_m_rd_clk_en = if_cfg_est_m.rd_clk_en;
	assign if_cfg_wst_s.rd_clk_en = if_cfg_wst_s_rd_clk_en;
	assign if_cfg_est_m.rd_data = if_cfg_est_m_rd_data;
	assign if_cfg_wst_s_rd_data = if_cfg_wst_s.rd_data;
	assign if_cfg_est_m.rd_data_valid = if_cfg_est_m_rd_data_valid;
	assign if_cfg_wst_s_rd_data_valid = if_cfg_wst_s.rd_data_valid;
	assign strm_wr_packet_w2e_wsti[91] = strm_wr_en_w2e_wsti;
	assign strm_wr_packet_w2e_wsti[90-:8] = strm_wr_strb_w2e_wsti;
	assign strm_wr_packet_w2e_wsti[82-:19] = strm_wr_addr_w2e_wsti;
	assign strm_wr_packet_w2e_wsti[63-:64] = strm_wr_data_w2e_wsti;
	assign strm_wr_en_w2e_esto = strm_wr_packet_w2e_esto[91];
	assign strm_wr_strb_w2e_esto = strm_wr_packet_w2e_esto[90-:8];
	assign strm_wr_addr_w2e_esto = strm_wr_packet_w2e_esto[82-:19];
	assign strm_wr_data_w2e_esto = strm_wr_packet_w2e_esto[63-:64];
	assign strm_wr_packet_e2w_esti[91] = strm_wr_en_e2w_esti;
	assign strm_wr_packet_e2w_esti[90-:8] = strm_wr_strb_e2w_esti;
	assign strm_wr_packet_e2w_esti[82-:19] = strm_wr_addr_e2w_esti;
	assign strm_wr_packet_e2w_esti[63-:64] = strm_wr_data_e2w_esti;
	assign strm_wr_en_e2w_wsto = strm_wr_packet_e2w_wsto[91];
	assign strm_wr_strb_e2w_wsto = strm_wr_packet_e2w_wsto[90-:8];
	assign strm_wr_addr_e2w_wsto = strm_wr_packet_e2w_wsto[82-:19];
	assign strm_wr_data_e2w_wsto = strm_wr_packet_e2w_wsto[63-:64];
	assign strm_rdrq_packet_w2e_wsti[19] = strm_rd_en_w2e_wsti;
	assign strm_rdrq_packet_w2e_wsti[18-:19] = strm_rd_addr_w2e_wsti;
	assign strm_rd_en_w2e_esto = strm_rdrq_packet_w2e_esto[19];
	assign strm_rd_addr_w2e_esto = strm_rdrq_packet_w2e_esto[18-:19];
	assign strm_rdrq_packet_e2w_esti[19] = strm_rd_en_e2w_esti;
	assign strm_rdrq_packet_e2w_esti[18-:19] = strm_rd_addr_e2w_esti;
	assign strm_rd_en_e2w_wsto = strm_rdrq_packet_e2w_wsto[19];
	assign strm_rd_addr_e2w_wsto = strm_rdrq_packet_e2w_wsto[18-:19];
	assign strm_rd_data_e2w_wsto = strm_rdrs_packet_e2w_wsto[64-:64];
	assign strm_rd_data_valid_e2w_wsto = strm_rdrs_packet_e2w_wsto[0];
	assign strm_rdrs_packet_e2w_esti[64-:64] = strm_rd_data_e2w_esti;
	assign strm_rdrs_packet_e2w_esti[0] = strm_rd_data_valid_e2w_esti;
	assign strm_rdrs_packet_w2e_wsti[64-:64] = strm_rd_data_w2e_wsti;
	assign strm_rdrs_packet_w2e_wsti[0] = strm_rd_data_valid_w2e_wsti;
	assign strm_rd_data_w2e_esto = strm_rdrs_packet_w2e_esto[64-:64];
	assign strm_rd_data_valid_w2e_esto = strm_rdrs_packet_w2e_esto[0];
	assign pcfg_rdrq_packet_w2e_wsti[19] = pcfg_rd_en_w2e_wsti;
	assign pcfg_rdrq_packet_w2e_wsti[18-:19] = pcfg_rd_addr_w2e_wsti;
	assign pcfg_rd_en_w2e_esto = pcfg_rdrq_packet_w2e_esto[19];
	assign pcfg_rd_addr_w2e_esto = pcfg_rdrq_packet_w2e_esto[18-:19];
	assign pcfg_rdrq_packet_e2w_esti[19] = pcfg_rd_en_e2w_esti;
	assign pcfg_rdrq_packet_e2w_esti[18-:19] = pcfg_rd_addr_e2w_esti;
	assign pcfg_rd_en_e2w_wsto = pcfg_rdrq_packet_e2w_wsto[19];
	assign pcfg_rd_addr_e2w_wsto = pcfg_rdrq_packet_e2w_wsto[18-:19];
	assign pcfg_rd_data_e2w_wsto = pcfg_rdrs_packet_e2w_wsto[64-:64];
	assign pcfg_rd_data_valid_e2w_wsto = pcfg_rdrs_packet_e2w_wsto[0];
	assign pcfg_rdrs_packet_e2w_esti[64-:64] = pcfg_rd_data_e2w_esti;
	assign pcfg_rdrs_packet_e2w_esti[0] = pcfg_rd_data_valid_e2w_esti;
	assign pcfg_rdrs_packet_w2e_wsti[64-:64] = pcfg_rd_data_w2e_wsti;
	assign pcfg_rdrs_packet_w2e_wsti[0] = pcfg_rd_data_valid_w2e_wsti;
	assign pcfg_rd_data_w2e_esto = pcfg_rdrs_packet_w2e_esto[64-:64];
	assign pcfg_rd_data_valid_w2e_esto = pcfg_rdrs_packet_w2e_esto[0];
	assign clk_en_cfg = if_cfg_wst_s.wr_clk_en | if_cfg_wst_s.rd_clk_en;
	assign glb_clk_gate_cfg_enable = clk_en_cfg | clk_en_master;
	assign glb_clk_gate_pcfg_broadcast_enable = clk_en_pcfg_broadcast | clk_en_master;
	assign clk_en_ld_dma = cfg_ld_dma_ctrl[7-:2] != 2'h0;
	assign glb_clk_gate_ld_dma_enable = clk_en_ld_dma | clk_en_master;
	assign clk_en_st_dma = cfg_st_dma_ctrl[6-:2] != 2'h0;
	assign glb_clk_gate_st_dma_enable = clk_en_st_dma | clk_en_master;
	assign clk_en_proc_switch = if_proc_wst_s.wr_clk_en | if_proc_wst_s.rd_clk_en;
	assign glb_clk_gate_proc_switch_enable = clk_en_proc_switch | clk_en_master;
	assign clk_en_pcfg_dma = cfg_pcfg_dma_ctrl[17] != 1'h0;
	assign glb_clk_gate_pcfg_dma_enable = clk_en_pcfg_dma | clk_en_master;
	assign clk_en_strm_switch = cfg_tile_connected_next | cfg_tile_connected_prev;
	assign glb_clk_gate_strm_switch_enable = clk_en_strm_switch | clk_en_master;
	assign clk_en_pcfg_switch = cfg_pcfg_tile_connected_next | cfg_pcfg_tile_connected_prev;
	assign glb_clk_gate_pcfg_switch_enable = clk_en_pcfg_switch | clk_en_master;
	assign clk_en_bank = ((((clk_en_lddma2bank | clk_en_stdma2bank) | clk_en_pcfgdma2bank) | clk_en_ring2bank) | clk_en_pcfgring2bank) | clk_en_procsw2bank;
	assign glb_clk_gate_bank_enable = (clk_en_bank | clk_en_master) | clk_en_bank_master;
	assign cfg_tile_connected_next = glb_cfg_cfg_data_network[6];
	assign cfg_tile_connected_prev = cfg_tile_connected_wsti;
	assign cfg_tile_connected_esto = cfg_tile_connected_next;
	assign cfg_pcfg_tile_connected_next = glb_cfg_cfg_pcfg_network[6];
	assign cfg_pcfg_tile_connected_prev = cfg_pcfg_tile_connected_wsti;
	assign cfg_pcfg_tile_connected_esto = cfg_pcfg_tile_connected_next;
	assign glb_strm_ring_switch_cfg_ld_dma_on = cfg_ld_dma_ctrl[7-:2] != 2'h0;
	assign glb_pcfg_ring_switch_cfg_ld_dma_on = cfg_pcfg_dma_ctrl[17] != 1'h0;
	assign rdrs_packet_bankarr2sw[0+:65] = glb_bank_0_rdrs_packet;
	assign rdrs_packet_bankarr2sw[65+:65] = glb_bank_1_rdrs_packet;
	assign cgra_cfg_g2f_cfg_wr_en[0] = cgra_cfg_g2f_cfg_w[64];
	assign cgra_cfg_g2f_cfg_rd_en[0] = cgra_cfg_g2f_cfg_w[65];
	assign cgra_cfg_g2f_cfg_addr[0+:32] = cgra_cfg_g2f_cfg_w[63-:32];
	assign cgra_cfg_g2f_cfg_data[0+:32] = cgra_cfg_g2f_cfg_w[31-:32];
	assign cgra_cfg_g2f_cfg_wr_en[1] = cgra_cfg_g2f_cfg_w[130];
	assign cgra_cfg_g2f_cfg_rd_en[1] = cgra_cfg_g2f_cfg_w[131];
	assign cgra_cfg_g2f_cfg_addr[32+:32] = cgra_cfg_g2f_cfg_w[129-:32];
	assign cgra_cfg_g2f_cfg_data[32+:32] = cgra_cfg_g2f_cfg_w[97-:32];
	assign glb_pcfg_broadcast_cgra_cfg_jtag_wsti[64] = cgra_cfg_jtag_wr_en_wsti;
	assign glb_pcfg_broadcast_cgra_cfg_jtag_wsti[65] = cgra_cfg_jtag_rd_en_wsti;
	assign glb_pcfg_broadcast_cgra_cfg_jtag_wsti[63-:32] = cgra_cfg_jtag_addr_wsti;
	assign glb_pcfg_broadcast_cgra_cfg_jtag_wsti[31-:32] = cgra_cfg_jtag_data_wsti;
	assign cgra_cfg_jtag_wr_en_esto = glb_pcfg_broadcast_cgra_cfg_jtag_esto[64];
	assign cgra_cfg_jtag_rd_en_esto = glb_pcfg_broadcast_cgra_cfg_jtag_esto[65];
	assign cgra_cfg_jtag_addr_esto = glb_pcfg_broadcast_cgra_cfg_jtag_esto[63-:32];
	assign cgra_cfg_jtag_data_esto = glb_pcfg_broadcast_cgra_cfg_jtag_esto[31-:32];
	assign glb_pcfg_broadcast_cgra_cfg_pcfg_wsti[64] = cgra_cfg_pcfg_wr_en_w2e_wsti;
	assign glb_pcfg_broadcast_cgra_cfg_pcfg_wsti[65] = cgra_cfg_pcfg_rd_en_w2e_wsti;
	assign glb_pcfg_broadcast_cgra_cfg_pcfg_wsti[63-:32] = cgra_cfg_pcfg_addr_w2e_wsti;
	assign glb_pcfg_broadcast_cgra_cfg_pcfg_wsti[31-:32] = cgra_cfg_pcfg_data_w2e_wsti;
	assign cgra_cfg_pcfg_wr_en_w2e_esto = glb_pcfg_broadcast_cgra_cfg_pcfg_esto[64];
	assign cgra_cfg_pcfg_rd_en_w2e_esto = glb_pcfg_broadcast_cgra_cfg_pcfg_esto[65];
	assign cgra_cfg_pcfg_addr_w2e_esto = glb_pcfg_broadcast_cgra_cfg_pcfg_esto[63-:32];
	assign cgra_cfg_pcfg_data_w2e_esto = glb_pcfg_broadcast_cgra_cfg_pcfg_esto[31-:32];
	assign glb_pcfg_broadcast_cgra_cfg_pcfg_esti[64] = cgra_cfg_pcfg_wr_en_e2w_esti;
	assign glb_pcfg_broadcast_cgra_cfg_pcfg_esti[65] = cgra_cfg_pcfg_rd_en_e2w_esti;
	assign glb_pcfg_broadcast_cgra_cfg_pcfg_esti[63-:32] = cgra_cfg_pcfg_addr_e2w_esti;
	assign glb_pcfg_broadcast_cgra_cfg_pcfg_esti[31-:32] = cgra_cfg_pcfg_data_e2w_esti;
	assign cgra_cfg_pcfg_wr_en_e2w_wsto = glb_pcfg_broadcast_cgra_cfg_pcfg_wsto[64];
	assign cgra_cfg_pcfg_rd_en_e2w_wsto = glb_pcfg_broadcast_cgra_cfg_pcfg_wsto[65];
	assign cgra_cfg_pcfg_addr_e2w_wsto = glb_pcfg_broadcast_cgra_cfg_pcfg_wsto[63-:32];
	assign cgra_cfg_pcfg_data_e2w_wsto = glb_pcfg_broadcast_cgra_cfg_pcfg_wsto[31-:32];
	clk_gate glb_clk_gate_cfg(
		.clk(clk),
		.enable(glb_clk_gate_cfg_enable),
		.gclk(gclk_cfg)
	);
	clk_gate glb_clk_gate_pcfg_broadcast(
		.clk(clk),
		.enable(glb_clk_gate_pcfg_broadcast_enable),
		.gclk(gclk_pcfg_broadcast)
	);
	clk_gate glb_clk_gate_ld_dma(
		.clk(clk),
		.enable(glb_clk_gate_ld_dma_enable),
		.gclk(gclk_ld_dma)
	);
	clk_gate glb_clk_gate_st_dma(
		.clk(clk),
		.enable(glb_clk_gate_st_dma_enable),
		.gclk(gclk_st_dma)
	);
	clk_gate glb_clk_gate_proc_switch(
		.clk(clk),
		.enable(glb_clk_gate_proc_switch_enable),
		.gclk(gclk_proc_switch)
	);
	clk_gate glb_clk_gate_pcfg_dma(
		.clk(clk),
		.enable(glb_clk_gate_pcfg_dma_enable),
		.gclk(gclk_pcfg_dma)
	);
	clk_gate glb_clk_gate_strm_switch(
		.clk(clk),
		.enable(glb_clk_gate_strm_switch_enable),
		.gclk(gclk_strm_switch)
	);
	clk_gate glb_clk_gate_pcfg_switch(
		.clk(clk),
		.enable(glb_clk_gate_pcfg_switch_enable),
		.gclk(gclk_pcfg_switch)
	);
	clk_gate glb_clk_gate_bank(
		.clk(clk),
		.enable(glb_clk_gate_bank_enable),
		.gclk(gclk_bank)
	);
	generate
		if (1) begin : glb_cfg
			wire gclk;
			wire glb_tile_id;
			wire mclk;
			wire reset;
			wire [6:0] cfg_data_network;
			wire [7:0] cfg_ld_dma_ctrl;
			wire [582:0] cfg_ld_dma_header;
			wire [5:0] cfg_pcfg_broadcast_mux;
			wire [17:0] cfg_pcfg_dma_ctrl;
			wire [34:0] cfg_pcfg_dma_header;
			wire [6:0] cfg_pcfg_network;
			wire [6:0] cfg_st_dma_ctrl;
			wire [514:0] cfg_st_dma_header;
			wire [31:0] cfg_st_dma_num_blocks;
			wire [8:0] glb_cfg_ctrl_h2d_pio_dec_address;
			wire glb_pio_d2h_dec_pio_ack;
			wire glb_pio_d2h_dec_pio_nack;
			wire [31:0] glb_pio_d2h_dec_pio_read_data;
			wire [5:0] glb_pio_h2d_pio_dec_address;
			wire glb_pio_h2d_pio_dec_read;
			wire glb_pio_h2d_pio_dec_write;
			wire [31:0] glb_pio_h2d_pio_dec_write_data;
			wire glb_pio_l2h_data_network_ctrl_connected_r;
			wire [5:0] glb_pio_l2h_data_network_latency_value_r;
			wire [1:0] glb_pio_l2h_ld_dma_ctrl_data_mux_r;
			wire glb_pio_l2h_ld_dma_ctrl_flush_mode_r;
			wire [1:0] glb_pio_l2h_ld_dma_ctrl_mode_r;
			wire glb_pio_l2h_ld_dma_ctrl_num_repeat_r;
			wire [1:0] glb_pio_l2h_ld_dma_ctrl_valid_mode_r;
			wire [15:0] glb_pio_l2h_ld_dma_header_0_cycle_start_addr_cycle_start_addr_r;
			wire [15:0] glb_pio_l2h_ld_dma_header_0_cycle_stride_0_cycle_stride_r;
			wire [15:0] glb_pio_l2h_ld_dma_header_0_cycle_stride_1_cycle_stride_r;
			wire [15:0] glb_pio_l2h_ld_dma_header_0_cycle_stride_2_cycle_stride_r;
			wire [15:0] glb_pio_l2h_ld_dma_header_0_cycle_stride_3_cycle_stride_r;
			wire [15:0] glb_pio_l2h_ld_dma_header_0_cycle_stride_4_cycle_stride_r;
			wire [15:0] glb_pio_l2h_ld_dma_header_0_cycle_stride_5_cycle_stride_r;
			wire [15:0] glb_pio_l2h_ld_dma_header_0_cycle_stride_6_cycle_stride_r;
			wire [15:0] glb_pio_l2h_ld_dma_header_0_cycle_stride_7_cycle_stride_r;
			wire [3:0] glb_pio_l2h_ld_dma_header_0_dim_dim_r;
			wire [31:0] glb_pio_l2h_ld_dma_header_0_range_0_range_r;
			wire [31:0] glb_pio_l2h_ld_dma_header_0_range_1_range_r;
			wire [31:0] glb_pio_l2h_ld_dma_header_0_range_2_range_r;
			wire [31:0] glb_pio_l2h_ld_dma_header_0_range_3_range_r;
			wire [31:0] glb_pio_l2h_ld_dma_header_0_range_4_range_r;
			wire [31:0] glb_pio_l2h_ld_dma_header_0_range_5_range_r;
			wire [31:0] glb_pio_l2h_ld_dma_header_0_range_6_range_r;
			wire [31:0] glb_pio_l2h_ld_dma_header_0_range_7_range_r;
			wire [18:0] glb_pio_l2h_ld_dma_header_0_start_addr_start_addr_r;
			wire [19:0] glb_pio_l2h_ld_dma_header_0_stride_0_stride_r;
			wire [19:0] glb_pio_l2h_ld_dma_header_0_stride_1_stride_r;
			wire [19:0] glb_pio_l2h_ld_dma_header_0_stride_2_stride_r;
			wire [19:0] glb_pio_l2h_ld_dma_header_0_stride_3_stride_r;
			wire [19:0] glb_pio_l2h_ld_dma_header_0_stride_4_stride_r;
			wire [19:0] glb_pio_l2h_ld_dma_header_0_stride_5_stride_r;
			wire [19:0] glb_pio_l2h_ld_dma_header_0_stride_6_stride_r;
			wire [19:0] glb_pio_l2h_ld_dma_header_0_stride_7_stride_r;
			wire [1:0] glb_pio_l2h_pcfg_broadcast_mux_east_r;
			wire [1:0] glb_pio_l2h_pcfg_broadcast_mux_south_r;
			wire [1:0] glb_pio_l2h_pcfg_broadcast_mux_west_r;
			wire glb_pio_l2h_pcfg_dma_ctrl_mode_r;
			wire glb_pio_l2h_pcfg_dma_ctrl_relocation_is_msb_r;
			wire [15:0] glb_pio_l2h_pcfg_dma_ctrl_relocation_value_r;
			wire [15:0] glb_pio_l2h_pcfg_dma_header_num_cfg_num_cfg_r;
			wire [18:0] glb_pio_l2h_pcfg_dma_header_start_addr_start_addr_r;
			wire glb_pio_l2h_pcfg_network_ctrl_connected_r;
			wire [5:0] glb_pio_l2h_pcfg_network_latency_value_r;
			wire [1:0] glb_pio_l2h_st_dma_ctrl_data_mux_r;
			wire [1:0] glb_pio_l2h_st_dma_ctrl_mode_r;
			wire glb_pio_l2h_st_dma_ctrl_num_repeat_r;
			wire [1:0] glb_pio_l2h_st_dma_ctrl_valid_mode_r;
			wire [15:0] glb_pio_l2h_st_dma_header_0_cycle_start_addr_cycle_start_addr_r;
			wire [15:0] glb_pio_l2h_st_dma_header_0_cycle_stride_0_cycle_stride_r;
			wire [15:0] glb_pio_l2h_st_dma_header_0_cycle_stride_1_cycle_stride_r;
			wire [15:0] glb_pio_l2h_st_dma_header_0_cycle_stride_2_cycle_stride_r;
			wire [15:0] glb_pio_l2h_st_dma_header_0_cycle_stride_3_cycle_stride_r;
			wire [15:0] glb_pio_l2h_st_dma_header_0_cycle_stride_4_cycle_stride_r;
			wire [15:0] glb_pio_l2h_st_dma_header_0_cycle_stride_5_cycle_stride_r;
			wire [15:0] glb_pio_l2h_st_dma_header_0_cycle_stride_6_cycle_stride_r;
			wire [3:0] glb_pio_l2h_st_dma_header_0_dim_dim_r;
			wire [31:0] glb_pio_l2h_st_dma_header_0_range_0_range_r;
			wire [31:0] glb_pio_l2h_st_dma_header_0_range_1_range_r;
			wire [31:0] glb_pio_l2h_st_dma_header_0_range_2_range_r;
			wire [31:0] glb_pio_l2h_st_dma_header_0_range_3_range_r;
			wire [31:0] glb_pio_l2h_st_dma_header_0_range_4_range_r;
			wire [31:0] glb_pio_l2h_st_dma_header_0_range_5_range_r;
			wire [31:0] glb_pio_l2h_st_dma_header_0_range_6_range_r;
			wire [18:0] glb_pio_l2h_st_dma_header_0_start_addr_start_addr_r;
			wire [19:0] glb_pio_l2h_st_dma_header_0_stride_0_stride_r;
			wire [19:0] glb_pio_l2h_st_dma_header_0_stride_1_stride_r;
			wire [19:0] glb_pio_l2h_st_dma_header_0_stride_2_stride_r;
			wire [19:0] glb_pio_l2h_st_dma_header_0_stride_3_stride_r;
			wire [19:0] glb_pio_l2h_st_dma_header_0_stride_4_stride_r;
			wire [19:0] glb_pio_l2h_st_dma_header_0_stride_5_stride_r;
			wire [19:0] glb_pio_l2h_st_dma_header_0_stride_6_stride_r;
			assign cfg_data_network[6] = glb_pio_l2h_data_network_ctrl_connected_r;
			assign cfg_data_network[5-:6] = glb_pio_l2h_data_network_latency_value_r;
			assign cfg_pcfg_network[6] = glb_pio_l2h_pcfg_network_ctrl_connected_r;
			assign cfg_pcfg_network[5-:6] = glb_pio_l2h_pcfg_network_latency_value_r;
			assign cfg_st_dma_ctrl[2-:2] = glb_pio_l2h_st_dma_ctrl_data_mux_r;
			assign cfg_st_dma_ctrl[6-:2] = glb_pio_l2h_st_dma_ctrl_mode_r;
			assign cfg_st_dma_ctrl[4-:2] = glb_pio_l2h_st_dma_ctrl_valid_mode_r;
			assign cfg_st_dma_ctrl[0] = glb_pio_l2h_st_dma_ctrl_num_repeat_r;
			assign cfg_st_dma_header[514-:19] = glb_pio_l2h_st_dma_header_0_start_addr_start_addr_r;
			assign cfg_st_dma_header[495-:16] = glb_pio_l2h_st_dma_header_0_cycle_start_addr_cycle_start_addr_r;
			assign cfg_st_dma_header[479-:4] = glb_pio_l2h_st_dma_header_0_dim_dim_r;
			assign cfg_st_dma_header[423-:16] = glb_pio_l2h_st_dma_header_0_cycle_stride_0_cycle_stride_r;
			assign cfg_st_dma_header[443-:20] = glb_pio_l2h_st_dma_header_0_stride_0_stride_r;
			assign cfg_st_dma_header[475-:32] = glb_pio_l2h_st_dma_header_0_range_0_range_r;
			assign cfg_st_dma_header[355-:16] = glb_pio_l2h_st_dma_header_0_cycle_stride_1_cycle_stride_r;
			assign cfg_st_dma_header[375-:20] = glb_pio_l2h_st_dma_header_0_stride_1_stride_r;
			assign cfg_st_dma_header[407-:32] = glb_pio_l2h_st_dma_header_0_range_1_range_r;
			assign cfg_st_dma_header[287-:16] = glb_pio_l2h_st_dma_header_0_cycle_stride_2_cycle_stride_r;
			assign cfg_st_dma_header[307-:20] = glb_pio_l2h_st_dma_header_0_stride_2_stride_r;
			assign cfg_st_dma_header[339-:32] = glb_pio_l2h_st_dma_header_0_range_2_range_r;
			assign cfg_st_dma_header[219-:16] = glb_pio_l2h_st_dma_header_0_cycle_stride_3_cycle_stride_r;
			assign cfg_st_dma_header[239-:20] = glb_pio_l2h_st_dma_header_0_stride_3_stride_r;
			assign cfg_st_dma_header[271-:32] = glb_pio_l2h_st_dma_header_0_range_3_range_r;
			assign cfg_st_dma_header[151-:16] = glb_pio_l2h_st_dma_header_0_cycle_stride_4_cycle_stride_r;
			assign cfg_st_dma_header[171-:20] = glb_pio_l2h_st_dma_header_0_stride_4_stride_r;
			assign cfg_st_dma_header[203-:32] = glb_pio_l2h_st_dma_header_0_range_4_range_r;
			assign cfg_st_dma_header[83-:16] = glb_pio_l2h_st_dma_header_0_cycle_stride_5_cycle_stride_r;
			assign cfg_st_dma_header[103-:20] = glb_pio_l2h_st_dma_header_0_stride_5_stride_r;
			assign cfg_st_dma_header[135-:32] = glb_pio_l2h_st_dma_header_0_range_5_range_r;
			assign cfg_st_dma_header[15-:16] = glb_pio_l2h_st_dma_header_0_cycle_stride_6_cycle_stride_r;
			assign cfg_st_dma_header[35-:20] = glb_pio_l2h_st_dma_header_0_stride_6_stride_r;
			assign cfg_st_dma_header[67-:32] = glb_pio_l2h_st_dma_header_0_range_6_range_r;
			assign cfg_ld_dma_ctrl[2-:2] = glb_pio_l2h_ld_dma_ctrl_data_mux_r;
			assign cfg_ld_dma_ctrl[7-:2] = glb_pio_l2h_ld_dma_ctrl_mode_r;
			assign cfg_ld_dma_ctrl[5-:2] = glb_pio_l2h_ld_dma_ctrl_valid_mode_r;
			assign cfg_ld_dma_ctrl[3] = glb_pio_l2h_ld_dma_ctrl_flush_mode_r;
			assign cfg_ld_dma_ctrl[0] = glb_pio_l2h_ld_dma_ctrl_num_repeat_r;
			assign cfg_ld_dma_header[582-:19] = glb_pio_l2h_ld_dma_header_0_start_addr_start_addr_r;
			assign cfg_ld_dma_header[563-:16] = glb_pio_l2h_ld_dma_header_0_cycle_start_addr_cycle_start_addr_r;
			assign cfg_ld_dma_header[547-:4] = glb_pio_l2h_ld_dma_header_0_dim_dim_r;
			assign cfg_ld_dma_header[491-:16] = glb_pio_l2h_ld_dma_header_0_cycle_stride_0_cycle_stride_r;
			assign cfg_ld_dma_header[511-:20] = glb_pio_l2h_ld_dma_header_0_stride_0_stride_r;
			assign cfg_ld_dma_header[543-:32] = glb_pio_l2h_ld_dma_header_0_range_0_range_r;
			assign cfg_ld_dma_header[423-:16] = glb_pio_l2h_ld_dma_header_0_cycle_stride_1_cycle_stride_r;
			assign cfg_ld_dma_header[443-:20] = glb_pio_l2h_ld_dma_header_0_stride_1_stride_r;
			assign cfg_ld_dma_header[475-:32] = glb_pio_l2h_ld_dma_header_0_range_1_range_r;
			assign cfg_ld_dma_header[355-:16] = glb_pio_l2h_ld_dma_header_0_cycle_stride_2_cycle_stride_r;
			assign cfg_ld_dma_header[375-:20] = glb_pio_l2h_ld_dma_header_0_stride_2_stride_r;
			assign cfg_ld_dma_header[407-:32] = glb_pio_l2h_ld_dma_header_0_range_2_range_r;
			assign cfg_ld_dma_header[287-:16] = glb_pio_l2h_ld_dma_header_0_cycle_stride_3_cycle_stride_r;
			assign cfg_ld_dma_header[307-:20] = glb_pio_l2h_ld_dma_header_0_stride_3_stride_r;
			assign cfg_ld_dma_header[339-:32] = glb_pio_l2h_ld_dma_header_0_range_3_range_r;
			assign cfg_ld_dma_header[219-:16] = glb_pio_l2h_ld_dma_header_0_cycle_stride_4_cycle_stride_r;
			assign cfg_ld_dma_header[239-:20] = glb_pio_l2h_ld_dma_header_0_stride_4_stride_r;
			assign cfg_ld_dma_header[271-:32] = glb_pio_l2h_ld_dma_header_0_range_4_range_r;
			assign cfg_ld_dma_header[151-:16] = glb_pio_l2h_ld_dma_header_0_cycle_stride_5_cycle_stride_r;
			assign cfg_ld_dma_header[171-:20] = glb_pio_l2h_ld_dma_header_0_stride_5_stride_r;
			assign cfg_ld_dma_header[203-:32] = glb_pio_l2h_ld_dma_header_0_range_5_range_r;
			assign cfg_ld_dma_header[83-:16] = glb_pio_l2h_ld_dma_header_0_cycle_stride_6_cycle_stride_r;
			assign cfg_ld_dma_header[103-:20] = glb_pio_l2h_ld_dma_header_0_stride_6_stride_r;
			assign cfg_ld_dma_header[135-:32] = glb_pio_l2h_ld_dma_header_0_range_6_range_r;
			assign cfg_ld_dma_header[15-:16] = glb_pio_l2h_ld_dma_header_0_cycle_stride_7_cycle_stride_r;
			assign cfg_ld_dma_header[35-:20] = glb_pio_l2h_ld_dma_header_0_stride_7_stride_r;
			assign cfg_ld_dma_header[67-:32] = glb_pio_l2h_ld_dma_header_0_range_7_range_r;
			assign cfg_pcfg_dma_ctrl[17] = glb_pio_l2h_pcfg_dma_ctrl_mode_r;
			assign cfg_pcfg_dma_ctrl[16-:16] = glb_pio_l2h_pcfg_dma_ctrl_relocation_value_r;
			assign cfg_pcfg_dma_ctrl[0] = glb_pio_l2h_pcfg_dma_ctrl_relocation_is_msb_r;
			assign cfg_pcfg_dma_header[34-:19] = glb_pio_l2h_pcfg_dma_header_start_addr_start_addr_r;
			assign cfg_pcfg_dma_header[15-:16] = glb_pio_l2h_pcfg_dma_header_num_cfg_num_cfg_r;
			assign cfg_pcfg_broadcast_mux[5-:2] = glb_pio_l2h_pcfg_broadcast_mux_west_r;
			assign cfg_pcfg_broadcast_mux[3-:2] = glb_pio_l2h_pcfg_broadcast_mux_east_r;
			assign cfg_pcfg_broadcast_mux[1-:2] = glb_pio_l2h_pcfg_broadcast_mux_south_r;
			assign glb_pio_h2d_pio_dec_address = glb_cfg_ctrl_h2d_pio_dec_address[5:0];
			glb_pio glb_pio(
				.clk(gclk),
				.h2d_pio_dec_address(glb_pio_h2d_pio_dec_address),
				.h2d_pio_dec_read(glb_pio_h2d_pio_dec_read),
				.h2d_pio_dec_write(glb_pio_h2d_pio_dec_write),
				.h2d_pio_dec_write_data(glb_pio_h2d_pio_dec_write_data),
				.reset(reset),
				.d2h_dec_pio_ack(glb_pio_d2h_dec_pio_ack),
				.d2h_dec_pio_nack(glb_pio_d2h_dec_pio_nack),
				.d2h_dec_pio_read_data(glb_pio_d2h_dec_pio_read_data),
				.l2h_data_network_ctrl_connected_r(glb_pio_l2h_data_network_ctrl_connected_r),
				.l2h_data_network_latency_value_r(glb_pio_l2h_data_network_latency_value_r),
				.l2h_ld_dma_ctrl_data_mux_r(glb_pio_l2h_ld_dma_ctrl_data_mux_r),
				.l2h_ld_dma_ctrl_flush_mode_r(glb_pio_l2h_ld_dma_ctrl_flush_mode_r),
				.l2h_ld_dma_ctrl_mode_r(glb_pio_l2h_ld_dma_ctrl_mode_r),
				.l2h_ld_dma_ctrl_num_repeat_r(glb_pio_l2h_ld_dma_ctrl_num_repeat_r),
				.l2h_ld_dma_ctrl_valid_mode_r(glb_pio_l2h_ld_dma_ctrl_valid_mode_r),
				.l2h_ld_dma_header_0_cycle_start_addr_cycle_start_addr_r(glb_pio_l2h_ld_dma_header_0_cycle_start_addr_cycle_start_addr_r),
				.l2h_ld_dma_header_0_cycle_stride_0_cycle_stride_r(glb_pio_l2h_ld_dma_header_0_cycle_stride_0_cycle_stride_r),
				.l2h_ld_dma_header_0_cycle_stride_1_cycle_stride_r(glb_pio_l2h_ld_dma_header_0_cycle_stride_1_cycle_stride_r),
				.l2h_ld_dma_header_0_cycle_stride_2_cycle_stride_r(glb_pio_l2h_ld_dma_header_0_cycle_stride_2_cycle_stride_r),
				.l2h_ld_dma_header_0_cycle_stride_3_cycle_stride_r(glb_pio_l2h_ld_dma_header_0_cycle_stride_3_cycle_stride_r),
				.l2h_ld_dma_header_0_cycle_stride_4_cycle_stride_r(glb_pio_l2h_ld_dma_header_0_cycle_stride_4_cycle_stride_r),
				.l2h_ld_dma_header_0_cycle_stride_5_cycle_stride_r(glb_pio_l2h_ld_dma_header_0_cycle_stride_5_cycle_stride_r),
				.l2h_ld_dma_header_0_cycle_stride_6_cycle_stride_r(glb_pio_l2h_ld_dma_header_0_cycle_stride_6_cycle_stride_r),
				.l2h_ld_dma_header_0_cycle_stride_7_cycle_stride_r(glb_pio_l2h_ld_dma_header_0_cycle_stride_7_cycle_stride_r),
				.l2h_ld_dma_header_0_dim_dim_r(glb_pio_l2h_ld_dma_header_0_dim_dim_r),
				.l2h_ld_dma_header_0_range_0_range_r(glb_pio_l2h_ld_dma_header_0_range_0_range_r),
				.l2h_ld_dma_header_0_range_1_range_r(glb_pio_l2h_ld_dma_header_0_range_1_range_r),
				.l2h_ld_dma_header_0_range_2_range_r(glb_pio_l2h_ld_dma_header_0_range_2_range_r),
				.l2h_ld_dma_header_0_range_3_range_r(glb_pio_l2h_ld_dma_header_0_range_3_range_r),
				.l2h_ld_dma_header_0_range_4_range_r(glb_pio_l2h_ld_dma_header_0_range_4_range_r),
				.l2h_ld_dma_header_0_range_5_range_r(glb_pio_l2h_ld_dma_header_0_range_5_range_r),
				.l2h_ld_dma_header_0_range_6_range_r(glb_pio_l2h_ld_dma_header_0_range_6_range_r),
				.l2h_ld_dma_header_0_range_7_range_r(glb_pio_l2h_ld_dma_header_0_range_7_range_r),
				.l2h_ld_dma_header_0_start_addr_start_addr_r(glb_pio_l2h_ld_dma_header_0_start_addr_start_addr_r),
				.l2h_ld_dma_header_0_stride_0_stride_r(glb_pio_l2h_ld_dma_header_0_stride_0_stride_r),
				.l2h_ld_dma_header_0_stride_1_stride_r(glb_pio_l2h_ld_dma_header_0_stride_1_stride_r),
				.l2h_ld_dma_header_0_stride_2_stride_r(glb_pio_l2h_ld_dma_header_0_stride_2_stride_r),
				.l2h_ld_dma_header_0_stride_3_stride_r(glb_pio_l2h_ld_dma_header_0_stride_3_stride_r),
				.l2h_ld_dma_header_0_stride_4_stride_r(glb_pio_l2h_ld_dma_header_0_stride_4_stride_r),
				.l2h_ld_dma_header_0_stride_5_stride_r(glb_pio_l2h_ld_dma_header_0_stride_5_stride_r),
				.l2h_ld_dma_header_0_stride_6_stride_r(glb_pio_l2h_ld_dma_header_0_stride_6_stride_r),
				.l2h_ld_dma_header_0_stride_7_stride_r(glb_pio_l2h_ld_dma_header_0_stride_7_stride_r),
				.l2h_pcfg_broadcast_mux_east_r(glb_pio_l2h_pcfg_broadcast_mux_east_r),
				.l2h_pcfg_broadcast_mux_south_r(glb_pio_l2h_pcfg_broadcast_mux_south_r),
				.l2h_pcfg_broadcast_mux_west_r(glb_pio_l2h_pcfg_broadcast_mux_west_r),
				.l2h_pcfg_dma_ctrl_mode_r(glb_pio_l2h_pcfg_dma_ctrl_mode_r),
				.l2h_pcfg_dma_ctrl_relocation_is_msb_r(glb_pio_l2h_pcfg_dma_ctrl_relocation_is_msb_r),
				.l2h_pcfg_dma_ctrl_relocation_value_r(glb_pio_l2h_pcfg_dma_ctrl_relocation_value_r),
				.l2h_pcfg_dma_header_num_cfg_num_cfg_r(glb_pio_l2h_pcfg_dma_header_num_cfg_num_cfg_r),
				.l2h_pcfg_dma_header_start_addr_start_addr_r(glb_pio_l2h_pcfg_dma_header_start_addr_start_addr_r),
				.l2h_pcfg_network_ctrl_connected_r(glb_pio_l2h_pcfg_network_ctrl_connected_r),
				.l2h_pcfg_network_latency_value_r(glb_pio_l2h_pcfg_network_latency_value_r),
				.l2h_st_dma_ctrl_data_mux_r(glb_pio_l2h_st_dma_ctrl_data_mux_r),
				.l2h_st_dma_ctrl_mode_r(glb_pio_l2h_st_dma_ctrl_mode_r),
				.l2h_st_dma_ctrl_num_repeat_r(glb_pio_l2h_st_dma_ctrl_num_repeat_r),
				.l2h_st_dma_ctrl_valid_mode_r(glb_pio_l2h_st_dma_ctrl_valid_mode_r),
				.l2h_st_dma_header_0_cycle_start_addr_cycle_start_addr_r(glb_pio_l2h_st_dma_header_0_cycle_start_addr_cycle_start_addr_r),
				.l2h_st_dma_header_0_cycle_stride_0_cycle_stride_r(glb_pio_l2h_st_dma_header_0_cycle_stride_0_cycle_stride_r),
				.l2h_st_dma_header_0_cycle_stride_1_cycle_stride_r(glb_pio_l2h_st_dma_header_0_cycle_stride_1_cycle_stride_r),
				.l2h_st_dma_header_0_cycle_stride_2_cycle_stride_r(glb_pio_l2h_st_dma_header_0_cycle_stride_2_cycle_stride_r),
				.l2h_st_dma_header_0_cycle_stride_3_cycle_stride_r(glb_pio_l2h_st_dma_header_0_cycle_stride_3_cycle_stride_r),
				.l2h_st_dma_header_0_cycle_stride_4_cycle_stride_r(glb_pio_l2h_st_dma_header_0_cycle_stride_4_cycle_stride_r),
				.l2h_st_dma_header_0_cycle_stride_5_cycle_stride_r(glb_pio_l2h_st_dma_header_0_cycle_stride_5_cycle_stride_r),
				.l2h_st_dma_header_0_cycle_stride_6_cycle_stride_r(glb_pio_l2h_st_dma_header_0_cycle_stride_6_cycle_stride_r),
				.l2h_st_dma_header_0_dim_dim_r(glb_pio_l2h_st_dma_header_0_dim_dim_r),
				.l2h_st_dma_header_0_range_0_range_r(glb_pio_l2h_st_dma_header_0_range_0_range_r),
				.l2h_st_dma_header_0_range_1_range_r(glb_pio_l2h_st_dma_header_0_range_1_range_r),
				.l2h_st_dma_header_0_range_2_range_r(glb_pio_l2h_st_dma_header_0_range_2_range_r),
				.l2h_st_dma_header_0_range_3_range_r(glb_pio_l2h_st_dma_header_0_range_3_range_r),
				.l2h_st_dma_header_0_range_4_range_r(glb_pio_l2h_st_dma_header_0_range_4_range_r),
				.l2h_st_dma_header_0_range_5_range_r(glb_pio_l2h_st_dma_header_0_range_5_range_r),
				.l2h_st_dma_header_0_range_6_range_r(glb_pio_l2h_st_dma_header_0_range_6_range_r),
				.l2h_st_dma_header_0_start_addr_start_addr_r(glb_pio_l2h_st_dma_header_0_start_addr_start_addr_r),
				.l2h_st_dma_header_0_stride_0_stride_r(glb_pio_l2h_st_dma_header_0_stride_0_stride_r),
				.l2h_st_dma_header_0_stride_1_stride_r(glb_pio_l2h_st_dma_header_0_stride_1_stride_r),
				.l2h_st_dma_header_0_stride_2_stride_r(glb_pio_l2h_st_dma_header_0_stride_2_stride_r),
				.l2h_st_dma_header_0_stride_3_stride_r(glb_pio_l2h_st_dma_header_0_stride_3_stride_r),
				.l2h_st_dma_header_0_stride_4_stride_r(glb_pio_l2h_st_dma_header_0_stride_4_stride_r),
				.l2h_st_dma_header_0_stride_5_stride_r(glb_pio_l2h_st_dma_header_0_stride_5_stride_r),
				.l2h_st_dma_header_0_stride_6_stride_r(glb_pio_l2h_st_dma_header_0_stride_6_stride_r),
				.l2h_st_dma_num_blocks_value_r(cfg_st_dma_num_blocks)
			);
			if (1) begin : glb_cfg_ctrl
				wire d2h_dec_pio_ack;
				wire d2h_dec_pio_nack;
				wire [31:0] d2h_dec_pio_read_data;
				wire gclk;
				wire glb_tile_id;
				wire mclk;
				wire reset;
				wire [8:0] h2d_pio_dec_address;
				wire h2d_pio_dec_read;
				wire h2d_pio_dec_write;
				wire [31:0] h2d_pio_dec_write_data;
				reg [8:0] addr_internal;
				reg if_cfg_est_m_rd_clk_en_sel;
				reg if_cfg_est_m_rd_clk_en_sel_first_cycle;
				reg if_cfg_est_m_rd_clk_en_sel_latch;
				reg if_cfg_est_m_wr_clk_en_sel;
				reg if_cfg_est_m_wr_clk_en_sel_first_cycle;
				reg if_cfg_est_m_wr_clk_en_sel_latch;
				reg if_cfg_wst_s_rd_clk_en_d;
				reg if_cfg_wst_s_wr_clk_en_d;
				reg [31:0] rd_data_internal;
				reg rd_data_valid_internal;
				reg rd_en_d1;
				reg rd_en_d2;
				reg rd_tile_id_match;
				reg read_internal;
				reg [31:0] wr_data_internal;
				reg wr_tile_id_match;
				reg write_internal;
				always @(*) begin
					wr_tile_id_match = glb_tile_id == glb_tile.if_cfg_wst_s.wr_addr[11];
					rd_tile_id_match = glb_tile_id == glb_tile.if_cfg_wst_s.rd_addr[11];
				end
				always @(*) begin
					wr_data_internal = 32'h00000000;
					addr_internal = 9'h000;
					read_internal = 1'h0;
					write_internal = 1'h0;
					if (glb_tile.if_cfg_wst_s.rd_en && rd_tile_id_match) begin
						addr_internal = glb_tile.if_cfg_wst_s.rd_addr[10:2];
						read_internal = 1'h1;
					end
					if (glb_tile.if_cfg_wst_s.wr_en && wr_tile_id_match) begin
						addr_internal = glb_tile.if_cfg_wst_s.wr_addr[10:2];
						wr_data_internal = glb_tile.if_cfg_wst_s.wr_data;
						write_internal = 1'h1;
					end
				end
				always @(posedge gclk or posedge reset)
					if (reset) begin
						glb_tile.if_cfg_est_m.wr_en <= 1'h0;
						glb_tile.if_cfg_est_m.wr_addr <= 12'h000;
						glb_tile.if_cfg_est_m.wr_data <= 32'h00000000;
					end
					else if (~(wr_tile_id_match && (glb_tile.if_cfg_wst_s.wr_en == 1'h1))) begin
						glb_tile.if_cfg_est_m.wr_en <= glb_tile.if_cfg_wst_s.wr_en;
						glb_tile.if_cfg_est_m.wr_addr <= glb_tile.if_cfg_wst_s.wr_addr;
						glb_tile.if_cfg_est_m.wr_data <= glb_tile.if_cfg_wst_s.wr_data;
					end
					else begin
						glb_tile.if_cfg_est_m.wr_en <= 1'h0;
						glb_tile.if_cfg_est_m.wr_addr <= 12'h000;
						glb_tile.if_cfg_est_m.wr_data <= 32'h00000000;
					end
				always @(posedge gclk or posedge reset)
					if (reset) begin
						glb_tile.if_cfg_est_m.rd_en <= 1'h0;
						glb_tile.if_cfg_est_m.rd_addr <= 12'h000;
					end
					else if (~(rd_tile_id_match && (glb_tile.if_cfg_wst_s.rd_en == 1'h1))) begin
						glb_tile.if_cfg_est_m.rd_en <= glb_tile.if_cfg_wst_s.rd_en;
						glb_tile.if_cfg_est_m.rd_addr <= glb_tile.if_cfg_wst_s.rd_addr;
					end
					else begin
						glb_tile.if_cfg_est_m.rd_en <= 1'h0;
						glb_tile.if_cfg_est_m.rd_addr <= 12'h000;
					end
				always @(posedge gclk or posedge reset)
					if (reset) begin
						glb_tile.if_cfg_wst_s.rd_data <= 32'h00000000;
						glb_tile.if_cfg_wst_s.rd_data_valid <= 1'h0;
					end
					else if (rd_data_valid_internal) begin
						glb_tile.if_cfg_wst_s.rd_data <= rd_data_internal;
						glb_tile.if_cfg_wst_s.rd_data_valid <= rd_data_valid_internal;
					end
					else begin
						glb_tile.if_cfg_wst_s.rd_data <= glb_tile.if_cfg_est_m.rd_data;
						glb_tile.if_cfg_wst_s.rd_data_valid <= glb_tile.if_cfg_est_m.rd_data_valid;
					end
				always @(posedge gclk or posedge reset)
					if (reset) begin
						rd_en_d1 <= 1'h0;
						rd_en_d2 <= 1'h0;
					end
					else begin
						rd_en_d1 <= read_internal;
						rd_en_d2 <= rd_en_d1;
					end
				always @(posedge gclk or posedge reset)
					if (reset) begin
						rd_data_valid_internal <= 1'h0;
						rd_data_internal <= 32'h00000000;
					end
					else if ((rd_en_d2 == 1'h1) & (d2h_dec_pio_ack | d2h_dec_pio_nack)) begin
						rd_data_valid_internal <= 1'h1;
						rd_data_internal <= d2h_dec_pio_read_data;
					end
					else begin
						rd_data_valid_internal <= 1'h0;
						rd_data_internal <= 32'h00000000;
					end
				always @(posedge mclk or posedge reset)
					if (reset) begin
						if_cfg_wst_s_wr_clk_en_d <= 1'h0;
						if_cfg_wst_s_rd_clk_en_d <= 1'h0;
					end
					else begin
						if_cfg_wst_s_wr_clk_en_d <= glb_tile.if_cfg_wst_s.wr_clk_en;
						if_cfg_wst_s_rd_clk_en_d <= glb_tile.if_cfg_wst_s.rd_clk_en;
					end
				always @(*) begin
					if_cfg_est_m_wr_clk_en_sel_first_cycle = glb_tile.if_cfg_wst_s.wr_en & ~wr_tile_id_match;
					if_cfg_est_m_rd_clk_en_sel_first_cycle = glb_tile.if_cfg_wst_s.rd_en & ~rd_tile_id_match;
				end
				always @(posedge mclk or posedge reset)
					if (reset)
						if_cfg_est_m_wr_clk_en_sel_latch <= 1'h0;
					else if (glb_tile.if_cfg_wst_s.wr_en == 1'h1) begin
						if (wr_tile_id_match)
							if_cfg_est_m_wr_clk_en_sel_latch <= 1'h0;
						else
							if_cfg_est_m_wr_clk_en_sel_latch <= 1'h1;
					end
					else if (glb_tile.if_cfg_wst_s.wr_clk_en == 1'h0)
						if_cfg_est_m_wr_clk_en_sel_latch <= 1'h0;
				always @(posedge mclk or posedge reset)
					if (reset)
						if_cfg_est_m_rd_clk_en_sel_latch <= 1'h0;
					else if (glb_tile.if_cfg_wst_s.rd_en == 1'h1) begin
						if (rd_tile_id_match)
							if_cfg_est_m_rd_clk_en_sel_latch <= 1'h0;
						else
							if_cfg_est_m_rd_clk_en_sel_latch <= 1'h1;
					end
					else if (glb_tile.if_cfg_wst_s.rd_clk_en == 1'h0)
						if_cfg_est_m_rd_clk_en_sel_latch <= 1'h0;
				always @(*) begin
					if_cfg_est_m_wr_clk_en_sel = if_cfg_est_m_wr_clk_en_sel_first_cycle | if_cfg_est_m_wr_clk_en_sel_latch;
					if_cfg_est_m_rd_clk_en_sel = if_cfg_est_m_rd_clk_en_sel_first_cycle | if_cfg_est_m_rd_clk_en_sel_latch;
				end
				always @(*)
					if (if_cfg_est_m_wr_clk_en_sel)
						glb_tile.if_cfg_est_m.wr_clk_en = if_cfg_wst_s_wr_clk_en_d;
					else
						glb_tile.if_cfg_est_m.wr_clk_en = 1'h0;
				always @(*)
					if (if_cfg_est_m_rd_clk_en_sel)
						glb_tile.if_cfg_est_m.rd_clk_en = if_cfg_wst_s_rd_clk_en_d;
					else
						glb_tile.if_cfg_est_m.rd_clk_en = 1'h0;
				assign h2d_pio_dec_write_data = wr_data_internal;
				assign h2d_pio_dec_address = addr_internal;
				assign h2d_pio_dec_read = read_internal;
				assign h2d_pio_dec_write = write_internal;
			end
			assign glb_cfg_ctrl.d2h_dec_pio_ack = glb_pio_d2h_dec_pio_ack;
			assign glb_cfg_ctrl.d2h_dec_pio_nack = glb_pio_d2h_dec_pio_nack;
			assign glb_cfg_ctrl.d2h_dec_pio_read_data = glb_pio_d2h_dec_pio_read_data;
			assign glb_cfg_ctrl.gclk = gclk;
			assign glb_cfg_ctrl.glb_tile_id = glb_tile_id;
			assign glb_cfg_ctrl.mclk = mclk;
			assign glb_cfg_ctrl.reset = reset;
			assign glb_cfg_ctrl_h2d_pio_dec_address = glb_cfg_ctrl.h2d_pio_dec_address;
			assign glb_pio_h2d_pio_dec_read = glb_cfg_ctrl.h2d_pio_dec_read;
			assign glb_pio_h2d_pio_dec_write = glb_cfg_ctrl.h2d_pio_dec_write;
			assign glb_pio_h2d_pio_dec_write_data = glb_cfg_ctrl.h2d_pio_dec_write_data;
		end
	endgenerate
	assign glb_cfg.gclk = gclk_cfg;
	assign glb_cfg.glb_tile_id = glb_tile_id;
	assign glb_cfg.mclk = clk;
	assign glb_cfg.reset = reset;
	assign glb_cfg_cfg_data_network = glb_cfg.cfg_data_network;
	assign cfg_ld_dma_ctrl = glb_cfg.cfg_ld_dma_ctrl;
	assign cfg_ld_dma_header = glb_cfg.cfg_ld_dma_header;
	assign cfg_pcfg_broadcast_mux = glb_cfg.cfg_pcfg_broadcast_mux;
	assign cfg_pcfg_dma_ctrl = glb_cfg.cfg_pcfg_dma_ctrl;
	assign cfg_pcfg_dma_header = glb_cfg.cfg_pcfg_dma_header;
	assign glb_cfg_cfg_pcfg_network = glb_cfg.cfg_pcfg_network;
	assign cfg_st_dma_ctrl = glb_cfg.cfg_st_dma_ctrl;
	assign cfg_st_dma_header = glb_cfg.cfg_st_dma_header;
	assign cfg_st_dma_num_blocks = glb_cfg.cfg_st_dma_num_blocks;
	glb_pcfg_broadcast glb_pcfg_broadcast(
		.cfg_pcfg_broadcast_mux(cfg_pcfg_broadcast_mux),
		.cgra_cfg_dma2mux(cgra_cfg_pcfgdma2mux),
		.cgra_cfg_jtag_addr_bypass_wsti(cgra_cfg_jtag_addr_bypass_wsti),
		.cgra_cfg_jtag_rd_en_bypass_wsti(cgra_cfg_jtag_rd_en_bypass_wsti),
		.cgra_cfg_jtag_wsti(glb_pcfg_broadcast_cgra_cfg_jtag_wsti),
		.cgra_cfg_pcfg_esti(glb_pcfg_broadcast_cgra_cfg_pcfg_esti),
		.cgra_cfg_pcfg_wsti(glb_pcfg_broadcast_cgra_cfg_pcfg_wsti),
		.clk(gclk_pcfg_broadcast),
		.reset(reset),
		.cgra_cfg_g2f(cgra_cfg_g2f_cfg_w),
		.cgra_cfg_jtag_addr_bypass_esto(cgra_cfg_jtag_addr_bypass_esto),
		.cgra_cfg_jtag_esto(glb_pcfg_broadcast_cgra_cfg_jtag_esto),
		.cgra_cfg_jtag_rd_en_bypass_esto(cgra_cfg_jtag_rd_en_bypass_esto),
		.cgra_cfg_pcfg_esto(glb_pcfg_broadcast_cgra_cfg_pcfg_esto),
		.cgra_cfg_pcfg_wsto(glb_pcfg_broadcast_cgra_cfg_pcfg_wsto)
	);
	glb_store_dma glb_store_dma(
		.cfg_data_network_f2g_mux(cfg_st_dma_ctrl[2-:2]),
		.cfg_data_network_latency(glb_cfg_cfg_data_network[5-:6]),
		.cfg_st_dma_ctrl_mode(cfg_st_dma_ctrl[6-:2]),
		.cfg_st_dma_ctrl_valid_mode(cfg_st_dma_ctrl[4-:2]),
		.cfg_st_dma_header(cfg_st_dma_header),
		.cfg_st_dma_num_blocks(cfg_st_dma_num_blocks),
		.cfg_st_dma_num_repeat(cfg_st_dma_ctrl[0]),
		.cfg_tile_connected_next(cfg_tile_connected_next),
		.cfg_tile_connected_prev(cfg_tile_connected_prev),
		.clk(gclk_st_dma),
		.ctrl_f2g(strm_ctrl_f2g),
		.data_f2g(strm_data_f2g),
		.data_f2g_vld(strm_data_f2g_vld),
		.reset(reset),
		.st_dma_start_pulse(strm_f2g_start_pulse),
		.clk_en_dma2bank(clk_en_stdma2bank),
		.data_f2g_rdy(strm_data_f2g_rdy),
		.st_dma_done_interrupt(strm_f2g_interrupt_pulse),
		.wr_packet_dma2bank(wr_packet_dma2bank),
		.wr_packet_dma2ring(wr_packet_dma2ring)
	);
	glb_load_dma glb_load_dma(
		.cfg_data_network_g2f_mux(cfg_ld_dma_ctrl[2-:2]),
		.cfg_data_network_latency(glb_cfg_cfg_data_network[5-:6]),
		.cfg_ld_dma_ctrl_flush_mode(cfg_ld_dma_ctrl[3]),
		.cfg_ld_dma_ctrl_mode(cfg_ld_dma_ctrl[7-:2]),
		.cfg_ld_dma_ctrl_valid_mode(cfg_ld_dma_ctrl[5-:2]),
		.cfg_ld_dma_header(cfg_ld_dma_header),
		.cfg_ld_dma_num_repeat(cfg_ld_dma_ctrl[0]),
		.cfg_tile_connected_next(cfg_tile_connected_next),
		.cfg_tile_connected_prev(cfg_tile_connected_prev),
		.clk(gclk_ld_dma),
		.data_g2f_rdy(strm_data_g2f_rdy),
		.glb_tile_id(glb_tile_id),
		.ld_dma_start_pulse(strm_g2f_start_pulse),
		.rdrs_packet_bank2dma(rdrs_packet_bank2dma),
		.rdrs_packet_ring2dma(rdrs_packet_ring2dma),
		.reset(reset),
		.clk_en_dma2bank(clk_en_lddma2bank),
		.ctrl_g2f(strm_ctrl_g2f),
		.data_flush(data_flush),
		.data_g2f(strm_data_g2f),
		.data_g2f_vld(strm_data_g2f_vld),
		.ld_dma_done_interrupt(strm_g2f_interrupt_pulse),
		.rdrq_packet_dma2bank(rdrq_packet_dma2bank),
		.rdrq_packet_dma2ring(rdrq_packet_dma2ring)
	);
	glb_pcfg_dma glb_pcfg_dma(
		.cfg_pcfg_dma_ctrl_mode(cfg_pcfg_dma_ctrl[17]),
		.cfg_pcfg_dma_ctrl_relocation_is_msb(cfg_pcfg_dma_ctrl[0]),
		.cfg_pcfg_dma_ctrl_relocation_value(cfg_pcfg_dma_ctrl[16-:16]),
		.cfg_pcfg_dma_header(cfg_pcfg_dma_header),
		.cfg_pcfg_network_latency(glb_cfg_cfg_pcfg_network[5-:6]),
		.cfg_pcfg_tile_connected_next(cfg_pcfg_tile_connected_next),
		.cfg_pcfg_tile_connected_prev(cfg_pcfg_tile_connected_prev),
		.clk(gclk_pcfg_dma),
		.glb_tile_id(glb_tile_id),
		.pcfg_dma_start_pulse(pcfg_start_pulse),
		.rdrs_packet_bank2dma(rdrs_packet_bank2pcfgdma),
		.rdrs_packet_ring2dma(rdrs_packet_pcfgring2dma),
		.reset(reset),
		.cgra_cfg_pcfg(cgra_cfg_pcfgdma2mux),
		.clk_en_dma2bank(clk_en_pcfgdma2bank),
		.pcfg_dma_done_interrupt(pcfg_g2f_interrupt_pulse),
		.rdrq_packet_dma2bank(rdrq_packet_pcfgdma2bank),
		.rdrq_packet_dma2ring(rdrq_packet_pcfgdma2ring)
	);
	glb_bank_mux glb_bank_mux(
		.cfg_pcfg_tile_connected_next(cfg_pcfg_tile_connected_next),
		.cfg_pcfg_tile_connected_prev(cfg_pcfg_tile_connected_prev),
		.cfg_tile_connected_next(cfg_tile_connected_next),
		.cfg_tile_connected_prev(cfg_tile_connected_prev),
		.clk(gclk_bank),
		.glb_tile_id(glb_tile_id),
		.rdrq_packet_dma2bank(rdrq_packet_dma2bank),
		.rdrq_packet_pcfgdma2bank(rdrq_packet_pcfgdma2bank),
		.rdrq_packet_pcfgring2bank(rdrq_packet_pcfgring2bank),
		.rdrq_packet_procsw2bank(rdrq_packet_procsw2bank),
		.rdrq_packet_ring2bank(rdrq_packet_ring2bank),
		.rdrs_packet_bankarr2sw(rdrs_packet_bankarr2sw),
		.reset(reset),
		.wr_packet_dma2bank(wr_packet_dma2bank),
		.wr_packet_procsw2bank(wr_packet_procsw2bank),
		.wr_packet_ring2bank(wr_packet_ring2bank),
		.rdrq_packet_sw2bankarr(rdrq_packet_sw2bankarr),
		.rdrs_packet_bank2dma(rdrs_packet_bank2dma),
		.rdrs_packet_bank2pcfgdma(rdrs_packet_bank2pcfgdma),
		.rdrs_packet_bank2pcfgring(rdrs_packet_bank2pcfgring),
		.rdrs_packet_bank2procsw(rdrs_packet_bank2procsw),
		.rdrs_packet_bank2ring(rdrs_packet_bank2ring),
		.wr_packet_sw2bankarr(wr_packet_sw2bankarr)
	);
	generate
		if (1) begin : glb_proc_switch
			wire gclk;
			wire glb_tile_id;
			wire mclk;
			wire [64:0] rdrs_packet;
			wire reset;
			wire clk_en_sw2bank;
			reg [19:0] rdrq_packet;
			reg [91:0] wr_packet;
			reg [18:0] bank_rd_addr;
			reg bank_rd_en;
			reg [18:0] bank_wr_addr;
			reg [63:0] bank_wr_data;
			reg bank_wr_en;
			reg [7:0] bank_wr_strb;
			reg [18:0] if_est_m_rd_addr_w;
			reg if_est_m_rd_clk_en_sel;
			reg if_est_m_rd_clk_en_sel_first_cycle;
			reg if_est_m_rd_clk_en_sel_latch;
			reg if_est_m_rd_en_w;
			reg [18:0] if_est_m_wr_addr_w;
			reg if_est_m_wr_clk_en_sel;
			reg if_est_m_wr_clk_en_sel_first_cycle;
			reg if_est_m_wr_clk_en_sel_latch;
			reg [63:0] if_est_m_wr_data_w;
			reg if_est_m_wr_en_w;
			reg [7:0] if_est_m_wr_strb_w;
			reg if_wst_s_rd_clk_en_d;
			reg if_wst_s_wr_clk_en_d;
			reg rd_data_valid_w;
			reg [63:0] rd_data_w;
			reg rd_tile_id_match;
			wire sw2bank_rd_clk_en;
			wire sw2bank_rd_clk_en_gen_enable;
			wire sw2bank_wr_clk_en;
			wire sw2bank_wr_clk_en_gen_enable;
			reg wr_tile_id_match;
			always @(*) begin
				wr_tile_id_match = glb_tile_id == glb_tile.if_proc_wst_s.wr_addr[18];
				rd_tile_id_match = glb_tile_id == glb_tile.if_proc_wst_s.rd_addr[18];
			end
			always @(*)
				if (glb_tile.if_proc_wst_s.wr_en) begin
					if (wr_tile_id_match) begin
						if_est_m_wr_en_w = 1'h0;
						if_est_m_wr_addr_w = 19'h00000;
						if_est_m_wr_data_w = 64'h0000000000000000;
						if_est_m_wr_strb_w = 8'h00;
						bank_wr_en = 1'h1;
						bank_wr_addr = glb_tile.if_proc_wst_s.wr_addr;
						bank_wr_data = glb_tile.if_proc_wst_s.wr_data;
						bank_wr_strb = glb_tile.if_proc_wst_s.wr_strb;
					end
					else begin
						if_est_m_wr_en_w = glb_tile.if_proc_wst_s.wr_en;
						if_est_m_wr_addr_w = glb_tile.if_proc_wst_s.wr_addr;
						if_est_m_wr_data_w = glb_tile.if_proc_wst_s.wr_data;
						if_est_m_wr_strb_w = glb_tile.if_proc_wst_s.wr_strb;
						bank_wr_en = 1'h0;
						bank_wr_addr = 19'h00000;
						bank_wr_data = 64'h0000000000000000;
						bank_wr_strb = 8'h00;
					end
				end
				else begin
					if_est_m_wr_en_w = 1'h0;
					if_est_m_wr_addr_w = 19'h00000;
					if_est_m_wr_data_w = 64'h0000000000000000;
					if_est_m_wr_strb_w = 8'h00;
					bank_wr_en = 1'h0;
					bank_wr_addr = 19'h00000;
					bank_wr_data = 64'h0000000000000000;
					bank_wr_strb = 8'h00;
				end
			always @(*)
				if (glb_tile.if_proc_wst_s.rd_en) begin
					if (rd_tile_id_match) begin
						if_est_m_rd_en_w = 1'h0;
						if_est_m_rd_addr_w = 19'h00000;
						bank_rd_en = 1'h1;
						bank_rd_addr = glb_tile.if_proc_wst_s.rd_addr;
					end
					else begin
						if_est_m_rd_en_w = glb_tile.if_proc_wst_s.rd_en;
						if_est_m_rd_addr_w = glb_tile.if_proc_wst_s.rd_addr;
						bank_rd_en = 1'h0;
						bank_rd_addr = 19'h00000;
					end
				end
				else begin
					if_est_m_rd_en_w = 1'h0;
					if_est_m_rd_addr_w = 19'h00000;
					bank_rd_en = 1'h0;
					bank_rd_addr = 19'h00000;
				end
			always @(*) begin
				rd_data_w = 64'h0000000000000000;
				rd_data_valid_w = 1'h0;
				if (rdrs_packet[0] == 1'h1) begin
					rd_data_w = rdrs_packet[64-:64];
					rd_data_valid_w = 1'h1;
				end
				else if (glb_tile.if_proc_est_m.rd_data_valid == 1'h1) begin
					rd_data_w = glb_tile.if_proc_est_m.rd_data;
					rd_data_valid_w = 1'h1;
				end
			end
			always @(posedge gclk or posedge reset)
				if (reset) begin
					glb_tile.if_proc_est_m.wr_en <= 1'h0;
					glb_tile.if_proc_est_m.wr_strb <= 8'h00;
					glb_tile.if_proc_est_m.wr_addr <= 19'h00000;
					glb_tile.if_proc_est_m.wr_data <= 64'h0000000000000000;
					glb_tile.if_proc_est_m.rd_en <= 1'h0;
					glb_tile.if_proc_est_m.rd_addr <= 19'h00000;
					glb_tile.if_proc_wst_s.rd_data <= 64'h0000000000000000;
					glb_tile.if_proc_wst_s.rd_data_valid <= 1'h0;
					wr_packet[91] <= 1'h0;
					wr_packet[90-:8] <= 8'h00;
					wr_packet[82-:19] <= 19'h00000;
					wr_packet[63-:64] <= 64'h0000000000000000;
					rdrq_packet[19] <= 1'h0;
					rdrq_packet[18-:19] <= 19'h00000;
				end
				else begin
					glb_tile.if_proc_est_m.wr_en <= if_est_m_wr_en_w;
					glb_tile.if_proc_est_m.wr_strb <= if_est_m_wr_strb_w;
					glb_tile.if_proc_est_m.wr_addr <= if_est_m_wr_addr_w;
					glb_tile.if_proc_est_m.wr_data <= if_est_m_wr_data_w;
					glb_tile.if_proc_est_m.rd_en <= if_est_m_rd_en_w;
					glb_tile.if_proc_est_m.rd_addr <= if_est_m_rd_addr_w;
					glb_tile.if_proc_wst_s.rd_data <= rd_data_w;
					glb_tile.if_proc_wst_s.rd_data_valid <= rd_data_valid_w;
					wr_packet[91] <= bank_wr_en;
					wr_packet[90-:8] <= bank_wr_strb;
					wr_packet[82-:19] <= bank_wr_addr;
					wr_packet[63-:64] <= bank_wr_data;
					rdrq_packet[19] <= bank_rd_en;
					rdrq_packet[18-:19] <= bank_rd_addr;
				end
			always @(posedge mclk or posedge reset)
				if (reset) begin
					if_wst_s_wr_clk_en_d <= 1'h0;
					if_wst_s_rd_clk_en_d <= 1'h0;
				end
				else begin
					if_wst_s_wr_clk_en_d <= glb_tile.if_proc_wst_s.wr_clk_en;
					if_wst_s_rd_clk_en_d <= glb_tile.if_proc_wst_s.rd_clk_en;
				end
			always @(*) begin
				if_est_m_wr_clk_en_sel_first_cycle = glb_tile.if_proc_wst_s.wr_en & ~wr_tile_id_match;
				if_est_m_rd_clk_en_sel_first_cycle = glb_tile.if_proc_wst_s.rd_en & ~rd_tile_id_match;
			end
			always @(posedge mclk or posedge reset)
				if (reset)
					if_est_m_wr_clk_en_sel_latch <= 1'h0;
				else if (glb_tile.if_proc_wst_s.wr_en == 1'h1) begin
					if (wr_tile_id_match)
						if_est_m_wr_clk_en_sel_latch <= 1'h0;
					else
						if_est_m_wr_clk_en_sel_latch <= 1'h1;
				end
				else if (glb_tile.if_proc_wst_s.wr_clk_en == 1'h0)
					if_est_m_wr_clk_en_sel_latch <= 1'h0;
			always @(posedge mclk or posedge reset)
				if (reset)
					if_est_m_rd_clk_en_sel_latch <= 1'h0;
				else if (glb_tile.if_proc_wst_s.rd_en == 1'h1) begin
					if (rd_tile_id_match)
						if_est_m_rd_clk_en_sel_latch <= 1'h0;
					else
						if_est_m_rd_clk_en_sel_latch <= 1'h1;
				end
				else if (glb_tile.if_proc_wst_s.rd_clk_en == 1'h0)
					if_est_m_rd_clk_en_sel_latch <= 1'h0;
			always @(*) begin
				if_est_m_wr_clk_en_sel = if_est_m_wr_clk_en_sel_first_cycle | if_est_m_wr_clk_en_sel_latch;
				if_est_m_rd_clk_en_sel = if_est_m_rd_clk_en_sel_first_cycle | if_est_m_rd_clk_en_sel_latch;
			end
			always @(*)
				if (if_est_m_wr_clk_en_sel)
					glb_tile.if_proc_est_m.wr_clk_en = if_wst_s_wr_clk_en_d;
				else
					glb_tile.if_proc_est_m.wr_clk_en = 1'h0;
			always @(*)
				if (if_est_m_rd_clk_en_sel)
					glb_tile.if_proc_est_m.rd_clk_en = if_wst_s_rd_clk_en_d;
				else
					glb_tile.if_proc_est_m.rd_clk_en = 1'h0;
			assign sw2bank_wr_clk_en_gen_enable = glb_tile.if_proc_wst_s.wr_en & wr_tile_id_match;
			assign sw2bank_rd_clk_en_gen_enable = glb_tile.if_proc_wst_s.rd_en & rd_tile_id_match;
			assign clk_en_sw2bank = sw2bank_wr_clk_en | sw2bank_rd_clk_en;
			glb_clk_en_gen_4 #(.cnt(32'h00000004)) sw2bank_wr_clk_en_gen(
				.clk(mclk),
				.enable(sw2bank_wr_clk_en_gen_enable),
				.reset(reset),
				.clk_en(sw2bank_wr_clk_en)
			);
			glb_clk_en_gen_6 #(.cnt(32'h00000006)) sw2bank_rd_clk_en_gen(
				.clk(mclk),
				.enable(sw2bank_rd_clk_en_gen_enable),
				.reset(reset),
				.clk_en(sw2bank_rd_clk_en)
			);
		end
	endgenerate
	assign glb_proc_switch.gclk = gclk_proc_switch;
	assign glb_proc_switch.glb_tile_id = glb_tile_id;
	assign glb_proc_switch.mclk = clk;
	assign glb_proc_switch.rdrs_packet = rdrs_packet_bank2procsw;
	assign glb_proc_switch.reset = reset;
	assign clk_en_procsw2bank = glb_proc_switch.clk_en_sw2bank;
	assign rdrq_packet_procsw2bank = glb_proc_switch.rdrq_packet;
	assign wr_packet_procsw2bank = glb_proc_switch.wr_packet;
	glb_ring_switch_WR_RD glb_strm_ring_switch(
		.cfg_ld_dma_on(glb_strm_ring_switch_cfg_ld_dma_on),
		.cfg_tile_connected_next(cfg_tile_connected_next),
		.cfg_tile_connected_prev(cfg_tile_connected_prev),
		.clk(gclk_strm_switch),
		.glb_tile_id(glb_tile_id),
		.rdrq_packet_dma2ring(rdrq_packet_dma2ring),
		.rdrq_packet_e2w_esti(strm_rdrq_packet_e2w_esti),
		.rdrq_packet_w2e_wsti(strm_rdrq_packet_w2e_wsti),
		.rdrs_packet_bank2ring(rdrs_packet_bank2ring),
		.rdrs_packet_e2w_esti(strm_rdrs_packet_e2w_esti),
		.rdrs_packet_w2e_wsti(strm_rdrs_packet_w2e_wsti),
		.reset(reset),
		.wr_packet_dma2ring(wr_packet_dma2ring),
		.wr_packet_e2w_esti(strm_wr_packet_e2w_esti),
		.wr_packet_w2e_wsti(strm_wr_packet_w2e_wsti),
		.clk_en_ring2bank(clk_en_ring2bank),
		.rdrq_packet_e2w_wsto(strm_rdrq_packet_e2w_wsto),
		.rdrq_packet_ring2bank(rdrq_packet_ring2bank),
		.rdrq_packet_w2e_esto(strm_rdrq_packet_w2e_esto),
		.rdrs_packet_e2w_wsto(strm_rdrs_packet_e2w_wsto),
		.rdrs_packet_ring2dma(rdrs_packet_ring2dma),
		.rdrs_packet_w2e_esto(strm_rdrs_packet_w2e_esto),
		.wr_packet_e2w_wsto(strm_wr_packet_e2w_wsto),
		.wr_packet_ring2bank(wr_packet_ring2bank),
		.wr_packet_w2e_esto(strm_wr_packet_w2e_esto)
	);
	glb_ring_switch_RD glb_pcfg_ring_switch(
		.cfg_ld_dma_on(glb_pcfg_ring_switch_cfg_ld_dma_on),
		.cfg_tile_connected_next(cfg_pcfg_tile_connected_next),
		.cfg_tile_connected_prev(cfg_pcfg_tile_connected_prev),
		.clk(gclk_pcfg_switch),
		.glb_tile_id(glb_tile_id),
		.rdrq_packet_dma2ring(rdrq_packet_pcfgdma2ring),
		.rdrq_packet_e2w_esti(pcfg_rdrq_packet_e2w_esti),
		.rdrq_packet_w2e_wsti(pcfg_rdrq_packet_w2e_wsti),
		.rdrs_packet_bank2ring(rdrs_packet_bank2pcfgring),
		.rdrs_packet_e2w_esti(pcfg_rdrs_packet_e2w_esti),
		.rdrs_packet_w2e_wsti(pcfg_rdrs_packet_w2e_wsti),
		.reset(reset),
		.clk_en_ring2bank(clk_en_pcfgring2bank),
		.rdrq_packet_e2w_wsto(pcfg_rdrq_packet_e2w_wsto),
		.rdrq_packet_ring2bank(rdrq_packet_pcfgring2bank),
		.rdrq_packet_w2e_esto(pcfg_rdrq_packet_w2e_esto),
		.rdrs_packet_e2w_wsto(pcfg_rdrs_packet_e2w_wsto),
		.rdrs_packet_ring2dma(rdrs_packet_pcfgring2dma),
		.rdrs_packet_w2e_esto(pcfg_rdrs_packet_w2e_esto)
	);
	glb_bank glb_bank_0(
		.clk(gclk_bank),
		.rdrq_packet(rdrq_packet_sw2bankarr[0+:18]),
		.reset(reset),
		.wr_packet(wr_packet_sw2bankarr[0+:90]),
		.rdrs_packet(glb_bank_0_rdrs_packet)
	);
	glb_bank glb_bank_1(
		.clk(gclk_bank),
		.rdrq_packet(rdrq_packet_sw2bankarr[18+:18]),
		.reset(reset),
		.wr_packet(wr_packet_sw2bankarr[90+:90]),
		.rdrs_packet(glb_bank_1_rdrs_packet)
	);
endmodule
module global_buffer (
	cgra_cfg_jtag_gc2glb_addr,
	cgra_cfg_jtag_gc2glb_data,
	cgra_cfg_jtag_gc2glb_rd_en,
	cgra_cfg_jtag_gc2glb_wr_en,
	cgra_stall_in,
	clk,
	flush_crossbar_sel,
	glb_clk_en_bank_master,
	glb_clk_en_master,
	if_cfg_rd_addr,
	if_cfg_rd_clk_en,
	if_cfg_rd_en,
	if_cfg_wr_addr,
	if_cfg_wr_clk_en,
	if_cfg_wr_data,
	if_cfg_wr_en,
	if_sram_cfg_rd_addr,
	if_sram_cfg_rd_en,
	if_sram_cfg_wr_addr,
	if_sram_cfg_wr_data,
	if_sram_cfg_wr_en,
	pcfg_broadcast_stall,
	pcfg_start_pulse,
	proc_rd_addr,
	proc_rd_en,
	proc_wr_addr,
	proc_wr_data,
	proc_wr_en,
	proc_wr_strb,
	reset,
	strm_ctrl_f2g,
	strm_data_f2g,
	strm_data_f2g_vld,
	strm_data_g2f_rdy,
	strm_f2g_start_pulse,
	strm_g2f_start_pulse,
	cgra_cfg_g2f_cfg_addr,
	cgra_cfg_g2f_cfg_data,
	cgra_cfg_g2f_cfg_rd_en,
	cgra_cfg_g2f_cfg_wr_en,
	cgra_stall,
	if_cfg_rd_data,
	if_cfg_rd_data_valid,
	if_sram_cfg_rd_data,
	if_sram_cfg_rd_data_valid,
	pcfg_g2f_interrupt_pulse,
	proc_rd_data,
	proc_rd_data_valid,
	strm_ctrl_g2f,
	strm_data_f2g_rdy,
	strm_data_flush_g2f,
	strm_data_g2f,
	strm_data_g2f_vld,
	strm_f2g_interrupt_pulse,
	strm_g2f_interrupt_pulse
);
	input wire [31:0] cgra_cfg_jtag_gc2glb_addr;
	input wire [31:0] cgra_cfg_jtag_gc2glb_data;
	input wire cgra_cfg_jtag_gc2glb_rd_en;
	input wire cgra_cfg_jtag_gc2glb_wr_en;
	input wire [3:0] cgra_stall_in;
	input wire clk;
	input wire flush_crossbar_sel;
	input wire [1:0] glb_clk_en_bank_master;
	input wire [1:0] glb_clk_en_master;
	input wire [11:0] if_cfg_rd_addr;
	input wire if_cfg_rd_clk_en;
	input wire if_cfg_rd_en;
	input wire [11:0] if_cfg_wr_addr;
	input wire if_cfg_wr_clk_en;
	input wire [31:0] if_cfg_wr_data;
	input wire if_cfg_wr_en;
	input wire [18:0] if_sram_cfg_rd_addr;
	input wire if_sram_cfg_rd_en;
	input wire [18:0] if_sram_cfg_wr_addr;
	input wire [31:0] if_sram_cfg_wr_data;
	input wire if_sram_cfg_wr_en;
	input wire [1:0] pcfg_broadcast_stall;
	input wire [1:0] pcfg_start_pulse;
	input wire [18:0] proc_rd_addr;
	input wire proc_rd_en;
	input wire [18:0] proc_wr_addr;
	input wire [63:0] proc_wr_data;
	input wire proc_wr_en;
	input wire [7:0] proc_wr_strb;
	input wire reset;
	input wire [3:0] strm_ctrl_f2g;
	input wire [63:0] strm_data_f2g;
	input wire [3:0] strm_data_f2g_vld;
	input wire [3:0] strm_data_g2f_rdy;
	input wire [1:0] strm_f2g_start_pulse;
	input wire [1:0] strm_g2f_start_pulse;
	output wire [127:0] cgra_cfg_g2f_cfg_addr;
	output wire [127:0] cgra_cfg_g2f_cfg_data;
	output wire [3:0] cgra_cfg_g2f_cfg_rd_en;
	output wire [3:0] cgra_cfg_g2f_cfg_wr_en;
	output wire [3:0] cgra_stall;
	output wire [31:0] if_cfg_rd_data;
	output wire if_cfg_rd_data_valid;
	output reg [31:0] if_sram_cfg_rd_data;
	output reg if_sram_cfg_rd_data_valid;
	output wire [1:0] pcfg_g2f_interrupt_pulse;
	output reg [63:0] proc_rd_data;
	output reg proc_rd_data_valid;
	output wire [3:0] strm_ctrl_g2f;
	output wire [3:0] strm_data_f2g_rdy;
	output wire strm_data_flush_g2f;
	output wire [63:0] strm_data_g2f;
	output wire [3:0] strm_data_g2f_vld;
	output wire [1:0] strm_f2g_interrupt_pulse;
	output wire [1:0] strm_g2f_interrupt_pulse;
	wire [2:0] cfg_pcfg_tile_connected;
	wire [2:0] cfg_tile_connected;
	wire [63:0] cgra_cfg_jtag_addr_bypass_esto;
	reg [63:0] cgra_cfg_jtag_addr_bypass_wsti;
	wire [63:0] cgra_cfg_jtag_addr_esto;
	reg [63:0] cgra_cfg_jtag_addr_wsti;
	wire [63:0] cgra_cfg_jtag_data_esto;
	reg [63:0] cgra_cfg_jtag_data_wsti;
	reg [31:0] cgra_cfg_jtag_gc2glb_addr_d;
	reg [31:0] cgra_cfg_jtag_gc2glb_data_d;
	reg cgra_cfg_jtag_gc2glb_rd_en_d;
	reg cgra_cfg_jtag_gc2glb_wr_en_d;
	wire [1:0] cgra_cfg_jtag_rd_en_bypass_esto;
	reg [1:0] cgra_cfg_jtag_rd_en_bypass_wsti;
	wire [1:0] cgra_cfg_jtag_rd_en_esto;
	reg [1:0] cgra_cfg_jtag_rd_en_wsti;
	wire [1:0] cgra_cfg_jtag_wr_en_esto;
	reg [1:0] cgra_cfg_jtag_wr_en_wsti;
	reg [63:0] cgra_cfg_pcfg_addr_esti;
	wire [63:0] cgra_cfg_pcfg_addr_esto;
	reg [63:0] cgra_cfg_pcfg_addr_wsti;
	wire [63:0] cgra_cfg_pcfg_addr_wsto;
	reg [63:0] cgra_cfg_pcfg_data_esti;
	wire [63:0] cgra_cfg_pcfg_data_esto;
	reg [63:0] cgra_cfg_pcfg_data_wsti;
	wire [63:0] cgra_cfg_pcfg_data_wsto;
	reg [1:0] cgra_cfg_pcfg_rd_en_esti;
	wire [1:0] cgra_cfg_pcfg_rd_en_esto;
	reg [1:0] cgra_cfg_pcfg_rd_en_wsti;
	wire [1:0] cgra_cfg_pcfg_rd_en_wsto;
	reg [1:0] cgra_cfg_pcfg_wr_en_esti;
	wire [1:0] cgra_cfg_pcfg_wr_en_esto;
	reg [1:0] cgra_cfg_pcfg_wr_en_wsti;
	wire [1:0] cgra_cfg_pcfg_wr_en_wsto;
	wire [1:0] data_flush;
	wire [1:0] data_flush_d;
	wire [1:0] flush_crossbar_in;
	wire flush_crossbar_sel_w;
	wire glb_tile_gen_0_cfg_pcfg_tile_connected_esto;
	wire glb_tile_gen_0_cfg_tile_connected_esto;
	wire [63:0] glb_tile_gen_0_cgra_cfg_g2f_cfg_addr;
	wire [63:0] glb_tile_gen_0_cgra_cfg_g2f_cfg_data;
	wire [1:0] glb_tile_gen_0_cgra_cfg_g2f_cfg_rd_en;
	wire [1:0] glb_tile_gen_0_cgra_cfg_g2f_cfg_wr_en;
	wire [31:0] glb_tile_gen_0_cgra_cfg_jtag_addr_bypass_esto;
	wire [31:0] glb_tile_gen_0_cgra_cfg_jtag_addr_esto;
	wire [31:0] glb_tile_gen_0_cgra_cfg_jtag_data_esto;
	wire glb_tile_gen_0_cgra_cfg_jtag_rd_en_bypass_esto;
	wire glb_tile_gen_0_cgra_cfg_jtag_rd_en_esto;
	wire glb_tile_gen_0_cgra_cfg_jtag_wr_en_esto;
	wire [31:0] glb_tile_gen_0_cgra_cfg_pcfg_addr_e2w_wsto;
	wire [31:0] glb_tile_gen_0_cgra_cfg_pcfg_addr_w2e_esto;
	wire [31:0] glb_tile_gen_0_cgra_cfg_pcfg_data_e2w_wsto;
	wire [31:0] glb_tile_gen_0_cgra_cfg_pcfg_data_w2e_esto;
	wire glb_tile_gen_0_cgra_cfg_pcfg_rd_en_e2w_wsto;
	wire glb_tile_gen_0_cgra_cfg_pcfg_rd_en_w2e_esto;
	wire glb_tile_gen_0_cgra_cfg_pcfg_wr_en_e2w_wsto;
	wire glb_tile_gen_0_cgra_cfg_pcfg_wr_en_w2e_esto;
	wire glb_tile_gen_0_clk_en_bank_master;
	wire glb_tile_gen_0_clk_en_master;
	wire glb_tile_gen_0_clk_en_pcfg_broadcast;
	wire glb_tile_gen_0_data_flush;
	wire glb_tile_gen_0_pcfg_g2f_interrupt_pulse;
	wire [18:0] glb_tile_gen_0_pcfg_rd_addr_e2w_wsto;
	wire [18:0] glb_tile_gen_0_pcfg_rd_addr_w2e_esto;
	wire [63:0] glb_tile_gen_0_pcfg_rd_data_e2w_wsto;
	wire glb_tile_gen_0_pcfg_rd_data_valid_e2w_wsto;
	wire glb_tile_gen_0_pcfg_rd_data_valid_w2e_esto;
	wire [63:0] glb_tile_gen_0_pcfg_rd_data_w2e_esto;
	wire glb_tile_gen_0_pcfg_rd_en_e2w_wsto;
	wire glb_tile_gen_0_pcfg_rd_en_w2e_esto;
	wire [1:0] glb_tile_gen_0_strm_ctrl_g2f;
	wire [1:0] glb_tile_gen_0_strm_data_f2g_rdy;
	wire [31:0] glb_tile_gen_0_strm_data_g2f;
	wire [1:0] glb_tile_gen_0_strm_data_g2f_vld;
	wire glb_tile_gen_0_strm_f2g_interrupt_pulse;
	wire glb_tile_gen_0_strm_g2f_interrupt_pulse;
	wire [18:0] glb_tile_gen_0_strm_rd_addr_e2w_wsto;
	wire [18:0] glb_tile_gen_0_strm_rd_addr_w2e_esto;
	wire [63:0] glb_tile_gen_0_strm_rd_data_e2w_wsto;
	wire glb_tile_gen_0_strm_rd_data_valid_e2w_wsto;
	wire glb_tile_gen_0_strm_rd_data_valid_w2e_esto;
	wire [63:0] glb_tile_gen_0_strm_rd_data_w2e_esto;
	wire glb_tile_gen_0_strm_rd_en_e2w_wsto;
	wire glb_tile_gen_0_strm_rd_en_w2e_esto;
	wire [18:0] glb_tile_gen_0_strm_wr_addr_e2w_wsto;
	wire [18:0] glb_tile_gen_0_strm_wr_addr_w2e_esto;
	wire [63:0] glb_tile_gen_0_strm_wr_data_e2w_wsto;
	wire [63:0] glb_tile_gen_0_strm_wr_data_w2e_esto;
	wire glb_tile_gen_0_strm_wr_en_e2w_wsto;
	wire glb_tile_gen_0_strm_wr_en_w2e_esto;
	wire [7:0] glb_tile_gen_0_strm_wr_strb_e2w_wsto;
	wire [7:0] glb_tile_gen_0_strm_wr_strb_w2e_esto;
	wire glb_tile_gen_1_cfg_pcfg_tile_connected_esto;
	wire glb_tile_gen_1_cfg_tile_connected_esto;
	wire [63:0] glb_tile_gen_1_cgra_cfg_g2f_cfg_addr;
	wire [63:0] glb_tile_gen_1_cgra_cfg_g2f_cfg_data;
	wire [1:0] glb_tile_gen_1_cgra_cfg_g2f_cfg_rd_en;
	wire [1:0] glb_tile_gen_1_cgra_cfg_g2f_cfg_wr_en;
	wire [31:0] glb_tile_gen_1_cgra_cfg_jtag_addr_bypass_esto;
	wire [31:0] glb_tile_gen_1_cgra_cfg_jtag_addr_esto;
	wire [31:0] glb_tile_gen_1_cgra_cfg_jtag_data_esto;
	wire glb_tile_gen_1_cgra_cfg_jtag_rd_en_bypass_esto;
	wire glb_tile_gen_1_cgra_cfg_jtag_rd_en_esto;
	wire glb_tile_gen_1_cgra_cfg_jtag_wr_en_esto;
	wire [31:0] glb_tile_gen_1_cgra_cfg_pcfg_addr_e2w_wsto;
	wire [31:0] glb_tile_gen_1_cgra_cfg_pcfg_addr_w2e_esto;
	wire [31:0] glb_tile_gen_1_cgra_cfg_pcfg_data_e2w_wsto;
	wire [31:0] glb_tile_gen_1_cgra_cfg_pcfg_data_w2e_esto;
	wire glb_tile_gen_1_cgra_cfg_pcfg_rd_en_e2w_wsto;
	wire glb_tile_gen_1_cgra_cfg_pcfg_rd_en_w2e_esto;
	wire glb_tile_gen_1_cgra_cfg_pcfg_wr_en_e2w_wsto;
	wire glb_tile_gen_1_cgra_cfg_pcfg_wr_en_w2e_esto;
	wire glb_tile_gen_1_clk_en_bank_master;
	wire glb_tile_gen_1_clk_en_master;
	wire glb_tile_gen_1_clk_en_pcfg_broadcast;
	wire glb_tile_gen_1_data_flush;
	wire glb_tile_gen_1_pcfg_g2f_interrupt_pulse;
	wire [18:0] glb_tile_gen_1_pcfg_rd_addr_e2w_wsto;
	wire [18:0] glb_tile_gen_1_pcfg_rd_addr_w2e_esto;
	wire [63:0] glb_tile_gen_1_pcfg_rd_data_e2w_wsto;
	wire glb_tile_gen_1_pcfg_rd_data_valid_e2w_wsto;
	wire glb_tile_gen_1_pcfg_rd_data_valid_w2e_esto;
	wire [63:0] glb_tile_gen_1_pcfg_rd_data_w2e_esto;
	wire glb_tile_gen_1_pcfg_rd_en_e2w_wsto;
	wire glb_tile_gen_1_pcfg_rd_en_w2e_esto;
	wire [1:0] glb_tile_gen_1_strm_ctrl_g2f;
	wire [1:0] glb_tile_gen_1_strm_data_f2g_rdy;
	wire [31:0] glb_tile_gen_1_strm_data_g2f;
	wire [1:0] glb_tile_gen_1_strm_data_g2f_vld;
	wire glb_tile_gen_1_strm_f2g_interrupt_pulse;
	wire glb_tile_gen_1_strm_g2f_interrupt_pulse;
	wire [18:0] glb_tile_gen_1_strm_rd_addr_e2w_wsto;
	wire [18:0] glb_tile_gen_1_strm_rd_addr_w2e_esto;
	wire [63:0] glb_tile_gen_1_strm_rd_data_e2w_wsto;
	wire glb_tile_gen_1_strm_rd_data_valid_e2w_wsto;
	wire glb_tile_gen_1_strm_rd_data_valid_w2e_esto;
	wire [63:0] glb_tile_gen_1_strm_rd_data_w2e_esto;
	wire glb_tile_gen_1_strm_rd_en_e2w_wsto;
	wire glb_tile_gen_1_strm_rd_en_w2e_esto;
	wire [18:0] glb_tile_gen_1_strm_wr_addr_e2w_wsto;
	wire [18:0] glb_tile_gen_1_strm_wr_addr_w2e_esto;
	wire [63:0] glb_tile_gen_1_strm_wr_data_e2w_wsto;
	wire [63:0] glb_tile_gen_1_strm_wr_data_w2e_esto;
	wire glb_tile_gen_1_strm_wr_en_e2w_wsto;
	wire glb_tile_gen_1_strm_wr_en_w2e_esto;
	wire [7:0] glb_tile_gen_1_strm_wr_strb_e2w_wsto;
	wire [7:0] glb_tile_gen_1_strm_wr_strb_w2e_esto;
	reg if_sram_cfg_rd_data_valid_w;
	reg [31:0] if_sram_cfg_rd_data_w;
	reg [1:0] pcfg_g2f_interrupt_pulse_d;
	wire [1:0] pcfg_g2f_interrupt_pulse_w;
	wire [169:0] pcfg_packet_e2w_esti;
	wire [169:0] pcfg_packet_e2w_wsto;
	wire [169:0] pcfg_packet_w2e_esto;
	wire [169:0] pcfg_packet_w2e_wsti;
	reg [18:0] proc_rd_addr_d;
	reg proc_rd_addr_sel;
	wire proc_rd_clk_en;
	wire proc_rd_clk_en_gen_enable;
	reg proc_rd_data_valid_w;
	reg [63:0] proc_rd_data_w;
	reg proc_rd_en_d;
	reg proc_rd_type;
	reg [18:0] proc_wr_addr_d;
	wire proc_wr_clk_en;
	wire proc_wr_clk_en_gen_enable;
	reg [63:0] proc_wr_data_d;
	reg proc_wr_en_d;
	reg [7:0] proc_wr_strb_d;
	reg [18:0] sram_cfg_rd_addr_d;
	reg sram_cfg_rd_en_d;
	reg [18:0] sram_cfg_wr_addr_d;
	reg [63:0] sram_cfg_wr_data_d;
	reg sram_cfg_wr_en_d;
	reg [7:0] sram_cfg_wr_strb_d;
	reg [1:0] strm_f2g_interrupt_pulse_d;
	wire [1:0] strm_f2g_interrupt_pulse_w;
	reg [1:0] strm_g2f_interrupt_pulse_d;
	wire [1:0] strm_g2f_interrupt_pulse_w;
	wire [353:0] strm_packet_e2w_esti;
	wire [353:0] strm_packet_e2w_wsto;
	wire [353:0] strm_packet_w2e_esto;
	wire [353:0] strm_packet_w2e_wsti;
	generate
		if (1) begin : if_cfg_tile2tile_0
			reg [11:0] rd_addr;
			reg rd_clk_en;
			wire [31:0] rd_data;
			wire rd_data_valid;
			reg rd_en;
			reg [11:0] wr_addr;
			reg wr_clk_en;
			reg [31:0] wr_data;
			reg wr_en;
		end
		if (1) begin : if_cfg_tile2tile_1
			wire [11:0] rd_addr;
			wire rd_clk_en;
			wire [31:0] rd_data;
			wire rd_data_valid;
			wire rd_en;
			wire [11:0] wr_addr;
			wire wr_clk_en;
			wire [31:0] wr_data;
			wire wr_en;
		end
		if (1) begin : if_cfg_tile2tile_2
			wire [11:0] rd_addr;
			wire rd_clk_en;
			wire [31:0] rd_data;
			wire rd_data_valid;
			wire rd_en;
			wire [11:0] wr_addr;
			wire wr_clk_en;
			wire [31:0] wr_data;
			wire wr_en;
		end
		if (1) begin : if_proc_tile2tile_0
			reg [18:0] rd_addr;
			wire rd_clk_en;
			wire [63:0] rd_data;
			wire rd_data_valid;
			reg rd_en;
			reg [18:0] wr_addr;
			wire wr_clk_en;
			reg [63:0] wr_data;
			reg wr_en;
			reg [7:0] wr_strb;
		end
		if (1) begin : if_proc_tile2tile_1
			wire [18:0] rd_addr;
			wire rd_clk_en;
			wire [63:0] rd_data;
			wire rd_data_valid;
			wire rd_en;
			wire [18:0] wr_addr;
			wire wr_clk_en;
			wire [63:0] wr_data;
			wire wr_en;
			wire [7:0] wr_strb;
		end
		if (1) begin : if_proc_tile2tile_2
			wire [18:0] rd_addr;
			wire rd_clk_en;
			wire [63:0] rd_data;
			wire rd_data_valid;
			wire rd_en;
			wire [18:0] wr_addr;
			wire wr_clk_en;
			wire [63:0] wr_data;
			wire wr_en;
			wire [7:0] wr_strb;
		end
		if (1) begin : if_sram_cfg_tile2tile_0
			wire [18:0] rd_addr;
			wire rd_clk_en;
			wire [31:0] rd_data;
			wire rd_data_valid;
			wire rd_en;
			wire [18:0] wr_addr;
			wire wr_clk_en;
			wire [31:0] wr_data;
			wire wr_en;
		end
		if (1) begin : if_sram_cfg_tile2tile_1
			wire [18:0] rd_addr;
			wire rd_clk_en;
			wire [31:0] rd_data;
			wire rd_data_valid;
			wire rd_en;
			wire [18:0] wr_addr;
			wire wr_clk_en;
			wire [31:0] wr_data;
			wire wr_en;
		end
		if (1) begin : if_sram_cfg_tile2tile_2
			wire [18:0] rd_addr;
			wire rd_clk_en;
			wire [31:0] rd_data;
			wire rd_data_valid;
			wire rd_en;
			wire [18:0] wr_addr;
			wire wr_clk_en;
			wire [31:0] wr_data;
			wire wr_en;
		end
	endgenerate
	assign cfg_tile_connected[0] = 1'h0;
	assign cfg_pcfg_tile_connected[0] = 1'h0;
	assign strm_f2g_interrupt_pulse = strm_f2g_interrupt_pulse_d;
	assign strm_g2f_interrupt_pulse = strm_g2f_interrupt_pulse_d;
	assign pcfg_g2f_interrupt_pulse = pcfg_g2f_interrupt_pulse_d;
	assign cgra_stall = cgra_stall_in;
	assign if_sram_cfg_tile2tile_2.rd_data = 32'h00000000;
	assign if_sram_cfg_tile2tile_2.rd_data_valid = 1'h0;
	assign glb_tile_gen_0_clk_en_pcfg_broadcast = ~pcfg_broadcast_stall[0];
	assign glb_tile_gen_0_clk_en_master = glb_clk_en_master[0];
	assign glb_tile_gen_0_clk_en_bank_master = glb_clk_en_bank_master[0];
	assign strm_packet_w2e_esto[176] = glb_tile_gen_0_strm_wr_en_w2e_esto;
	assign strm_packet_w2e_esto[175-:8] = glb_tile_gen_0_strm_wr_strb_w2e_esto;
	assign strm_packet_w2e_esto[167-:19] = glb_tile_gen_0_strm_wr_addr_w2e_esto;
	assign strm_packet_w2e_esto[148-:64] = glb_tile_gen_0_strm_wr_data_w2e_esto;
	assign strm_packet_w2e_esto[84] = glb_tile_gen_0_strm_rd_en_w2e_esto;
	assign strm_packet_w2e_esto[83-:19] = glb_tile_gen_0_strm_rd_addr_w2e_esto;
	assign strm_packet_w2e_esto[64-:64] = glb_tile_gen_0_strm_rd_data_w2e_esto;
	assign strm_packet_w2e_esto[0] = glb_tile_gen_0_strm_rd_data_valid_w2e_esto;
	assign strm_packet_e2w_wsto[176] = glb_tile_gen_0_strm_wr_en_e2w_wsto;
	assign strm_packet_e2w_wsto[175-:8] = glb_tile_gen_0_strm_wr_strb_e2w_wsto;
	assign strm_packet_e2w_wsto[167-:19] = glb_tile_gen_0_strm_wr_addr_e2w_wsto;
	assign strm_packet_e2w_wsto[148-:64] = glb_tile_gen_0_strm_wr_data_e2w_wsto;
	assign strm_packet_e2w_wsto[84] = glb_tile_gen_0_strm_rd_en_e2w_wsto;
	assign strm_packet_e2w_wsto[83-:19] = glb_tile_gen_0_strm_rd_addr_e2w_wsto;
	assign strm_packet_e2w_wsto[64-:64] = glb_tile_gen_0_strm_rd_data_e2w_wsto;
	assign strm_packet_e2w_wsto[0] = glb_tile_gen_0_strm_rd_data_valid_e2w_wsto;
	assign pcfg_packet_w2e_esto[84] = glb_tile_gen_0_pcfg_rd_en_w2e_esto;
	assign pcfg_packet_w2e_esto[83-:19] = glb_tile_gen_0_pcfg_rd_addr_w2e_esto;
	assign pcfg_packet_w2e_esto[64-:64] = glb_tile_gen_0_pcfg_rd_data_w2e_esto;
	assign pcfg_packet_w2e_esto[0] = glb_tile_gen_0_pcfg_rd_data_valid_w2e_esto;
	assign pcfg_packet_e2w_wsto[84] = glb_tile_gen_0_pcfg_rd_en_e2w_wsto;
	assign pcfg_packet_e2w_wsto[83-:19] = glb_tile_gen_0_pcfg_rd_addr_e2w_wsto;
	assign pcfg_packet_e2w_wsto[64-:64] = glb_tile_gen_0_pcfg_rd_data_e2w_wsto;
	assign pcfg_packet_e2w_wsto[0] = glb_tile_gen_0_pcfg_rd_data_valid_e2w_wsto;
	assign cfg_tile_connected[1] = glb_tile_gen_0_cfg_tile_connected_esto;
	assign cfg_pcfg_tile_connected[1] = glb_tile_gen_0_cfg_pcfg_tile_connected_esto;
	assign strm_data_f2g_rdy[0+:2] = glb_tile_gen_0_strm_data_f2g_rdy;
	assign strm_data_g2f[0+:32] = glb_tile_gen_0_strm_data_g2f;
	assign strm_data_g2f_vld[0+:2] = glb_tile_gen_0_strm_data_g2f_vld;
	assign strm_ctrl_g2f[0+:2] = glb_tile_gen_0_strm_ctrl_g2f;
	assign data_flush[0] = glb_tile_gen_0_data_flush;
	assign cgra_cfg_g2f_cfg_wr_en[0+:2] = glb_tile_gen_0_cgra_cfg_g2f_cfg_wr_en;
	assign cgra_cfg_g2f_cfg_rd_en[0+:2] = glb_tile_gen_0_cgra_cfg_g2f_cfg_rd_en;
	assign cgra_cfg_g2f_cfg_addr[0+:64] = glb_tile_gen_0_cgra_cfg_g2f_cfg_addr;
	assign cgra_cfg_g2f_cfg_data[0+:64] = glb_tile_gen_0_cgra_cfg_g2f_cfg_data;
	assign cgra_cfg_pcfg_wr_en_esto[0] = glb_tile_gen_0_cgra_cfg_pcfg_wr_en_w2e_esto;
	assign cgra_cfg_pcfg_rd_en_esto[0] = glb_tile_gen_0_cgra_cfg_pcfg_rd_en_w2e_esto;
	assign cgra_cfg_pcfg_addr_esto[0+:32] = glb_tile_gen_0_cgra_cfg_pcfg_addr_w2e_esto;
	assign cgra_cfg_pcfg_data_esto[0+:32] = glb_tile_gen_0_cgra_cfg_pcfg_data_w2e_esto;
	assign cgra_cfg_pcfg_wr_en_wsto[0] = glb_tile_gen_0_cgra_cfg_pcfg_wr_en_e2w_wsto;
	assign cgra_cfg_pcfg_rd_en_wsto[0] = glb_tile_gen_0_cgra_cfg_pcfg_rd_en_e2w_wsto;
	assign cgra_cfg_pcfg_addr_wsto[0+:32] = glb_tile_gen_0_cgra_cfg_pcfg_addr_e2w_wsto;
	assign cgra_cfg_pcfg_data_wsto[0+:32] = glb_tile_gen_0_cgra_cfg_pcfg_data_e2w_wsto;
	assign cgra_cfg_jtag_wr_en_esto[0] = glb_tile_gen_0_cgra_cfg_jtag_wr_en_esto;
	assign cgra_cfg_jtag_rd_en_esto[0] = glb_tile_gen_0_cgra_cfg_jtag_rd_en_esto;
	assign cgra_cfg_jtag_addr_esto[0+:32] = glb_tile_gen_0_cgra_cfg_jtag_addr_esto;
	assign cgra_cfg_jtag_data_esto[0+:32] = glb_tile_gen_0_cgra_cfg_jtag_data_esto;
	assign cgra_cfg_jtag_rd_en_bypass_esto[0] = glb_tile_gen_0_cgra_cfg_jtag_rd_en_bypass_esto;
	assign cgra_cfg_jtag_addr_bypass_esto[0+:32] = glb_tile_gen_0_cgra_cfg_jtag_addr_bypass_esto;
	assign strm_f2g_interrupt_pulse_w[0] = glb_tile_gen_0_strm_f2g_interrupt_pulse;
	assign strm_g2f_interrupt_pulse_w[0] = glb_tile_gen_0_strm_g2f_interrupt_pulse;
	assign pcfg_g2f_interrupt_pulse_w[0] = glb_tile_gen_0_pcfg_g2f_interrupt_pulse;
	assign glb_tile_gen_1_clk_en_pcfg_broadcast = ~pcfg_broadcast_stall[1];
	assign glb_tile_gen_1_clk_en_master = glb_clk_en_master[1];
	assign glb_tile_gen_1_clk_en_bank_master = glb_clk_en_bank_master[1];
	assign strm_packet_w2e_esto[353] = glb_tile_gen_1_strm_wr_en_w2e_esto;
	assign strm_packet_w2e_esto[352-:8] = glb_tile_gen_1_strm_wr_strb_w2e_esto;
	assign strm_packet_w2e_esto[344-:19] = glb_tile_gen_1_strm_wr_addr_w2e_esto;
	assign strm_packet_w2e_esto[325-:64] = glb_tile_gen_1_strm_wr_data_w2e_esto;
	assign strm_packet_w2e_esto[261] = glb_tile_gen_1_strm_rd_en_w2e_esto;
	assign strm_packet_w2e_esto[260-:19] = glb_tile_gen_1_strm_rd_addr_w2e_esto;
	assign strm_packet_w2e_esto[241-:64] = glb_tile_gen_1_strm_rd_data_w2e_esto;
	assign strm_packet_w2e_esto[177] = glb_tile_gen_1_strm_rd_data_valid_w2e_esto;
	assign strm_packet_e2w_wsto[353] = glb_tile_gen_1_strm_wr_en_e2w_wsto;
	assign strm_packet_e2w_wsto[352-:8] = glb_tile_gen_1_strm_wr_strb_e2w_wsto;
	assign strm_packet_e2w_wsto[344-:19] = glb_tile_gen_1_strm_wr_addr_e2w_wsto;
	assign strm_packet_e2w_wsto[325-:64] = glb_tile_gen_1_strm_wr_data_e2w_wsto;
	assign strm_packet_e2w_wsto[261] = glb_tile_gen_1_strm_rd_en_e2w_wsto;
	assign strm_packet_e2w_wsto[260-:19] = glb_tile_gen_1_strm_rd_addr_e2w_wsto;
	assign strm_packet_e2w_wsto[241-:64] = glb_tile_gen_1_strm_rd_data_e2w_wsto;
	assign strm_packet_e2w_wsto[177] = glb_tile_gen_1_strm_rd_data_valid_e2w_wsto;
	assign pcfg_packet_w2e_esto[169] = glb_tile_gen_1_pcfg_rd_en_w2e_esto;
	assign pcfg_packet_w2e_esto[168-:19] = glb_tile_gen_1_pcfg_rd_addr_w2e_esto;
	assign pcfg_packet_w2e_esto[149-:64] = glb_tile_gen_1_pcfg_rd_data_w2e_esto;
	assign pcfg_packet_w2e_esto[85] = glb_tile_gen_1_pcfg_rd_data_valid_w2e_esto;
	assign pcfg_packet_e2w_wsto[169] = glb_tile_gen_1_pcfg_rd_en_e2w_wsto;
	assign pcfg_packet_e2w_wsto[168-:19] = glb_tile_gen_1_pcfg_rd_addr_e2w_wsto;
	assign pcfg_packet_e2w_wsto[149-:64] = glb_tile_gen_1_pcfg_rd_data_e2w_wsto;
	assign pcfg_packet_e2w_wsto[85] = glb_tile_gen_1_pcfg_rd_data_valid_e2w_wsto;
	assign cfg_tile_connected[2] = glb_tile_gen_1_cfg_tile_connected_esto;
	assign cfg_pcfg_tile_connected[2] = glb_tile_gen_1_cfg_pcfg_tile_connected_esto;
	assign strm_data_f2g_rdy[2+:2] = glb_tile_gen_1_strm_data_f2g_rdy;
	assign strm_data_g2f[32+:32] = glb_tile_gen_1_strm_data_g2f;
	assign strm_data_g2f_vld[2+:2] = glb_tile_gen_1_strm_data_g2f_vld;
	assign strm_ctrl_g2f[2+:2] = glb_tile_gen_1_strm_ctrl_g2f;
	assign data_flush[1] = glb_tile_gen_1_data_flush;
	assign cgra_cfg_g2f_cfg_wr_en[2+:2] = glb_tile_gen_1_cgra_cfg_g2f_cfg_wr_en;
	assign cgra_cfg_g2f_cfg_rd_en[2+:2] = glb_tile_gen_1_cgra_cfg_g2f_cfg_rd_en;
	assign cgra_cfg_g2f_cfg_addr[64+:64] = glb_tile_gen_1_cgra_cfg_g2f_cfg_addr;
	assign cgra_cfg_g2f_cfg_data[64+:64] = glb_tile_gen_1_cgra_cfg_g2f_cfg_data;
	assign cgra_cfg_pcfg_wr_en_esto[1] = glb_tile_gen_1_cgra_cfg_pcfg_wr_en_w2e_esto;
	assign cgra_cfg_pcfg_rd_en_esto[1] = glb_tile_gen_1_cgra_cfg_pcfg_rd_en_w2e_esto;
	assign cgra_cfg_pcfg_addr_esto[32+:32] = glb_tile_gen_1_cgra_cfg_pcfg_addr_w2e_esto;
	assign cgra_cfg_pcfg_data_esto[32+:32] = glb_tile_gen_1_cgra_cfg_pcfg_data_w2e_esto;
	assign cgra_cfg_pcfg_wr_en_wsto[1] = glb_tile_gen_1_cgra_cfg_pcfg_wr_en_e2w_wsto;
	assign cgra_cfg_pcfg_rd_en_wsto[1] = glb_tile_gen_1_cgra_cfg_pcfg_rd_en_e2w_wsto;
	assign cgra_cfg_pcfg_addr_wsto[32+:32] = glb_tile_gen_1_cgra_cfg_pcfg_addr_e2w_wsto;
	assign cgra_cfg_pcfg_data_wsto[32+:32] = glb_tile_gen_1_cgra_cfg_pcfg_data_e2w_wsto;
	assign cgra_cfg_jtag_wr_en_esto[1] = glb_tile_gen_1_cgra_cfg_jtag_wr_en_esto;
	assign cgra_cfg_jtag_rd_en_esto[1] = glb_tile_gen_1_cgra_cfg_jtag_rd_en_esto;
	assign cgra_cfg_jtag_addr_esto[32+:32] = glb_tile_gen_1_cgra_cfg_jtag_addr_esto;
	assign cgra_cfg_jtag_data_esto[32+:32] = glb_tile_gen_1_cgra_cfg_jtag_data_esto;
	assign cgra_cfg_jtag_rd_en_bypass_esto[1] = glb_tile_gen_1_cgra_cfg_jtag_rd_en_bypass_esto;
	assign cgra_cfg_jtag_addr_bypass_esto[32+:32] = glb_tile_gen_1_cgra_cfg_jtag_addr_bypass_esto;
	assign strm_f2g_interrupt_pulse_w[1] = glb_tile_gen_1_strm_f2g_interrupt_pulse;
	assign strm_g2f_interrupt_pulse_w[1] = glb_tile_gen_1_strm_g2f_interrupt_pulse;
	assign pcfg_g2f_interrupt_pulse_w[1] = glb_tile_gen_1_pcfg_g2f_interrupt_pulse;
	always @(posedge clk or posedge reset)
		if (reset) begin
			proc_wr_en_d <= 1'h0;
			proc_wr_strb_d <= 8'h00;
			proc_wr_addr_d <= 19'h00000;
			proc_wr_data_d <= 64'h0000000000000000;
			proc_rd_en_d <= 1'h0;
			proc_rd_addr_d <= 19'h00000;
		end
		else begin
			proc_wr_en_d <= proc_wr_en;
			proc_wr_strb_d <= proc_wr_strb;
			proc_wr_addr_d <= proc_wr_addr;
			proc_wr_data_d <= proc_wr_data;
			proc_rd_en_d <= proc_rd_en;
			proc_rd_addr_d <= proc_rd_addr;
		end
	always @(posedge clk or posedge reset)
		if (reset) begin
			sram_cfg_wr_en_d <= 1'h0;
			sram_cfg_wr_strb_d <= 8'h00;
			sram_cfg_wr_addr_d <= 19'h00000;
			sram_cfg_wr_data_d <= 64'h0000000000000000;
			sram_cfg_rd_en_d <= 1'h0;
			sram_cfg_rd_addr_d <= 19'h00000;
		end
		else begin
			sram_cfg_wr_en_d <= if_sram_cfg_wr_en;
			sram_cfg_wr_addr_d <= if_sram_cfg_wr_addr;
			if (if_sram_cfg_wr_addr[2] == 1'h0) begin
				sram_cfg_wr_data_d <= {32'h00000000, if_sram_cfg_wr_data};
				sram_cfg_wr_strb_d <= 8'h0f;
			end
			else begin
				sram_cfg_wr_data_d <= {if_sram_cfg_wr_data[31:0], 32'h00000000};
				sram_cfg_wr_strb_d <= 8'hf0;
			end
			sram_cfg_rd_en_d <= if_sram_cfg_rd_en;
			sram_cfg_rd_addr_d <= if_sram_cfg_rd_addr;
		end
	always @(posedge clk or posedge reset)
		if (reset) begin
			if_proc_tile2tile_0.wr_en <= 1'h0;
			if_proc_tile2tile_0.wr_strb <= 8'h00;
			if_proc_tile2tile_0.wr_addr <= 19'h00000;
			if_proc_tile2tile_0.wr_data <= 64'h0000000000000000;
		end
		else if (proc_wr_en_d) begin
			if_proc_tile2tile_0.wr_en <= proc_wr_en_d;
			if_proc_tile2tile_0.wr_strb <= proc_wr_strb_d;
			if_proc_tile2tile_0.wr_addr <= proc_wr_addr_d;
			if_proc_tile2tile_0.wr_data <= proc_wr_data_d;
		end
		else if (sram_cfg_wr_en_d) begin
			if_proc_tile2tile_0.wr_en <= sram_cfg_wr_en_d;
			if_proc_tile2tile_0.wr_strb <= sram_cfg_wr_strb_d;
			if_proc_tile2tile_0.wr_addr <= sram_cfg_wr_addr_d;
			if_proc_tile2tile_0.wr_data <= sram_cfg_wr_data_d;
		end
		else begin
			if_proc_tile2tile_0.wr_en <= proc_wr_en_d;
			if_proc_tile2tile_0.wr_strb <= proc_wr_strb_d;
			if_proc_tile2tile_0.wr_addr <= proc_wr_addr_d;
			if_proc_tile2tile_0.wr_data <= proc_wr_data_d;
		end
	always @(posedge clk or posedge reset)
		if (reset) begin
			if_proc_tile2tile_0.rd_en <= 1'h0;
			if_proc_tile2tile_0.rd_addr <= 19'h00000;
			proc_rd_type <= 1'h0;
			proc_rd_addr_sel <= 1'h0;
		end
		else if (proc_rd_en_d) begin
			if_proc_tile2tile_0.rd_en <= proc_rd_en_d;
			if_proc_tile2tile_0.rd_addr <= proc_rd_addr_d;
			proc_rd_type <= 1'h0;
			proc_rd_addr_sel <= 1'h0;
		end
		else if (sram_cfg_rd_en_d) begin
			if_proc_tile2tile_0.rd_en <= sram_cfg_rd_en_d;
			if_proc_tile2tile_0.rd_addr <= sram_cfg_rd_addr_d;
			proc_rd_addr_sel <= sram_cfg_rd_addr_d[2];
			proc_rd_type <= 1'h1;
		end
		else begin
			if_proc_tile2tile_0.rd_en <= proc_rd_en_d;
			if_proc_tile2tile_0.rd_addr <= proc_rd_addr_d;
			proc_rd_type <= proc_rd_type;
			proc_rd_addr_sel <= proc_rd_addr_sel;
		end
	always @(*)
		if (proc_rd_type == 1'h0) begin
			proc_rd_data_w = if_proc_tile2tile_0.rd_data;
			proc_rd_data_valid_w = if_proc_tile2tile_0.rd_data_valid;
			if_sram_cfg_rd_data_w = 32'h00000000;
			if_sram_cfg_rd_data_valid_w = 1'h0;
		end
		else if (proc_rd_type == 1'h1) begin
			proc_rd_data_w = 64'h0000000000000000;
			proc_rd_data_valid_w = 1'h0;
			if (proc_rd_addr_sel == 1'h0)
				if_sram_cfg_rd_data_w = if_proc_tile2tile_0.rd_data[31:0];
			else
				if_sram_cfg_rd_data_w = if_proc_tile2tile_0.rd_data[63:32];
			if_sram_cfg_rd_data_valid_w = if_proc_tile2tile_0.rd_data_valid;
		end
		else begin
			proc_rd_data_w = if_proc_tile2tile_0.rd_data;
			proc_rd_data_valid_w = if_proc_tile2tile_0.rd_data_valid;
			if_sram_cfg_rd_data_w = 32'h00000000;
			if_sram_cfg_rd_data_valid_w = 1'h0;
		end
	always @(posedge clk or posedge reset)
		if (reset) begin
			proc_rd_data <= 64'h0000000000000000;
			proc_rd_data_valid <= 1'h0;
			if_sram_cfg_rd_data <= 32'h00000000;
			if_sram_cfg_rd_data_valid <= 1'h0;
		end
		else begin
			proc_rd_data <= proc_rd_data_w;
			proc_rd_data_valid <= proc_rd_data_valid_w;
			if_sram_cfg_rd_data <= if_sram_cfg_rd_data_w;
			if_sram_cfg_rd_data_valid <= if_sram_cfg_rd_data_valid_w;
		end
	assign proc_wr_clk_en_gen_enable = proc_wr_en_d | sram_cfg_wr_en_d;
	assign if_proc_tile2tile_0.wr_clk_en = proc_wr_clk_en;
	assign proc_rd_clk_en_gen_enable = proc_rd_en_d | sram_cfg_rd_en_d;
	assign if_proc_tile2tile_0.rd_clk_en = proc_rd_clk_en;
	always @(posedge clk or posedge reset)
		if (reset) begin
			if_cfg_tile2tile_0.wr_en <= 1'h0;
			if_cfg_tile2tile_0.wr_clk_en <= 1'h0;
			if_cfg_tile2tile_0.wr_addr <= 12'h000;
			if_cfg_tile2tile_0.wr_data <= 32'h00000000;
			if_cfg_tile2tile_0.rd_en <= 1'h0;
			if_cfg_tile2tile_0.rd_clk_en <= 1'h0;
			if_cfg_tile2tile_0.rd_addr <= 12'h000;
		end
		else begin
			if_cfg_tile2tile_0.wr_en <= if_cfg_wr_en;
			if_cfg_tile2tile_0.wr_clk_en <= if_cfg_wr_clk_en;
			if_cfg_tile2tile_0.wr_addr <= if_cfg_wr_addr;
			if_cfg_tile2tile_0.wr_data <= if_cfg_wr_data;
			if_cfg_tile2tile_0.rd_en <= if_cfg_rd_en;
			if_cfg_tile2tile_0.rd_clk_en <= if_cfg_rd_clk_en;
			if_cfg_tile2tile_0.rd_addr <= if_cfg_rd_addr;
		end
	always @(posedge clk or posedge reset)
		if (reset) begin
			cgra_cfg_jtag_gc2glb_wr_en_d <= 1'h0;
			cgra_cfg_jtag_gc2glb_rd_en_d <= 1'h0;
			cgra_cfg_jtag_gc2glb_addr_d <= 32'h00000000;
			cgra_cfg_jtag_gc2glb_data_d <= 32'h00000000;
		end
		else begin
			cgra_cfg_jtag_gc2glb_wr_en_d <= cgra_cfg_jtag_gc2glb_wr_en;
			cgra_cfg_jtag_gc2glb_rd_en_d <= cgra_cfg_jtag_gc2glb_rd_en;
			cgra_cfg_jtag_gc2glb_addr_d <= cgra_cfg_jtag_gc2glb_addr;
			cgra_cfg_jtag_gc2glb_data_d <= cgra_cfg_jtag_gc2glb_data;
		end
	assign strm_packet_e2w_esti[177+:177] = 177'h000000000000000000000000000000000000000000000;
	assign pcfg_packet_e2w_esti[85+:85] = 85'h0000000000000000000000;
	assign strm_packet_e2w_esti[0+:177] = strm_packet_e2w_wsto[177+:177];
	assign pcfg_packet_e2w_esti[0+:85] = pcfg_packet_e2w_wsto[85+:85];
	assign strm_packet_w2e_wsti[0+:177] = 177'h000000000000000000000000000000000000000000000;
	assign pcfg_packet_w2e_wsti[0+:85] = 85'h0000000000000000000000;
	assign strm_packet_w2e_wsti[177+:177] = strm_packet_w2e_esto[0+:177];
	assign pcfg_packet_w2e_wsti[85+:85] = pcfg_packet_w2e_esto[0+:85];
	always @(*) begin
		cgra_cfg_jtag_rd_en_wsti[0] = 1'h0;
		cgra_cfg_jtag_wr_en_wsti[0] = cgra_cfg_jtag_gc2glb_wr_en_d;
		cgra_cfg_jtag_addr_wsti[0+:32] = cgra_cfg_jtag_gc2glb_addr_d;
		cgra_cfg_jtag_data_wsti[0+:32] = cgra_cfg_jtag_gc2glb_data_d;
		cgra_cfg_jtag_rd_en_bypass_wsti[0] = cgra_cfg_jtag_gc2glb_rd_en_d;
		cgra_cfg_jtag_addr_bypass_wsti[0+:32] = cgra_cfg_jtag_gc2glb_addr_d;
		cgra_cfg_pcfg_rd_en_wsti[0] = 1'h0;
		cgra_cfg_pcfg_wr_en_wsti[0] = 1'h0;
		cgra_cfg_pcfg_addr_wsti[0+:32] = 32'h00000000;
		cgra_cfg_pcfg_data_wsti[0+:32] = 32'h00000000;
		cgra_cfg_jtag_rd_en_wsti[1] = cgra_cfg_jtag_rd_en_esto[0];
		cgra_cfg_jtag_wr_en_wsti[1] = cgra_cfg_jtag_wr_en_esto[0];
		cgra_cfg_jtag_addr_wsti[32+:32] = cgra_cfg_jtag_addr_esto[0+:32];
		cgra_cfg_jtag_data_wsti[32+:32] = cgra_cfg_jtag_data_esto[0+:32];
		cgra_cfg_jtag_rd_en_bypass_wsti[1] = cgra_cfg_jtag_rd_en_bypass_esto[0];
		cgra_cfg_jtag_addr_bypass_wsti[32+:32] = cgra_cfg_jtag_addr_bypass_esto[0+:32];
		cgra_cfg_pcfg_rd_en_wsti[1] = cgra_cfg_pcfg_rd_en_esto[0];
		cgra_cfg_pcfg_wr_en_wsti[1] = cgra_cfg_pcfg_wr_en_esto[0];
		cgra_cfg_pcfg_addr_wsti[32+:32] = cgra_cfg_pcfg_addr_esto[0+:32];
		cgra_cfg_pcfg_data_wsti[32+:32] = cgra_cfg_pcfg_data_esto[0+:32];
	end
	always @(*) begin
		cgra_cfg_pcfg_rd_en_esti[0] = cgra_cfg_pcfg_rd_en_wsto[1];
		cgra_cfg_pcfg_wr_en_esti[0] = cgra_cfg_pcfg_wr_en_wsto[1];
		cgra_cfg_pcfg_addr_esti[0+:32] = cgra_cfg_pcfg_addr_wsto[32+:32];
		cgra_cfg_pcfg_data_esti[0+:32] = cgra_cfg_pcfg_data_wsto[32+:32];
		cgra_cfg_pcfg_rd_en_esti[1] = 1'h0;
		cgra_cfg_pcfg_wr_en_esti[1] = 1'h0;
		cgra_cfg_pcfg_addr_esti[32+:32] = 32'h00000000;
		cgra_cfg_pcfg_data_esti[32+:32] = 32'h00000000;
	end
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	always @(posedge clk or posedge reset)
		if (reset) begin : sv2v_autoblock_1
			reg [31:0] i;
			for (i = 0; i < 2; i = i + 1)
				begin
					strm_f2g_interrupt_pulse_d[sv2v_cast_1(i)] <= 1'h0;
					strm_g2f_interrupt_pulse_d[sv2v_cast_1(i)] <= 1'h0;
					pcfg_g2f_interrupt_pulse_d[sv2v_cast_1(i)] <= 1'h0;
				end
		end
		else begin : sv2v_autoblock_2
			reg [31:0] i;
			for (i = 0; i < 2; i = i + 1)
				begin
					strm_f2g_interrupt_pulse_d[sv2v_cast_1(i)] <= strm_f2g_interrupt_pulse_w[sv2v_cast_1(i)];
					strm_g2f_interrupt_pulse_d[sv2v_cast_1(i)] <= strm_g2f_interrupt_pulse_w[sv2v_cast_1(i)];
					pcfg_g2f_interrupt_pulse_d[sv2v_cast_1(i)] <= pcfg_g2f_interrupt_pulse_w[sv2v_cast_1(i)];
				end
		end
	assign if_cfg_rd_data = if_cfg_tile2tile_0.rd_data;
	assign if_cfg_rd_data_valid = if_cfg_tile2tile_0.rd_data_valid;
	assign flush_crossbar_in[0] = data_flush_d[0];
	assign flush_crossbar_in[1] = data_flush_d[1];
	assign flush_crossbar_sel_w = flush_crossbar_sel;
	glb_tile glb_tile_gen_0(
		.cfg_pcfg_tile_connected_wsti(cfg_pcfg_tile_connected[0]),
		.cfg_tile_connected_wsti(cfg_tile_connected[0]),
		.cgra_cfg_jtag_addr_bypass_wsti(cgra_cfg_jtag_addr_bypass_wsti[0+:32]),
		.cgra_cfg_jtag_addr_wsti(cgra_cfg_jtag_addr_wsti[0+:32]),
		.cgra_cfg_jtag_data_wsti(cgra_cfg_jtag_data_wsti[0+:32]),
		.cgra_cfg_jtag_rd_en_bypass_wsti(cgra_cfg_jtag_rd_en_bypass_wsti[0]),
		.cgra_cfg_jtag_rd_en_wsti(cgra_cfg_jtag_rd_en_wsti[0]),
		.cgra_cfg_jtag_wr_en_wsti(cgra_cfg_jtag_wr_en_wsti[0]),
		.cgra_cfg_pcfg_addr_e2w_esti(cgra_cfg_pcfg_addr_esti[0+:32]),
		.cgra_cfg_pcfg_addr_w2e_wsti(cgra_cfg_pcfg_addr_wsti[0+:32]),
		.cgra_cfg_pcfg_data_e2w_esti(cgra_cfg_pcfg_data_esti[0+:32]),
		.cgra_cfg_pcfg_data_w2e_wsti(cgra_cfg_pcfg_data_wsti[0+:32]),
		.cgra_cfg_pcfg_rd_en_e2w_esti(cgra_cfg_pcfg_rd_en_esti[0]),
		.cgra_cfg_pcfg_rd_en_w2e_wsti(cgra_cfg_pcfg_rd_en_wsti[0]),
		.cgra_cfg_pcfg_wr_en_e2w_esti(cgra_cfg_pcfg_wr_en_esti[0]),
		.cgra_cfg_pcfg_wr_en_w2e_wsti(cgra_cfg_pcfg_wr_en_wsti[0]),
		.clk(clk),
		.clk_en_bank_master(glb_tile_gen_0_clk_en_bank_master),
		.clk_en_master(glb_tile_gen_0_clk_en_master),
		.clk_en_pcfg_broadcast(glb_tile_gen_0_clk_en_pcfg_broadcast),
		.glb_tile_id(1'h0),
		.if_cfg_est_m_rd_data(if_cfg_tile2tile_1.rd_data),
		.if_cfg_est_m_rd_data_valid(if_cfg_tile2tile_1.rd_data_valid),
		.if_cfg_wst_s_rd_addr(if_cfg_tile2tile_0.rd_addr),
		.if_cfg_wst_s_rd_clk_en(if_cfg_tile2tile_0.rd_clk_en),
		.if_cfg_wst_s_rd_en(if_cfg_tile2tile_0.rd_en),
		.if_cfg_wst_s_wr_addr(if_cfg_tile2tile_0.wr_addr),
		.if_cfg_wst_s_wr_clk_en(if_cfg_tile2tile_0.wr_clk_en),
		.if_cfg_wst_s_wr_data(if_cfg_tile2tile_0.wr_data),
		.if_cfg_wst_s_wr_en(if_cfg_tile2tile_0.wr_en),
		.if_proc_est_m_rd_data(if_proc_tile2tile_1.rd_data),
		.if_proc_est_m_rd_data_valid(if_proc_tile2tile_1.rd_data_valid),
		.if_proc_wst_s_rd_addr(if_proc_tile2tile_0.rd_addr),
		.if_proc_wst_s_rd_clk_en(if_proc_tile2tile_0.rd_clk_en),
		.if_proc_wst_s_rd_en(if_proc_tile2tile_0.rd_en),
		.if_proc_wst_s_wr_addr(if_proc_tile2tile_0.wr_addr),
		.if_proc_wst_s_wr_clk_en(if_proc_tile2tile_0.wr_clk_en),
		.if_proc_wst_s_wr_data(if_proc_tile2tile_0.wr_data),
		.if_proc_wst_s_wr_en(if_proc_tile2tile_0.wr_en),
		.if_proc_wst_s_wr_strb(if_proc_tile2tile_0.wr_strb),
		.pcfg_rd_addr_e2w_esti(pcfg_packet_e2w_esti[83-:19]),
		.pcfg_rd_addr_w2e_wsti(pcfg_packet_w2e_wsti[83-:19]),
		.pcfg_rd_data_e2w_esti(pcfg_packet_e2w_esti[64-:64]),
		.pcfg_rd_data_valid_e2w_esti(pcfg_packet_e2w_esti[0]),
		.pcfg_rd_data_valid_w2e_wsti(pcfg_packet_w2e_wsti[0]),
		.pcfg_rd_data_w2e_wsti(pcfg_packet_w2e_wsti[64-:64]),
		.pcfg_rd_en_e2w_esti(pcfg_packet_e2w_esti[84]),
		.pcfg_rd_en_w2e_wsti(pcfg_packet_w2e_wsti[84]),
		.pcfg_start_pulse(pcfg_start_pulse[0]),
		.reset(reset),
		.strm_ctrl_f2g(strm_ctrl_f2g[0+:2]),
		.strm_data_f2g(strm_data_f2g[0+:32]),
		.strm_data_f2g_vld(strm_data_f2g_vld[0+:2]),
		.strm_data_g2f_rdy(strm_data_g2f_rdy[0+:2]),
		.strm_f2g_start_pulse(strm_f2g_start_pulse[0]),
		.strm_g2f_start_pulse(strm_g2f_start_pulse[0]),
		.strm_rd_addr_e2w_esti(strm_packet_e2w_esti[83-:19]),
		.strm_rd_addr_w2e_wsti(strm_packet_w2e_wsti[83-:19]),
		.strm_rd_data_e2w_esti(strm_packet_e2w_esti[64-:64]),
		.strm_rd_data_valid_e2w_esti(strm_packet_e2w_esti[0]),
		.strm_rd_data_valid_w2e_wsti(strm_packet_w2e_wsti[0]),
		.strm_rd_data_w2e_wsti(strm_packet_w2e_wsti[64-:64]),
		.strm_rd_en_e2w_esti(strm_packet_e2w_esti[84]),
		.strm_rd_en_w2e_wsti(strm_packet_w2e_wsti[84]),
		.strm_wr_addr_e2w_esti(strm_packet_e2w_esti[167-:19]),
		.strm_wr_addr_w2e_wsti(strm_packet_w2e_wsti[167-:19]),
		.strm_wr_data_e2w_esti(strm_packet_e2w_esti[148-:64]),
		.strm_wr_data_w2e_wsti(strm_packet_w2e_wsti[148-:64]),
		.strm_wr_en_e2w_esti(strm_packet_e2w_esti[176]),
		.strm_wr_en_w2e_wsti(strm_packet_w2e_wsti[176]),
		.strm_wr_strb_e2w_esti(strm_packet_e2w_esti[175-:8]),
		.strm_wr_strb_w2e_wsti(strm_packet_w2e_wsti[175-:8]),
		.cfg_pcfg_tile_connected_esto(glb_tile_gen_0_cfg_pcfg_tile_connected_esto),
		.cfg_tile_connected_esto(glb_tile_gen_0_cfg_tile_connected_esto),
		.cgra_cfg_g2f_cfg_addr(glb_tile_gen_0_cgra_cfg_g2f_cfg_addr),
		.cgra_cfg_g2f_cfg_data(glb_tile_gen_0_cgra_cfg_g2f_cfg_data),
		.cgra_cfg_g2f_cfg_rd_en(glb_tile_gen_0_cgra_cfg_g2f_cfg_rd_en),
		.cgra_cfg_g2f_cfg_wr_en(glb_tile_gen_0_cgra_cfg_g2f_cfg_wr_en),
		.cgra_cfg_jtag_addr_bypass_esto(glb_tile_gen_0_cgra_cfg_jtag_addr_bypass_esto),
		.cgra_cfg_jtag_addr_esto(glb_tile_gen_0_cgra_cfg_jtag_addr_esto),
		.cgra_cfg_jtag_data_esto(glb_tile_gen_0_cgra_cfg_jtag_data_esto),
		.cgra_cfg_jtag_rd_en_bypass_esto(glb_tile_gen_0_cgra_cfg_jtag_rd_en_bypass_esto),
		.cgra_cfg_jtag_rd_en_esto(glb_tile_gen_0_cgra_cfg_jtag_rd_en_esto),
		.cgra_cfg_jtag_wr_en_esto(glb_tile_gen_0_cgra_cfg_jtag_wr_en_esto),
		.cgra_cfg_pcfg_addr_e2w_wsto(glb_tile_gen_0_cgra_cfg_pcfg_addr_e2w_wsto),
		.cgra_cfg_pcfg_addr_w2e_esto(glb_tile_gen_0_cgra_cfg_pcfg_addr_w2e_esto),
		.cgra_cfg_pcfg_data_e2w_wsto(glb_tile_gen_0_cgra_cfg_pcfg_data_e2w_wsto),
		.cgra_cfg_pcfg_data_w2e_esto(glb_tile_gen_0_cgra_cfg_pcfg_data_w2e_esto),
		.cgra_cfg_pcfg_rd_en_e2w_wsto(glb_tile_gen_0_cgra_cfg_pcfg_rd_en_e2w_wsto),
		.cgra_cfg_pcfg_rd_en_w2e_esto(glb_tile_gen_0_cgra_cfg_pcfg_rd_en_w2e_esto),
		.cgra_cfg_pcfg_wr_en_e2w_wsto(glb_tile_gen_0_cgra_cfg_pcfg_wr_en_e2w_wsto),
		.cgra_cfg_pcfg_wr_en_w2e_esto(glb_tile_gen_0_cgra_cfg_pcfg_wr_en_w2e_esto),
		.data_flush(glb_tile_gen_0_data_flush),
		.if_cfg_est_m_rd_addr(if_cfg_tile2tile_1.rd_addr),
		.if_cfg_est_m_rd_clk_en(if_cfg_tile2tile_1.rd_clk_en),
		.if_cfg_est_m_rd_en(if_cfg_tile2tile_1.rd_en),
		.if_cfg_est_m_wr_addr(if_cfg_tile2tile_1.wr_addr),
		.if_cfg_est_m_wr_clk_en(if_cfg_tile2tile_1.wr_clk_en),
		.if_cfg_est_m_wr_data(if_cfg_tile2tile_1.wr_data),
		.if_cfg_est_m_wr_en(if_cfg_tile2tile_1.wr_en),
		.if_cfg_wst_s_rd_data(if_cfg_tile2tile_0.rd_data),
		.if_cfg_wst_s_rd_data_valid(if_cfg_tile2tile_0.rd_data_valid),
		.if_proc_est_m_rd_addr(if_proc_tile2tile_1.rd_addr),
		.if_proc_est_m_rd_clk_en(if_proc_tile2tile_1.rd_clk_en),
		.if_proc_est_m_rd_en(if_proc_tile2tile_1.rd_en),
		.if_proc_est_m_wr_addr(if_proc_tile2tile_1.wr_addr),
		.if_proc_est_m_wr_clk_en(if_proc_tile2tile_1.wr_clk_en),
		.if_proc_est_m_wr_data(if_proc_tile2tile_1.wr_data),
		.if_proc_est_m_wr_en(if_proc_tile2tile_1.wr_en),
		.if_proc_est_m_wr_strb(if_proc_tile2tile_1.wr_strb),
		.if_proc_wst_s_rd_data(if_proc_tile2tile_0.rd_data),
		.if_proc_wst_s_rd_data_valid(if_proc_tile2tile_0.rd_data_valid),
		.pcfg_g2f_interrupt_pulse(glb_tile_gen_0_pcfg_g2f_interrupt_pulse),
		.pcfg_rd_addr_e2w_wsto(glb_tile_gen_0_pcfg_rd_addr_e2w_wsto),
		.pcfg_rd_addr_w2e_esto(glb_tile_gen_0_pcfg_rd_addr_w2e_esto),
		.pcfg_rd_data_e2w_wsto(glb_tile_gen_0_pcfg_rd_data_e2w_wsto),
		.pcfg_rd_data_valid_e2w_wsto(glb_tile_gen_0_pcfg_rd_data_valid_e2w_wsto),
		.pcfg_rd_data_valid_w2e_esto(glb_tile_gen_0_pcfg_rd_data_valid_w2e_esto),
		.pcfg_rd_data_w2e_esto(glb_tile_gen_0_pcfg_rd_data_w2e_esto),
		.pcfg_rd_en_e2w_wsto(glb_tile_gen_0_pcfg_rd_en_e2w_wsto),
		.pcfg_rd_en_w2e_esto(glb_tile_gen_0_pcfg_rd_en_w2e_esto),
		.strm_ctrl_g2f(glb_tile_gen_0_strm_ctrl_g2f),
		.strm_data_f2g_rdy(glb_tile_gen_0_strm_data_f2g_rdy),
		.strm_data_g2f(glb_tile_gen_0_strm_data_g2f),
		.strm_data_g2f_vld(glb_tile_gen_0_strm_data_g2f_vld),
		.strm_f2g_interrupt_pulse(glb_tile_gen_0_strm_f2g_interrupt_pulse),
		.strm_g2f_interrupt_pulse(glb_tile_gen_0_strm_g2f_interrupt_pulse),
		.strm_rd_addr_e2w_wsto(glb_tile_gen_0_strm_rd_addr_e2w_wsto),
		.strm_rd_addr_w2e_esto(glb_tile_gen_0_strm_rd_addr_w2e_esto),
		.strm_rd_data_e2w_wsto(glb_tile_gen_0_strm_rd_data_e2w_wsto),
		.strm_rd_data_valid_e2w_wsto(glb_tile_gen_0_strm_rd_data_valid_e2w_wsto),
		.strm_rd_data_valid_w2e_esto(glb_tile_gen_0_strm_rd_data_valid_w2e_esto),
		.strm_rd_data_w2e_esto(glb_tile_gen_0_strm_rd_data_w2e_esto),
		.strm_rd_en_e2w_wsto(glb_tile_gen_0_strm_rd_en_e2w_wsto),
		.strm_rd_en_w2e_esto(glb_tile_gen_0_strm_rd_en_w2e_esto),
		.strm_wr_addr_e2w_wsto(glb_tile_gen_0_strm_wr_addr_e2w_wsto),
		.strm_wr_addr_w2e_esto(glb_tile_gen_0_strm_wr_addr_w2e_esto),
		.strm_wr_data_e2w_wsto(glb_tile_gen_0_strm_wr_data_e2w_wsto),
		.strm_wr_data_w2e_esto(glb_tile_gen_0_strm_wr_data_w2e_esto),
		.strm_wr_en_e2w_wsto(glb_tile_gen_0_strm_wr_en_e2w_wsto),
		.strm_wr_en_w2e_esto(glb_tile_gen_0_strm_wr_en_w2e_esto),
		.strm_wr_strb_e2w_wsto(glb_tile_gen_0_strm_wr_strb_e2w_wsto),
		.strm_wr_strb_w2e_esto(glb_tile_gen_0_strm_wr_strb_w2e_esto)
	);
	glb_tile glb_tile_gen_1(
		.cfg_pcfg_tile_connected_wsti(cfg_pcfg_tile_connected[1]),
		.cfg_tile_connected_wsti(cfg_tile_connected[1]),
		.cgra_cfg_jtag_addr_bypass_wsti(cgra_cfg_jtag_addr_bypass_wsti[32+:32]),
		.cgra_cfg_jtag_addr_wsti(cgra_cfg_jtag_addr_wsti[32+:32]),
		.cgra_cfg_jtag_data_wsti(cgra_cfg_jtag_data_wsti[32+:32]),
		.cgra_cfg_jtag_rd_en_bypass_wsti(cgra_cfg_jtag_rd_en_bypass_wsti[1]),
		.cgra_cfg_jtag_rd_en_wsti(cgra_cfg_jtag_rd_en_wsti[1]),
		.cgra_cfg_jtag_wr_en_wsti(cgra_cfg_jtag_wr_en_wsti[1]),
		.cgra_cfg_pcfg_addr_e2w_esti(cgra_cfg_pcfg_addr_esti[32+:32]),
		.cgra_cfg_pcfg_addr_w2e_wsti(cgra_cfg_pcfg_addr_wsti[32+:32]),
		.cgra_cfg_pcfg_data_e2w_esti(cgra_cfg_pcfg_data_esti[32+:32]),
		.cgra_cfg_pcfg_data_w2e_wsti(cgra_cfg_pcfg_data_wsti[32+:32]),
		.cgra_cfg_pcfg_rd_en_e2w_esti(cgra_cfg_pcfg_rd_en_esti[1]),
		.cgra_cfg_pcfg_rd_en_w2e_wsti(cgra_cfg_pcfg_rd_en_wsti[1]),
		.cgra_cfg_pcfg_wr_en_e2w_esti(cgra_cfg_pcfg_wr_en_esti[1]),
		.cgra_cfg_pcfg_wr_en_w2e_wsti(cgra_cfg_pcfg_wr_en_wsti[1]),
		.clk(clk),
		.clk_en_bank_master(glb_tile_gen_1_clk_en_bank_master),
		.clk_en_master(glb_tile_gen_1_clk_en_master),
		.clk_en_pcfg_broadcast(glb_tile_gen_1_clk_en_pcfg_broadcast),
		.glb_tile_id(1'h1),
		.if_cfg_est_m_rd_data(32'h00000000),
		.if_cfg_est_m_rd_data_valid(1'h0),
		.if_cfg_wst_s_rd_addr(if_cfg_tile2tile_1.rd_addr),
		.if_cfg_wst_s_rd_clk_en(if_cfg_tile2tile_1.rd_clk_en),
		.if_cfg_wst_s_rd_en(if_cfg_tile2tile_1.rd_en),
		.if_cfg_wst_s_wr_addr(if_cfg_tile2tile_1.wr_addr),
		.if_cfg_wst_s_wr_clk_en(if_cfg_tile2tile_1.wr_clk_en),
		.if_cfg_wst_s_wr_data(if_cfg_tile2tile_1.wr_data),
		.if_cfg_wst_s_wr_en(if_cfg_tile2tile_1.wr_en),
		.if_proc_est_m_rd_data(64'h0000000000000000),
		.if_proc_est_m_rd_data_valid(1'h0),
		.if_proc_wst_s_rd_addr(if_proc_tile2tile_1.rd_addr),
		.if_proc_wst_s_rd_clk_en(if_proc_tile2tile_1.rd_clk_en),
		.if_proc_wst_s_rd_en(if_proc_tile2tile_1.rd_en),
		.if_proc_wst_s_wr_addr(if_proc_tile2tile_1.wr_addr),
		.if_proc_wst_s_wr_clk_en(if_proc_tile2tile_1.wr_clk_en),
		.if_proc_wst_s_wr_data(if_proc_tile2tile_1.wr_data),
		.if_proc_wst_s_wr_en(if_proc_tile2tile_1.wr_en),
		.if_proc_wst_s_wr_strb(if_proc_tile2tile_1.wr_strb),
		.pcfg_rd_addr_e2w_esti(pcfg_packet_e2w_esti[168-:19]),
		.pcfg_rd_addr_w2e_wsti(pcfg_packet_w2e_wsti[168-:19]),
		.pcfg_rd_data_e2w_esti(pcfg_packet_e2w_esti[149-:64]),
		.pcfg_rd_data_valid_e2w_esti(pcfg_packet_e2w_esti[85]),
		.pcfg_rd_data_valid_w2e_wsti(pcfg_packet_w2e_wsti[85]),
		.pcfg_rd_data_w2e_wsti(pcfg_packet_w2e_wsti[149-:64]),
		.pcfg_rd_en_e2w_esti(pcfg_packet_e2w_esti[169]),
		.pcfg_rd_en_w2e_wsti(pcfg_packet_w2e_wsti[169]),
		.pcfg_start_pulse(pcfg_start_pulse[1]),
		.reset(reset),
		.strm_ctrl_f2g(strm_ctrl_f2g[2+:2]),
		.strm_data_f2g(strm_data_f2g[32+:32]),
		.strm_data_f2g_vld(strm_data_f2g_vld[2+:2]),
		.strm_data_g2f_rdy(strm_data_g2f_rdy[2+:2]),
		.strm_f2g_start_pulse(strm_f2g_start_pulse[1]),
		.strm_g2f_start_pulse(strm_g2f_start_pulse[1]),
		.strm_rd_addr_e2w_esti(strm_packet_e2w_esti[260-:19]),
		.strm_rd_addr_w2e_wsti(strm_packet_w2e_wsti[260-:19]),
		.strm_rd_data_e2w_esti(strm_packet_e2w_esti[241-:64]),
		.strm_rd_data_valid_e2w_esti(strm_packet_e2w_esti[177]),
		.strm_rd_data_valid_w2e_wsti(strm_packet_w2e_wsti[177]),
		.strm_rd_data_w2e_wsti(strm_packet_w2e_wsti[241-:64]),
		.strm_rd_en_e2w_esti(strm_packet_e2w_esti[261]),
		.strm_rd_en_w2e_wsti(strm_packet_w2e_wsti[261]),
		.strm_wr_addr_e2w_esti(strm_packet_e2w_esti[344-:19]),
		.strm_wr_addr_w2e_wsti(strm_packet_w2e_wsti[344-:19]),
		.strm_wr_data_e2w_esti(strm_packet_e2w_esti[325-:64]),
		.strm_wr_data_w2e_wsti(strm_packet_w2e_wsti[325-:64]),
		.strm_wr_en_e2w_esti(strm_packet_e2w_esti[353]),
		.strm_wr_en_w2e_wsti(strm_packet_w2e_wsti[353]),
		.strm_wr_strb_e2w_esti(strm_packet_e2w_esti[352-:8]),
		.strm_wr_strb_w2e_wsti(strm_packet_w2e_wsti[352-:8]),
		.cfg_pcfg_tile_connected_esto(glb_tile_gen_1_cfg_pcfg_tile_connected_esto),
		.cfg_tile_connected_esto(glb_tile_gen_1_cfg_tile_connected_esto),
		.cgra_cfg_g2f_cfg_addr(glb_tile_gen_1_cgra_cfg_g2f_cfg_addr),
		.cgra_cfg_g2f_cfg_data(glb_tile_gen_1_cgra_cfg_g2f_cfg_data),
		.cgra_cfg_g2f_cfg_rd_en(glb_tile_gen_1_cgra_cfg_g2f_cfg_rd_en),
		.cgra_cfg_g2f_cfg_wr_en(glb_tile_gen_1_cgra_cfg_g2f_cfg_wr_en),
		.cgra_cfg_jtag_addr_bypass_esto(glb_tile_gen_1_cgra_cfg_jtag_addr_bypass_esto),
		.cgra_cfg_jtag_addr_esto(glb_tile_gen_1_cgra_cfg_jtag_addr_esto),
		.cgra_cfg_jtag_data_esto(glb_tile_gen_1_cgra_cfg_jtag_data_esto),
		.cgra_cfg_jtag_rd_en_bypass_esto(glb_tile_gen_1_cgra_cfg_jtag_rd_en_bypass_esto),
		.cgra_cfg_jtag_rd_en_esto(glb_tile_gen_1_cgra_cfg_jtag_rd_en_esto),
		.cgra_cfg_jtag_wr_en_esto(glb_tile_gen_1_cgra_cfg_jtag_wr_en_esto),
		.cgra_cfg_pcfg_addr_e2w_wsto(glb_tile_gen_1_cgra_cfg_pcfg_addr_e2w_wsto),
		.cgra_cfg_pcfg_addr_w2e_esto(glb_tile_gen_1_cgra_cfg_pcfg_addr_w2e_esto),
		.cgra_cfg_pcfg_data_e2w_wsto(glb_tile_gen_1_cgra_cfg_pcfg_data_e2w_wsto),
		.cgra_cfg_pcfg_data_w2e_esto(glb_tile_gen_1_cgra_cfg_pcfg_data_w2e_esto),
		.cgra_cfg_pcfg_rd_en_e2w_wsto(glb_tile_gen_1_cgra_cfg_pcfg_rd_en_e2w_wsto),
		.cgra_cfg_pcfg_rd_en_w2e_esto(glb_tile_gen_1_cgra_cfg_pcfg_rd_en_w2e_esto),
		.cgra_cfg_pcfg_wr_en_e2w_wsto(glb_tile_gen_1_cgra_cfg_pcfg_wr_en_e2w_wsto),
		.cgra_cfg_pcfg_wr_en_w2e_esto(glb_tile_gen_1_cgra_cfg_pcfg_wr_en_w2e_esto),
		.data_flush(glb_tile_gen_1_data_flush),
		.if_cfg_est_m_rd_addr(if_cfg_tile2tile_2.rd_addr),
		.if_cfg_est_m_rd_clk_en(if_cfg_tile2tile_2.rd_clk_en),
		.if_cfg_est_m_rd_en(if_cfg_tile2tile_2.rd_en),
		.if_cfg_est_m_wr_addr(if_cfg_tile2tile_2.wr_addr),
		.if_cfg_est_m_wr_clk_en(if_cfg_tile2tile_2.wr_clk_en),
		.if_cfg_est_m_wr_data(if_cfg_tile2tile_2.wr_data),
		.if_cfg_est_m_wr_en(if_cfg_tile2tile_2.wr_en),
		.if_cfg_wst_s_rd_data(if_cfg_tile2tile_1.rd_data),
		.if_cfg_wst_s_rd_data_valid(if_cfg_tile2tile_1.rd_data_valid),
		.if_proc_est_m_rd_addr(if_proc_tile2tile_2.rd_addr),
		.if_proc_est_m_rd_clk_en(if_proc_tile2tile_2.rd_clk_en),
		.if_proc_est_m_rd_en(if_proc_tile2tile_2.rd_en),
		.if_proc_est_m_wr_addr(if_proc_tile2tile_2.wr_addr),
		.if_proc_est_m_wr_clk_en(if_proc_tile2tile_2.wr_clk_en),
		.if_proc_est_m_wr_data(if_proc_tile2tile_2.wr_data),
		.if_proc_est_m_wr_en(if_proc_tile2tile_2.wr_en),
		.if_proc_est_m_wr_strb(if_proc_tile2tile_2.wr_strb),
		.if_proc_wst_s_rd_data(if_proc_tile2tile_1.rd_data),
		.if_proc_wst_s_rd_data_valid(if_proc_tile2tile_1.rd_data_valid),
		.pcfg_g2f_interrupt_pulse(glb_tile_gen_1_pcfg_g2f_interrupt_pulse),
		.pcfg_rd_addr_e2w_wsto(glb_tile_gen_1_pcfg_rd_addr_e2w_wsto),
		.pcfg_rd_addr_w2e_esto(glb_tile_gen_1_pcfg_rd_addr_w2e_esto),
		.pcfg_rd_data_e2w_wsto(glb_tile_gen_1_pcfg_rd_data_e2w_wsto),
		.pcfg_rd_data_valid_e2w_wsto(glb_tile_gen_1_pcfg_rd_data_valid_e2w_wsto),
		.pcfg_rd_data_valid_w2e_esto(glb_tile_gen_1_pcfg_rd_data_valid_w2e_esto),
		.pcfg_rd_data_w2e_esto(glb_tile_gen_1_pcfg_rd_data_w2e_esto),
		.pcfg_rd_en_e2w_wsto(glb_tile_gen_1_pcfg_rd_en_e2w_wsto),
		.pcfg_rd_en_w2e_esto(glb_tile_gen_1_pcfg_rd_en_w2e_esto),
		.strm_ctrl_g2f(glb_tile_gen_1_strm_ctrl_g2f),
		.strm_data_f2g_rdy(glb_tile_gen_1_strm_data_f2g_rdy),
		.strm_data_g2f(glb_tile_gen_1_strm_data_g2f),
		.strm_data_g2f_vld(glb_tile_gen_1_strm_data_g2f_vld),
		.strm_f2g_interrupt_pulse(glb_tile_gen_1_strm_f2g_interrupt_pulse),
		.strm_g2f_interrupt_pulse(glb_tile_gen_1_strm_g2f_interrupt_pulse),
		.strm_rd_addr_e2w_wsto(glb_tile_gen_1_strm_rd_addr_e2w_wsto),
		.strm_rd_addr_w2e_esto(glb_tile_gen_1_strm_rd_addr_w2e_esto),
		.strm_rd_data_e2w_wsto(glb_tile_gen_1_strm_rd_data_e2w_wsto),
		.strm_rd_data_valid_e2w_wsto(glb_tile_gen_1_strm_rd_data_valid_e2w_wsto),
		.strm_rd_data_valid_w2e_esto(glb_tile_gen_1_strm_rd_data_valid_w2e_esto),
		.strm_rd_data_w2e_esto(glb_tile_gen_1_strm_rd_data_w2e_esto),
		.strm_rd_en_e2w_wsto(glb_tile_gen_1_strm_rd_en_e2w_wsto),
		.strm_rd_en_w2e_esto(glb_tile_gen_1_strm_rd_en_w2e_esto),
		.strm_wr_addr_e2w_wsto(glb_tile_gen_1_strm_wr_addr_e2w_wsto),
		.strm_wr_addr_w2e_esto(glb_tile_gen_1_strm_wr_addr_w2e_esto),
		.strm_wr_data_e2w_wsto(glb_tile_gen_1_strm_wr_data_e2w_wsto),
		.strm_wr_data_w2e_esto(glb_tile_gen_1_strm_wr_data_w2e_esto),
		.strm_wr_en_e2w_wsto(glb_tile_gen_1_strm_wr_en_e2w_wsto),
		.strm_wr_en_w2e_esto(glb_tile_gen_1_strm_wr_en_w2e_esto),
		.strm_wr_strb_e2w_wsto(glb_tile_gen_1_strm_wr_strb_e2w_wsto),
		.strm_wr_strb_w2e_esto(glb_tile_gen_1_strm_wr_strb_w2e_esto)
	);
	glb_clk_en_gen_5 #(.cnt(32'h00000005)) proc_wr_clk_en_gen(
		.clk(clk),
		.enable(proc_wr_clk_en_gen_enable),
		.reset(reset),
		.clk_en(proc_wr_clk_en)
	);
	glb_clk_en_gen_11 #(.cnt(32'h0000000b)) proc_rd_clk_en_gen(
		.clk(clk),
		.enable(proc_rd_clk_en_gen_enable),
		.reset(reset),
		.clk_en(proc_rd_clk_en)
	);
	pipeline_w_2_d_1 flush_pipeline(
		.clk(clk),
		.clk_en(1'h1),
		.in_(data_flush),
		.reset(reset),
		.out_(data_flush_d)
	);
	glb_crossbar_I_2_O_1_W_1 flush_crossbar(
		.in_(flush_crossbar_in),
		.sel_(flush_crossbar_sel_w),
		.out_(strm_data_flush_g2f)
	);
endmodule
module global_buffer_W (
	cgra_cfg_jtag_gc2glb_addr,
	cgra_cfg_jtag_gc2glb_data,
	cgra_cfg_jtag_gc2glb_rd_en,
	cgra_cfg_jtag_gc2glb_wr_en,
	cgra_stall_in,
	clk,
	flush_crossbar_sel,
	glb_clk_en_bank_master,
	glb_clk_en_master,
	if_cfg_rd_addr,
	if_cfg_rd_clk_en,
	if_cfg_rd_en,
	if_cfg_wr_addr,
	if_cfg_wr_clk_en,
	if_cfg_wr_data,
	if_cfg_wr_en,
	if_sram_cfg_rd_addr,
	if_sram_cfg_rd_en,
	if_sram_cfg_wr_addr,
	if_sram_cfg_wr_data,
	if_sram_cfg_wr_en,
	pcfg_broadcast_stall,
	pcfg_start_pulse,
	proc_rd_addr,
	proc_rd_en,
	proc_wr_addr,
	proc_wr_data,
	proc_wr_en,
	proc_wr_strb,
	reset,
	strm_ctrl_f2g_0_0,
	strm_ctrl_f2g_0_1,
	strm_ctrl_f2g_1_0,
	strm_ctrl_f2g_1_1,
	strm_data_f2g_0_0,
	strm_data_f2g_0_1,
	strm_data_f2g_1_0,
	strm_data_f2g_1_1,
	strm_data_f2g_vld_0_0,
	strm_data_f2g_vld_0_1,
	strm_data_f2g_vld_1_0,
	strm_data_f2g_vld_1_1,
	strm_data_g2f_rdy_0_0,
	strm_data_g2f_rdy_0_1,
	strm_data_g2f_rdy_1_0,
	strm_data_g2f_rdy_1_1,
	strm_f2g_start_pulse,
	strm_g2f_start_pulse,
	cgra_cfg_g2f_cfg_addr_0_0,
	cgra_cfg_g2f_cfg_addr_0_1,
	cgra_cfg_g2f_cfg_addr_1_0,
	cgra_cfg_g2f_cfg_addr_1_1,
	cgra_cfg_g2f_cfg_data_0_0,
	cgra_cfg_g2f_cfg_data_0_1,
	cgra_cfg_g2f_cfg_data_1_0,
	cgra_cfg_g2f_cfg_data_1_1,
	cgra_cfg_g2f_cfg_rd_en_0_0,
	cgra_cfg_g2f_cfg_rd_en_0_1,
	cgra_cfg_g2f_cfg_rd_en_1_0,
	cgra_cfg_g2f_cfg_rd_en_1_1,
	cgra_cfg_g2f_cfg_wr_en_0_0,
	cgra_cfg_g2f_cfg_wr_en_0_1,
	cgra_cfg_g2f_cfg_wr_en_1_0,
	cgra_cfg_g2f_cfg_wr_en_1_1,
	cgra_stall,
	if_cfg_rd_data,
	if_cfg_rd_data_valid,
	if_sram_cfg_rd_data,
	if_sram_cfg_rd_data_valid,
	pcfg_g2f_interrupt_pulse,
	proc_rd_data,
	proc_rd_data_valid,
	strm_ctrl_g2f_0_0,
	strm_ctrl_g2f_0_1,
	strm_ctrl_g2f_1_0,
	strm_ctrl_g2f_1_1,
	strm_data_f2g_rdy_0_0,
	strm_data_f2g_rdy_0_1,
	strm_data_f2g_rdy_1_0,
	strm_data_f2g_rdy_1_1,
	strm_data_flush_g2f,
	strm_data_g2f_0_0,
	strm_data_g2f_0_1,
	strm_data_g2f_1_0,
	strm_data_g2f_1_1,
	strm_data_g2f_vld_0_0,
	strm_data_g2f_vld_0_1,
	strm_data_g2f_vld_1_0,
	strm_data_g2f_vld_1_1,
	strm_f2g_interrupt_pulse,
	strm_g2f_interrupt_pulse
);
	input wire [31:0] cgra_cfg_jtag_gc2glb_addr;
	input wire [31:0] cgra_cfg_jtag_gc2glb_data;
	input wire cgra_cfg_jtag_gc2glb_rd_en;
	input wire cgra_cfg_jtag_gc2glb_wr_en;
	input wire [3:0] cgra_stall_in;
	input wire clk;
	input wire flush_crossbar_sel;
	input wire [1:0] glb_clk_en_bank_master;
	input wire [1:0] glb_clk_en_master;
	input wire [11:0] if_cfg_rd_addr;
	input wire if_cfg_rd_clk_en;
	input wire if_cfg_rd_en;
	input wire [11:0] if_cfg_wr_addr;
	input wire if_cfg_wr_clk_en;
	input wire [31:0] if_cfg_wr_data;
	input wire if_cfg_wr_en;
	input wire [18:0] if_sram_cfg_rd_addr;
	input wire if_sram_cfg_rd_en;
	input wire [18:0] if_sram_cfg_wr_addr;
	input wire [31:0] if_sram_cfg_wr_data;
	input wire if_sram_cfg_wr_en;
	input wire [1:0] pcfg_broadcast_stall;
	input wire [1:0] pcfg_start_pulse;
	input wire [18:0] proc_rd_addr;
	input wire proc_rd_en;
	input wire [18:0] proc_wr_addr;
	input wire [63:0] proc_wr_data;
	input wire proc_wr_en;
	input wire [7:0] proc_wr_strb;
	input wire reset;
	input wire strm_ctrl_f2g_0_0;
	input wire strm_ctrl_f2g_0_1;
	input wire strm_ctrl_f2g_1_0;
	input wire strm_ctrl_f2g_1_1;
	input wire [15:0] strm_data_f2g_0_0;
	input wire [15:0] strm_data_f2g_0_1;
	input wire [15:0] strm_data_f2g_1_0;
	input wire [15:0] strm_data_f2g_1_1;
	input wire strm_data_f2g_vld_0_0;
	input wire strm_data_f2g_vld_0_1;
	input wire strm_data_f2g_vld_1_0;
	input wire strm_data_f2g_vld_1_1;
	input wire strm_data_g2f_rdy_0_0;
	input wire strm_data_g2f_rdy_0_1;
	input wire strm_data_g2f_rdy_1_0;
	input wire strm_data_g2f_rdy_1_1;
	input wire [1:0] strm_f2g_start_pulse;
	input wire [1:0] strm_g2f_start_pulse;
	output wire [31:0] cgra_cfg_g2f_cfg_addr_0_0;
	output wire [31:0] cgra_cfg_g2f_cfg_addr_0_1;
	output wire [31:0] cgra_cfg_g2f_cfg_addr_1_0;
	output wire [31:0] cgra_cfg_g2f_cfg_addr_1_1;
	output wire [31:0] cgra_cfg_g2f_cfg_data_0_0;
	output wire [31:0] cgra_cfg_g2f_cfg_data_0_1;
	output wire [31:0] cgra_cfg_g2f_cfg_data_1_0;
	output wire [31:0] cgra_cfg_g2f_cfg_data_1_1;
	output wire cgra_cfg_g2f_cfg_rd_en_0_0;
	output wire cgra_cfg_g2f_cfg_rd_en_0_1;
	output wire cgra_cfg_g2f_cfg_rd_en_1_0;
	output wire cgra_cfg_g2f_cfg_rd_en_1_1;
	output wire cgra_cfg_g2f_cfg_wr_en_0_0;
	output wire cgra_cfg_g2f_cfg_wr_en_0_1;
	output wire cgra_cfg_g2f_cfg_wr_en_1_0;
	output wire cgra_cfg_g2f_cfg_wr_en_1_1;
	output wire [3:0] cgra_stall;
	output wire [31:0] if_cfg_rd_data;
	output wire if_cfg_rd_data_valid;
	output wire [31:0] if_sram_cfg_rd_data;
	output wire if_sram_cfg_rd_data_valid;
	output wire [1:0] pcfg_g2f_interrupt_pulse;
	output wire [63:0] proc_rd_data;
	output wire proc_rd_data_valid;
	output wire strm_ctrl_g2f_0_0;
	output wire strm_ctrl_g2f_0_1;
	output wire strm_ctrl_g2f_1_0;
	output wire strm_ctrl_g2f_1_1;
	output wire strm_data_f2g_rdy_0_0;
	output wire strm_data_f2g_rdy_0_1;
	output wire strm_data_f2g_rdy_1_0;
	output wire strm_data_f2g_rdy_1_1;
	output wire strm_data_flush_g2f;
	output wire [15:0] strm_data_g2f_0_0;
	output wire [15:0] strm_data_g2f_0_1;
	output wire [15:0] strm_data_g2f_1_0;
	output wire [15:0] strm_data_g2f_1_1;
	output wire strm_data_g2f_vld_0_0;
	output wire strm_data_g2f_vld_0_1;
	output wire strm_data_g2f_vld_1_0;
	output wire strm_data_g2f_vld_1_1;
	output wire [1:0] strm_f2g_interrupt_pulse;
	output wire [1:0] strm_g2f_interrupt_pulse;
	wire [127:0] global_buffer_cgra_cfg_g2f_cfg_addr;
	wire [127:0] global_buffer_cgra_cfg_g2f_cfg_data;
	wire [3:0] global_buffer_cgra_cfg_g2f_cfg_rd_en;
	wire [3:0] global_buffer_cgra_cfg_g2f_cfg_wr_en;
	wire [3:0] global_buffer_strm_ctrl_f2g;
	wire [3:0] global_buffer_strm_ctrl_g2f;
	wire [63:0] global_buffer_strm_data_f2g;
	wire [3:0] global_buffer_strm_data_f2g_rdy;
	wire [3:0] global_buffer_strm_data_f2g_vld;
	wire [63:0] global_buffer_strm_data_g2f;
	wire [3:0] global_buffer_strm_data_g2f_rdy;
	wire [3:0] global_buffer_strm_data_g2f_vld;
	assign cgra_cfg_g2f_cfg_addr_0_0 = global_buffer_cgra_cfg_g2f_cfg_addr[0+:32];
	assign cgra_cfg_g2f_cfg_addr_0_1 = global_buffer_cgra_cfg_g2f_cfg_addr[32+:32];
	assign cgra_cfg_g2f_cfg_addr_1_0 = global_buffer_cgra_cfg_g2f_cfg_addr[64+:32];
	assign cgra_cfg_g2f_cfg_addr_1_1 = global_buffer_cgra_cfg_g2f_cfg_addr[96+:32];
	assign cgra_cfg_g2f_cfg_data_0_0 = global_buffer_cgra_cfg_g2f_cfg_data[0+:32];
	assign cgra_cfg_g2f_cfg_data_0_1 = global_buffer_cgra_cfg_g2f_cfg_data[32+:32];
	assign cgra_cfg_g2f_cfg_data_1_0 = global_buffer_cgra_cfg_g2f_cfg_data[64+:32];
	assign cgra_cfg_g2f_cfg_data_1_1 = global_buffer_cgra_cfg_g2f_cfg_data[96+:32];
	assign cgra_cfg_g2f_cfg_rd_en_0_0 = global_buffer_cgra_cfg_g2f_cfg_rd_en[0];
	assign cgra_cfg_g2f_cfg_rd_en_0_1 = global_buffer_cgra_cfg_g2f_cfg_rd_en[1];
	assign cgra_cfg_g2f_cfg_rd_en_1_0 = global_buffer_cgra_cfg_g2f_cfg_rd_en[2];
	assign cgra_cfg_g2f_cfg_rd_en_1_1 = global_buffer_cgra_cfg_g2f_cfg_rd_en[3];
	assign cgra_cfg_g2f_cfg_wr_en_0_0 = global_buffer_cgra_cfg_g2f_cfg_wr_en[0];
	assign cgra_cfg_g2f_cfg_wr_en_0_1 = global_buffer_cgra_cfg_g2f_cfg_wr_en[1];
	assign cgra_cfg_g2f_cfg_wr_en_1_0 = global_buffer_cgra_cfg_g2f_cfg_wr_en[2];
	assign cgra_cfg_g2f_cfg_wr_en_1_1 = global_buffer_cgra_cfg_g2f_cfg_wr_en[3];
	assign global_buffer_strm_ctrl_f2g[0] = strm_ctrl_f2g_0_0;
	assign global_buffer_strm_ctrl_f2g[1] = strm_ctrl_f2g_0_1;
	assign global_buffer_strm_ctrl_f2g[2] = strm_ctrl_f2g_1_0;
	assign global_buffer_strm_ctrl_f2g[3] = strm_ctrl_f2g_1_1;
	assign strm_ctrl_g2f_0_0 = global_buffer_strm_ctrl_g2f[0];
	assign strm_ctrl_g2f_0_1 = global_buffer_strm_ctrl_g2f[1];
	assign strm_ctrl_g2f_1_0 = global_buffer_strm_ctrl_g2f[2];
	assign strm_ctrl_g2f_1_1 = global_buffer_strm_ctrl_g2f[3];
	assign global_buffer_strm_data_f2g[0+:16] = strm_data_f2g_0_0;
	assign global_buffer_strm_data_f2g[16+:16] = strm_data_f2g_0_1;
	assign global_buffer_strm_data_f2g[32+:16] = strm_data_f2g_1_0;
	assign global_buffer_strm_data_f2g[48+:16] = strm_data_f2g_1_1;
	assign strm_data_f2g_rdy_0_0 = global_buffer_strm_data_f2g_rdy[0];
	assign strm_data_f2g_rdy_0_1 = global_buffer_strm_data_f2g_rdy[1];
	assign strm_data_f2g_rdy_1_0 = global_buffer_strm_data_f2g_rdy[2];
	assign strm_data_f2g_rdy_1_1 = global_buffer_strm_data_f2g_rdy[3];
	assign global_buffer_strm_data_f2g_vld[0] = strm_data_f2g_vld_0_0;
	assign global_buffer_strm_data_f2g_vld[1] = strm_data_f2g_vld_0_1;
	assign global_buffer_strm_data_f2g_vld[2] = strm_data_f2g_vld_1_0;
	assign global_buffer_strm_data_f2g_vld[3] = strm_data_f2g_vld_1_1;
	assign strm_data_g2f_0_0 = global_buffer_strm_data_g2f[0+:16];
	assign strm_data_g2f_0_1 = global_buffer_strm_data_g2f[16+:16];
	assign strm_data_g2f_1_0 = global_buffer_strm_data_g2f[32+:16];
	assign strm_data_g2f_1_1 = global_buffer_strm_data_g2f[48+:16];
	assign global_buffer_strm_data_g2f_rdy[0] = strm_data_g2f_rdy_0_0;
	assign global_buffer_strm_data_g2f_rdy[1] = strm_data_g2f_rdy_0_1;
	assign global_buffer_strm_data_g2f_rdy[2] = strm_data_g2f_rdy_1_0;
	assign global_buffer_strm_data_g2f_rdy[3] = strm_data_g2f_rdy_1_1;
	assign strm_data_g2f_vld_0_0 = global_buffer_strm_data_g2f_vld[0];
	assign strm_data_g2f_vld_0_1 = global_buffer_strm_data_g2f_vld[1];
	assign strm_data_g2f_vld_1_0 = global_buffer_strm_data_g2f_vld[2];
	assign strm_data_g2f_vld_1_1 = global_buffer_strm_data_g2f_vld[3];
	global_buffer global_buffer(
		.cgra_cfg_jtag_gc2glb_addr(cgra_cfg_jtag_gc2glb_addr),
		.cgra_cfg_jtag_gc2glb_data(cgra_cfg_jtag_gc2glb_data),
		.cgra_cfg_jtag_gc2glb_rd_en(cgra_cfg_jtag_gc2glb_rd_en),
		.cgra_cfg_jtag_gc2glb_wr_en(cgra_cfg_jtag_gc2glb_wr_en),
		.cgra_stall_in(cgra_stall_in),
		.clk(clk),
		.flush_crossbar_sel(flush_crossbar_sel),
		.glb_clk_en_bank_master(glb_clk_en_bank_master),
		.glb_clk_en_master(glb_clk_en_master),
		.if_cfg_rd_addr(if_cfg_rd_addr),
		.if_cfg_rd_clk_en(if_cfg_rd_clk_en),
		.if_cfg_rd_en(if_cfg_rd_en),
		.if_cfg_wr_addr(if_cfg_wr_addr),
		.if_cfg_wr_clk_en(if_cfg_wr_clk_en),
		.if_cfg_wr_data(if_cfg_wr_data),
		.if_cfg_wr_en(if_cfg_wr_en),
		.if_sram_cfg_rd_addr(if_sram_cfg_rd_addr),
		.if_sram_cfg_rd_en(if_sram_cfg_rd_en),
		.if_sram_cfg_wr_addr(if_sram_cfg_wr_addr),
		.if_sram_cfg_wr_data(if_sram_cfg_wr_data),
		.if_sram_cfg_wr_en(if_sram_cfg_wr_en),
		.pcfg_broadcast_stall(pcfg_broadcast_stall),
		.pcfg_start_pulse(pcfg_start_pulse),
		.proc_rd_addr(proc_rd_addr),
		.proc_rd_en(proc_rd_en),
		.proc_wr_addr(proc_wr_addr),
		.proc_wr_data(proc_wr_data),
		.proc_wr_en(proc_wr_en),
		.proc_wr_strb(proc_wr_strb),
		.reset(reset),
		.strm_ctrl_f2g(global_buffer_strm_ctrl_f2g),
		.strm_data_f2g(global_buffer_strm_data_f2g),
		.strm_data_f2g_vld(global_buffer_strm_data_f2g_vld),
		.strm_data_g2f_rdy(global_buffer_strm_data_g2f_rdy),
		.strm_f2g_start_pulse(strm_f2g_start_pulse),
		.strm_g2f_start_pulse(strm_g2f_start_pulse),
		.cgra_cfg_g2f_cfg_addr(global_buffer_cgra_cfg_g2f_cfg_addr),
		.cgra_cfg_g2f_cfg_data(global_buffer_cgra_cfg_g2f_cfg_data),
		.cgra_cfg_g2f_cfg_rd_en(global_buffer_cgra_cfg_g2f_cfg_rd_en),
		.cgra_cfg_g2f_cfg_wr_en(global_buffer_cgra_cfg_g2f_cfg_wr_en),
		.cgra_stall(cgra_stall),
		.if_cfg_rd_data(if_cfg_rd_data),
		.if_cfg_rd_data_valid(if_cfg_rd_data_valid),
		.if_sram_cfg_rd_data(if_sram_cfg_rd_data),
		.if_sram_cfg_rd_data_valid(if_sram_cfg_rd_data_valid),
		.pcfg_g2f_interrupt_pulse(pcfg_g2f_interrupt_pulse),
		.proc_rd_data(proc_rd_data),
		.proc_rd_data_valid(proc_rd_data_valid),
		.strm_ctrl_g2f(global_buffer_strm_ctrl_g2f),
		.strm_data_f2g_rdy(global_buffer_strm_data_f2g_rdy),
		.strm_data_flush_g2f(strm_data_flush_g2f),
		.strm_data_g2f(global_buffer_strm_data_g2f),
		.strm_data_g2f_vld(global_buffer_strm_data_g2f_vld),
		.strm_f2g_interrupt_pulse(strm_f2g_interrupt_pulse),
		.strm_g2f_interrupt_pulse(strm_g2f_interrupt_pulse)
	);
endmodule
module pipeline_w_144_d_0 (
	clk,
	clk_en,
	in_,
	reset,
	out_
);
	input wire clk;
	input wire clk_en;
	input wire [143:0] in_;
	input wire reset;
	output wire [143:0] out_;
	assign out_ = in_;
endmodule
module pipeline_w_18_d_0 (
	clk,
	clk_en,
	in_,
	reset,
	out_
);
	input wire clk;
	input wire clk_en;
	input wire [17:0] in_;
	input wire reset;
	output wire [17:0] out_;
	assign out_ = in_;
endmodule
module pipeline_w_1_d_0 (
	clk,
	clk_en,
	in_,
	reset,
	out_
);
	input wire clk;
	input wire clk_en;
	input wire in_;
	input wire reset;
	output wire out_;
	assign out_ = in_;
endmodule
module pipeline_w_1_d_1 (
	clk,
	clk_en,
	in_,
	reset,
	out_
);
	input wire clk;
	input wire clk_en;
	input wire in_;
	input wire reset;
	output wire out_;
	reg pipeline_r;
	assign out_ = pipeline_r;
	always @(posedge clk or posedge reset)
		if (reset)
			pipeline_r <= 1'h0;
		else if (clk_en)
			pipeline_r <= in_;
endmodule
module pipeline_w_1_d_12_array (
	clk,
	clk_en,
	in_,
	reset,
	out_
);
	input wire clk;
	input wire clk_en;
	input wire in_;
	input wire reset;
	output wire [11:0] out_;
	reg [11:0] pipeline_r;
	assign out_ = pipeline_r;
	always @(posedge clk or posedge reset)
		if (reset) begin
			pipeline_r[0] <= 1'h0;
			pipeline_r[1] <= 1'h0;
			pipeline_r[2] <= 1'h0;
			pipeline_r[3] <= 1'h0;
			pipeline_r[4] <= 1'h0;
			pipeline_r[5] <= 1'h0;
			pipeline_r[6] <= 1'h0;
			pipeline_r[7] <= 1'h0;
			pipeline_r[8] <= 1'h0;
			pipeline_r[9] <= 1'h0;
			pipeline_r[10] <= 1'h0;
			pipeline_r[11] <= 1'h0;
		end
		else if (clk_en) begin
			pipeline_r[0] <= in_;
			pipeline_r[1] <= pipeline_r[4'h0];
			pipeline_r[2] <= pipeline_r[4'h1];
			pipeline_r[3] <= pipeline_r[4'h2];
			pipeline_r[4] <= pipeline_r[4'h3];
			pipeline_r[5] <= pipeline_r[4'h4];
			pipeline_r[6] <= pipeline_r[4'h5];
			pipeline_r[7] <= pipeline_r[4'h6];
			pipeline_r[8] <= pipeline_r[4'h7];
			pipeline_r[9] <= pipeline_r[4'h8];
			pipeline_r[10] <= pipeline_r[4'h9];
			pipeline_r[11] <= pipeline_r[4'ha];
		end
endmodule
module pipeline_w_1_d_20_array (
	clk,
	clk_en,
	in_,
	reset,
	out_
);
	input wire clk;
	input wire clk_en;
	input wire in_;
	input wire reset;
	output wire [19:0] out_;
	reg [19:0] pipeline_r;
	assign out_ = pipeline_r;
	always @(posedge clk or posedge reset)
		if (reset) begin
			pipeline_r[0] <= 1'h0;
			pipeline_r[1] <= 1'h0;
			pipeline_r[2] <= 1'h0;
			pipeline_r[3] <= 1'h0;
			pipeline_r[4] <= 1'h0;
			pipeline_r[5] <= 1'h0;
			pipeline_r[6] <= 1'h0;
			pipeline_r[7] <= 1'h0;
			pipeline_r[8] <= 1'h0;
			pipeline_r[9] <= 1'h0;
			pipeline_r[10] <= 1'h0;
			pipeline_r[11] <= 1'h0;
			pipeline_r[12] <= 1'h0;
			pipeline_r[13] <= 1'h0;
			pipeline_r[14] <= 1'h0;
			pipeline_r[15] <= 1'h0;
			pipeline_r[16] <= 1'h0;
			pipeline_r[17] <= 1'h0;
			pipeline_r[18] <= 1'h0;
			pipeline_r[19] <= 1'h0;
		end
		else if (clk_en) begin
			pipeline_r[0] <= in_;
			pipeline_r[1] <= pipeline_r[5'h00];
			pipeline_r[2] <= pipeline_r[5'h01];
			pipeline_r[3] <= pipeline_r[5'h02];
			pipeline_r[4] <= pipeline_r[5'h03];
			pipeline_r[5] <= pipeline_r[5'h04];
			pipeline_r[6] <= pipeline_r[5'h05];
			pipeline_r[7] <= pipeline_r[5'h06];
			pipeline_r[8] <= pipeline_r[5'h07];
			pipeline_r[9] <= pipeline_r[5'h08];
			pipeline_r[10] <= pipeline_r[5'h09];
			pipeline_r[11] <= pipeline_r[5'h0a];
			pipeline_r[12] <= pipeline_r[5'h0b];
			pipeline_r[13] <= pipeline_r[5'h0c];
			pipeline_r[14] <= pipeline_r[5'h0d];
			pipeline_r[15] <= pipeline_r[5'h0e];
			pipeline_r[16] <= pipeline_r[5'h0f];
			pipeline_r[17] <= pipeline_r[5'h10];
			pipeline_r[18] <= pipeline_r[5'h11];
			pipeline_r[19] <= pipeline_r[5'h12];
		end
endmodule
module pipeline_w_1_d_22_array (
	clk,
	clk_en,
	in_,
	reset,
	out_
);
	input wire clk;
	input wire clk_en;
	input wire in_;
	input wire reset;
	output wire [21:0] out_;
	reg [21:0] pipeline_r;
	assign out_ = pipeline_r;
	always @(posedge clk or posedge reset)
		if (reset) begin
			pipeline_r[0] <= 1'h0;
			pipeline_r[1] <= 1'h0;
			pipeline_r[2] <= 1'h0;
			pipeline_r[3] <= 1'h0;
			pipeline_r[4] <= 1'h0;
			pipeline_r[5] <= 1'h0;
			pipeline_r[6] <= 1'h0;
			pipeline_r[7] <= 1'h0;
			pipeline_r[8] <= 1'h0;
			pipeline_r[9] <= 1'h0;
			pipeline_r[10] <= 1'h0;
			pipeline_r[11] <= 1'h0;
			pipeline_r[12] <= 1'h0;
			pipeline_r[13] <= 1'h0;
			pipeline_r[14] <= 1'h0;
			pipeline_r[15] <= 1'h0;
			pipeline_r[16] <= 1'h0;
			pipeline_r[17] <= 1'h0;
			pipeline_r[18] <= 1'h0;
			pipeline_r[19] <= 1'h0;
			pipeline_r[20] <= 1'h0;
			pipeline_r[21] <= 1'h0;
		end
		else if (clk_en) begin
			pipeline_r[0] <= in_;
			pipeline_r[1] <= pipeline_r[5'h00];
			pipeline_r[2] <= pipeline_r[5'h01];
			pipeline_r[3] <= pipeline_r[5'h02];
			pipeline_r[4] <= pipeline_r[5'h03];
			pipeline_r[5] <= pipeline_r[5'h04];
			pipeline_r[6] <= pipeline_r[5'h05];
			pipeline_r[7] <= pipeline_r[5'h06];
			pipeline_r[8] <= pipeline_r[5'h07];
			pipeline_r[9] <= pipeline_r[5'h08];
			pipeline_r[10] <= pipeline_r[5'h09];
			pipeline_r[11] <= pipeline_r[5'h0a];
			pipeline_r[12] <= pipeline_r[5'h0b];
			pipeline_r[13] <= pipeline_r[5'h0c];
			pipeline_r[14] <= pipeline_r[5'h0d];
			pipeline_r[15] <= pipeline_r[5'h0e];
			pipeline_r[16] <= pipeline_r[5'h0f];
			pipeline_r[17] <= pipeline_r[5'h10];
			pipeline_r[18] <= pipeline_r[5'h11];
			pipeline_r[19] <= pipeline_r[5'h12];
			pipeline_r[20] <= pipeline_r[5'h13];
			pipeline_r[21] <= pipeline_r[5'h14];
		end
endmodule
module pipeline_w_1_d_24_array (
	clk,
	clk_en,
	in_,
	reset,
	out_
);
	input wire clk;
	input wire clk_en;
	input wire in_;
	input wire reset;
	output wire [23:0] out_;
	reg [23:0] pipeline_r;
	assign out_ = pipeline_r;
	always @(posedge clk or posedge reset)
		if (reset) begin
			pipeline_r[0] <= 1'h0;
			pipeline_r[1] <= 1'h0;
			pipeline_r[2] <= 1'h0;
			pipeline_r[3] <= 1'h0;
			pipeline_r[4] <= 1'h0;
			pipeline_r[5] <= 1'h0;
			pipeline_r[6] <= 1'h0;
			pipeline_r[7] <= 1'h0;
			pipeline_r[8] <= 1'h0;
			pipeline_r[9] <= 1'h0;
			pipeline_r[10] <= 1'h0;
			pipeline_r[11] <= 1'h0;
			pipeline_r[12] <= 1'h0;
			pipeline_r[13] <= 1'h0;
			pipeline_r[14] <= 1'h0;
			pipeline_r[15] <= 1'h0;
			pipeline_r[16] <= 1'h0;
			pipeline_r[17] <= 1'h0;
			pipeline_r[18] <= 1'h0;
			pipeline_r[19] <= 1'h0;
			pipeline_r[20] <= 1'h0;
			pipeline_r[21] <= 1'h0;
			pipeline_r[22] <= 1'h0;
			pipeline_r[23] <= 1'h0;
		end
		else if (clk_en) begin
			pipeline_r[0] <= in_;
			pipeline_r[1] <= pipeline_r[5'h00];
			pipeline_r[2] <= pipeline_r[5'h01];
			pipeline_r[3] <= pipeline_r[5'h02];
			pipeline_r[4] <= pipeline_r[5'h03];
			pipeline_r[5] <= pipeline_r[5'h04];
			pipeline_r[6] <= pipeline_r[5'h05];
			pipeline_r[7] <= pipeline_r[5'h06];
			pipeline_r[8] <= pipeline_r[5'h07];
			pipeline_r[9] <= pipeline_r[5'h08];
			pipeline_r[10] <= pipeline_r[5'h09];
			pipeline_r[11] <= pipeline_r[5'h0a];
			pipeline_r[12] <= pipeline_r[5'h0b];
			pipeline_r[13] <= pipeline_r[5'h0c];
			pipeline_r[14] <= pipeline_r[5'h0d];
			pipeline_r[15] <= pipeline_r[5'h0e];
			pipeline_r[16] <= pipeline_r[5'h0f];
			pipeline_r[17] <= pipeline_r[5'h10];
			pipeline_r[18] <= pipeline_r[5'h11];
			pipeline_r[19] <= pipeline_r[5'h12];
			pipeline_r[20] <= pipeline_r[5'h13];
			pipeline_r[21] <= pipeline_r[5'h14];
			pipeline_r[22] <= pipeline_r[5'h15];
			pipeline_r[23] <= pipeline_r[5'h16];
		end
endmodule
module pipeline_w_1_d_5 (
	clk,
	clk_en,
	in_,
	reset,
	out_
);
	input wire clk;
	input wire clk_en;
	input wire in_;
	input wire reset;
	output wire out_;
	reg pipeline_r [4:0];
	assign out_ = pipeline_r[4];
	always @(posedge clk or posedge reset)
		if (reset) begin
			pipeline_r[0] <= 1'h0;
			pipeline_r[1] <= 1'h0;
			pipeline_r[2] <= 1'h0;
			pipeline_r[3] <= 1'h0;
			pipeline_r[4] <= 1'h0;
		end
		else if (clk_en) begin
			pipeline_r[0] <= in_;
			pipeline_r[1] <= pipeline_r[3'h0];
			pipeline_r[2] <= pipeline_r[3'h1];
			pipeline_r[3] <= pipeline_r[3'h2];
			pipeline_r[4] <= pipeline_r[3'h3];
		end
endmodule
module pipeline_w_2_d_1 (
	clk,
	clk_en,
	in_,
	reset,
	out_
);
	input wire clk;
	input wire clk_en;
	input wire [1:0] in_;
	input wire reset;
	output wire [1:0] out_;
	reg [1:0] pipeline_r [0:0];
	assign out_ = pipeline_r[0];
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	always @(posedge clk or posedge reset)
		if (reset) begin : sv2v_autoblock_1
			reg [31:0] i;
			for (i = 0; i < 1; i = i + 1)
				pipeline_r[sv2v_cast_1(i)] <= 2'h0;
		end
		else if (clk_en) begin : sv2v_autoblock_2
			reg [31:0] i;
			for (i = 0; i < 1; i = i + 1)
				if (i == 32'h00000000)
					pipeline_r[sv2v_cast_1(i)] <= in_;
				else
					pipeline_r[sv2v_cast_1(i)] <= pipeline_r[sv2v_cast_1(i - 32'h00000001)];
		end
endmodule
module pipeline_w_2_d_2 (
	clk,
	clk_en,
	in_,
	reset,
	out_
);
	input wire clk;
	input wire clk_en;
	input wire [1:0] in_;
	input wire reset;
	output wire [1:0] out_;
	reg [1:0] pipeline_r [1:0];
	assign out_ = pipeline_r[1];
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	always @(posedge clk or posedge reset)
		if (reset) begin : sv2v_autoblock_1
			reg [31:0] i;
			for (i = 0; i < 2; i = i + 1)
				pipeline_r[sv2v_cast_1(i)] <= 2'h0;
		end
		else if (clk_en) begin : sv2v_autoblock_2
			reg [31:0] i;
			for (i = 0; i < 2; i = i + 1)
				if (i == 32'h00000000)
					pipeline_r[sv2v_cast_1(i)] <= in_;
				else
					pipeline_r[sv2v_cast_1(i)] <= pipeline_r[sv2v_cast_1(i - 32'h00000001)];
		end
endmodule
module pipeline_w_2_d_22_array (
	clk,
	clk_en,
	in_,
	reset,
	out_
);
	input wire clk;
	input wire clk_en;
	input wire [1:0] in_;
	input wire reset;
	output wire [43:0] out_;
	reg [43:0] pipeline_r;
	assign out_ = pipeline_r;
	function automatic [4:0] sv2v_cast_5;
		input reg [4:0] inp;
		sv2v_cast_5 = inp;
	endfunction
	always @(posedge clk or posedge reset)
		if (reset) begin : sv2v_autoblock_1
			reg [31:0] i;
			for (i = 0; i < 22; i = i + 1)
				pipeline_r[sv2v_cast_5(i) * 2+:2] <= 2'h0;
		end
		else if (clk_en) begin : sv2v_autoblock_2
			reg [31:0] i;
			for (i = 0; i < 22; i = i + 1)
				if (i == 32'h00000000)
					pipeline_r[sv2v_cast_5(i) * 2+:2] <= in_;
				else
					pipeline_r[sv2v_cast_5(i) * 2+:2] <= pipeline_r[sv2v_cast_5(i - 32'h00000001) * 2+:2];
		end
endmodule
module pipeline_w_4_d_2 (
	clk,
	clk_en,
	in_,
	reset,
	out_
);
	input wire clk;
	input wire clk_en;
	input wire [3:0] in_;
	input wire reset;
	output wire [3:0] out_;
	reg [3:0] pipeline_r [1:0];
	assign out_ = pipeline_r[1];
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	always @(posedge clk or posedge reset)
		if (reset) begin : sv2v_autoblock_1
			reg [31:0] i;
			for (i = 0; i < 2; i = i + 1)
				pipeline_r[sv2v_cast_1(i)] <= 4'h0;
		end
		else if (clk_en) begin : sv2v_autoblock_2
			reg [31:0] i;
			for (i = 0; i < 2; i = i + 1)
				if (i == 32'h00000000)
					pipeline_r[sv2v_cast_1(i)] <= in_;
				else
					pipeline_r[sv2v_cast_1(i)] <= pipeline_r[sv2v_cast_1(i - 32'h00000001)];
		end
endmodule
module pipeline_w_64_d_0 (
	clk,
	clk_en,
	in_,
	reset,
	out_
);
	input wire clk;
	input wire clk_en;
	input wire [63:0] in_;
	input wire reset;
	output wire [63:0] out_;
	assign out_ = in_;
endmodule
module pipeline_w_65_d_1 (
	clk,
	clk_en,
	in_,
	reset,
	out_
);
	input wire clk;
	input wire clk_en;
	input wire [64:0] in_;
	input wire reset;
	output wire [64:0] out_;
	reg [64:0] pipeline_r [0:0];
	assign out_ = pipeline_r[0];
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	always @(posedge clk or posedge reset)
		if (reset) begin : sv2v_autoblock_1
			reg [31:0] i;
			for (i = 0; i < 1; i = i + 1)
				pipeline_r[sv2v_cast_1(i)] <= 65'h00000000000000000;
		end
		else if (clk_en) begin : sv2v_autoblock_2
			reg [31:0] i;
			for (i = 0; i < 1; i = i + 1)
				if (i == 32'h00000000)
					pipeline_r[sv2v_cast_1(i)] <= in_;
				else
					pipeline_r[sv2v_cast_1(i)] <= pipeline_r[sv2v_cast_1(i - 32'h00000001)];
		end
endmodule
module pipeline_w_74_d_0_reset_high (
	clk,
	clk_en,
	in_,
	reset,
	out_
);
	input wire clk;
	input wire clk_en;
	input wire [73:0] in_;
	input wire reset;
	output wire [73:0] out_;
	assign out_ = in_;
endmodule
module pipeline_w_78_d_0 (
	clk,
	clk_en,
	in_,
	reset,
	out_
);
	input wire clk;
	input wire clk_en;
	input wire [77:0] in_;
	input wire reset;
	output wire [77:0] out_;
	assign out_ = in_;
endmodule
module pipeline_w_90_d_0 (
	clk,
	clk_en,
	in_,
	reset,
	out_
);
	input wire clk;
	input wire clk_en;
	input wire [89:0] in_;
	input wire reset;
	output wire [89:0] out_;
	assign out_ = in_;
endmodule
module reg_fifo_d_19_w_16 (
	almost_empty_diff,
	almost_full_diff,
	clk,
	clk_en,
	data_in,
	flush,
	pop,
	push,
	reset,
	almost_empty,
	almost_full,
	data_out,
	empty,
	full
);
	parameter data_width = 16'h0010;
	input wire [4:0] almost_empty_diff;
	input wire [4:0] almost_full_diff;
	input wire clk;
	input wire clk_en;
	input wire [data_width - 1:0] data_in;
	input wire flush;
	input wire pop;
	input wire push;
	input wire reset;
	output reg almost_empty;
	output reg almost_full;
	output reg [data_width - 1:0] data_out;
	output wire empty;
	output wire full;
	reg [5:0] num_items;
	reg [4:0] rd_ptr;
	wire read;
	reg [(19 * data_width) - 1:0] reg_array;
	reg [4:0] wr_ptr;
	wire write;
	assign full = num_items == 6'h13;
	assign empty = num_items == 6'h00;
	assign read = pop & ~empty;
	assign write = push & ~full;
	function automatic [5:0] sv2v_cast_6;
		input reg [5:0] inp;
		sv2v_cast_6 = inp;
	endfunction
	always @(*) begin
		almost_full = (6'h13 - sv2v_cast_6(almost_full_diff)) <= num_items;
		almost_empty = sv2v_cast_6(almost_empty_diff) >= num_items;
	end
	always @(posedge clk or posedge reset)
		if (reset)
			num_items <= 6'h00;
		else if (clk_en) begin
			if (flush)
				num_items <= 6'h00;
			else if (write & ~read)
				num_items <= num_items + 6'h01;
			else if (~write & read)
				num_items <= num_items - 6'h01;
			else
				num_items <= num_items;
		end
	always @(posedge clk or posedge reset)
		if (reset)
			reg_array <= 304'h0;
		else if (clk_en) begin
			if (write)
				reg_array[wr_ptr * data_width+:data_width] <= data_in;
		end
	always @(posedge clk or posedge reset)
		if (reset)
			wr_ptr <= 5'h00;
		else if (clk_en) begin
			if (flush)
				wr_ptr <= 5'h00;
			else if (write) begin
				if (wr_ptr == 5'h12)
					wr_ptr <= 5'h00;
				else
					wr_ptr <= wr_ptr + 5'h01;
			end
		end
	always @(posedge clk or posedge reset)
		if (reset)
			rd_ptr <= 5'h00;
		else if (clk_en) begin
			if (flush)
				rd_ptr <= 5'h00;
			else if (read) begin
				if (rd_ptr == 5'h12)
					rd_ptr <= 5'h00;
				else
					rd_ptr <= rd_ptr + 5'h01;
			end
		end
	always @(*) data_out = reg_array[rd_ptr * data_width+:data_width];
endmodule
module reg_fifo_d_2_w_16 (
	almost_empty_diff,
	almost_full_diff,
	clk,
	clk_en,
	data_in,
	flush,
	pop,
	push,
	reset,
	almost_empty,
	almost_full,
	data_out,
	empty,
	full
);
	parameter data_width = 16'h0010;
	input wire almost_empty_diff;
	input wire almost_full_diff;
	input wire clk;
	input wire clk_en;
	input wire [data_width - 1:0] data_in;
	input wire flush;
	input wire pop;
	input wire push;
	input wire reset;
	output reg almost_empty;
	output reg almost_full;
	output reg [data_width - 1:0] data_out;
	output wire empty;
	output wire full;
	reg [1:0] num_items;
	reg rd_ptr;
	wire read;
	reg [(2 * data_width) - 1:0] reg_array;
	reg wr_ptr;
	wire write;
	assign full = num_items == 2'h2;
	assign empty = num_items == 2'h0;
	assign read = pop & ~empty;
	assign write = push & ~full;
	function automatic [1:0] sv2v_cast_2;
		input reg [1:0] inp;
		sv2v_cast_2 = inp;
	endfunction
	always @(*) begin
		almost_full = (2'h2 - sv2v_cast_2(almost_full_diff)) <= num_items;
		almost_empty = sv2v_cast_2(almost_empty_diff) >= num_items;
	end
	always @(posedge clk or posedge reset)
		if (reset)
			num_items <= 2'h0;
		else if (clk_en) begin
			if (flush)
				num_items <= 2'h0;
			else if (write & ~read)
				num_items <= num_items + 2'h1;
			else if (~write & read)
				num_items <= num_items - 2'h1;
			else
				num_items <= num_items;
		end
	always @(posedge clk or posedge reset)
		if (reset)
			reg_array <= 32'h00000000;
		else if (clk_en) begin
			if (write)
				reg_array[wr_ptr * data_width+:data_width] <= data_in;
		end
	always @(posedge clk or posedge reset)
		if (reset)
			wr_ptr <= 1'h0;
		else if (clk_en) begin
			if (flush)
				wr_ptr <= 1'h0;
			else if (write) begin
				if (wr_ptr == 1'h1)
					wr_ptr <= 1'h0;
				else
					wr_ptr <= wr_ptr + 1'h1;
			end
		end
	always @(posedge clk or posedge reset)
		if (reset)
			rd_ptr <= 1'h0;
		else if (clk_en) begin
			if (flush)
				rd_ptr <= 1'h0;
			else if (read) begin
				if (rd_ptr == 1'h1)
					rd_ptr <= 1'h0;
				else
					rd_ptr <= rd_ptr + 1'h1;
			end
		end
	always @(*) data_out = reg_array[rd_ptr * data_width+:data_width];
endmodule
module reg_fifo_d_4_w_16 (
	almost_empty_diff,
	almost_full_diff,
	clk,
	clk_en,
	data_in,
	flush,
	pop,
	push,
	reset,
	almost_empty,
	almost_full,
	data_out,
	empty,
	full
);
	parameter data_width = 16'h0010;
	input wire [1:0] almost_empty_diff;
	input wire [1:0] almost_full_diff;
	input wire clk;
	input wire clk_en;
	input wire [data_width - 1:0] data_in;
	input wire flush;
	input wire pop;
	input wire push;
	input wire reset;
	output reg almost_empty;
	output reg almost_full;
	output reg [data_width - 1:0] data_out;
	output wire empty;
	output wire full;
	reg [2:0] num_items;
	reg [1:0] rd_ptr;
	wire read;
	reg [(4 * data_width) - 1:0] reg_array;
	reg [1:0] wr_ptr;
	wire write;
	assign full = num_items == 3'h4;
	assign empty = num_items == 3'h0;
	assign read = pop & ~empty;
	assign write = push & ~full;
	function automatic [2:0] sv2v_cast_3;
		input reg [2:0] inp;
		sv2v_cast_3 = inp;
	endfunction
	always @(*) begin
		almost_full = (3'h4 - sv2v_cast_3(almost_full_diff)) <= num_items;
		almost_empty = sv2v_cast_3(almost_empty_diff) >= num_items;
	end
	always @(posedge clk or posedge reset)
		if (reset)
			num_items <= 3'h0;
		else if (clk_en) begin
			if (flush)
				num_items <= 3'h0;
			else if (write & ~read)
				num_items <= num_items + 3'h1;
			else if (~write & read)
				num_items <= num_items - 3'h1;
			else
				num_items <= num_items;
		end
	always @(posedge clk or posedge reset)
		if (reset)
			reg_array <= 64'h0000000000000000;
		else if (clk_en) begin
			if (write)
				reg_array[wr_ptr * data_width+:data_width] <= data_in;
		end
	always @(posedge clk or posedge reset)
		if (reset)
			wr_ptr <= 2'h0;
		else if (clk_en) begin
			if (flush)
				wr_ptr <= 2'h0;
			else if (write) begin
				if (wr_ptr == 2'h3)
					wr_ptr <= 2'h0;
				else
					wr_ptr <= wr_ptr + 2'h1;
			end
		end
	always @(posedge clk or posedge reset)
		if (reset)
			rd_ptr <= 2'h0;
		else if (clk_en) begin
			if (flush)
				rd_ptr <= 2'h0;
			else if (read) begin
				if (rd_ptr == 2'h3)
					rd_ptr <= 2'h0;
				else
					rd_ptr <= rd_ptr + 2'h1;
			end
		end
	always @(*) data_out = reg_array[rd_ptr * data_width+:data_width];
endmodule
module coreir_wrap (
	in,
	out
);
	input in;
	output wire out;
	assign out = in;
endmodule
module coreir_ult (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output wire out;
	assign out = in0 < in1;
endmodule
module coreir_reg (
	clk,
	in,
	out
);
	parameter width = 1;
	parameter clk_posedge = 1;
	parameter init = 1;
	input clk;
	input [width - 1:0] in;
	output wire [width - 1:0] out;
	reg [width - 1:0] outReg = init;
	wire real_clk;
	assign real_clk = (clk_posedge ? clk : ~clk);
	always @(posedge real_clk) outReg <= in;
	assign out = outReg;
endmodule
module coreir_orr (
	in,
	out
);
	parameter width = 1;
	input [width - 1:0] in;
	output wire out;
	assign out = |in;
endmodule
module coreir_or (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output wire [width - 1:0] out;
	assign out = in0 | in1;
endmodule
module coreir_not (
	in,
	out
);
	parameter width = 1;
	input [width - 1:0] in;
	output wire [width - 1:0] out;
	assign out = ~in;
endmodule
module coreir_mux (
	in0,
	in1,
	sel,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	input sel;
	output wire [width - 1:0] out;
	assign out = (sel ? in1 : in0);
endmodule
module coreir_eq (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output wire out;
	assign out = in0 == in1;
endmodule
module coreir_const (out);
	parameter width = 1;
	parameter value = 1;
	output wire [width - 1:0] out;
	assign out = value;
endmodule
module coreir_andr (
	in,
	out
);
	parameter width = 1;
	input [width - 1:0] in;
	output wire out;
	assign out = &in;
endmodule
module coreir_and (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output wire [width - 1:0] out;
	assign out = in0 & in1;
endmodule
module corebit_const (out);
	parameter value = 1;
	output wire out;
	assign out = value;
endmodule
module corebit_and (
	in0,
	in1,
	out
);
	input in0;
	input in1;
	output wire out;
	assign out = in0 & in1;
endmodule
module and_cell (
	A,
	B,
	Z
);
	input A;
	input B;
	output wire Z;
	AN_CELL inst(
		.A1(A),
		.A2(B),
		.Z(Z)
	);
endmodule
module SplitFifo_17 (
	clk,
	clk_en,
	data_in,
	end_fifo,
	fifo_en,
	ready1,
	rst,
	start_fifo,
	valid0,
	data_out,
	ready0,
	valid1
);
	input wire clk;
	input wire clk_en;
	input wire [16:0] data_in;
	input wire end_fifo;
	input wire fifo_en;
	input wire ready1;
	input wire rst;
	input wire start_fifo;
	input wire valid0;
	output wire [16:0] data_out;
	output wire ready0;
	output wire valid1;
	wire empty;
	reg empty_n;
	wire ready_in;
	wire valid_in;
	reg [16:0] value;
	assign empty = ~empty_n;
	assign ready_in = ready1 && ~start_fifo;
	assign ready0 = (fifo_en ? empty || ready_in : clk_en);
	assign valid_in = valid0 && ~end_fifo;
	assign valid1 = (fifo_en ? ~empty || valid_in : clk_en);
	assign data_out = (empty && fifo_en ? data_in : value);
	always @(posedge clk or posedge rst)
		if (rst)
			value <= 17'h00000;
		else if (clk_en) begin
			if (~fifo_en || ((valid0 && ready0) && ~((empty && ready1) && valid1)))
				value <= data_in;
		end
	always @(posedge clk or posedge rst)
		if (rst)
			empty_n <= 1'h0;
		else if (clk_en) begin
			if (fifo_en) begin
				if (valid1 && ready1) begin
					if (~(valid0 && ready0))
						empty_n <= 1'h0;
				end
				else if (valid0 && ready0)
					empty_n <= 1'h1;
			end
		end
endmodule
module SplitFifo_1 (
	clk,
	clk_en,
	data_in,
	end_fifo,
	fifo_en,
	ready1,
	rst,
	start_fifo,
	valid0,
	data_out,
	ready0,
	valid1
);
	input wire clk;
	input wire clk_en;
	input wire data_in;
	input wire end_fifo;
	input wire fifo_en;
	input wire ready1;
	input wire rst;
	input wire start_fifo;
	input wire valid0;
	output wire data_out;
	output wire ready0;
	output wire valid1;
	wire empty;
	reg empty_n;
	wire ready_in;
	wire valid_in;
	reg value;
	assign empty = ~empty_n;
	assign ready_in = ready1 && ~start_fifo;
	assign ready0 = (fifo_en ? empty || ready_in : clk_en);
	assign valid_in = valid0 && ~end_fifo;
	assign valid1 = (fifo_en ? ~empty || valid_in : clk_en);
	assign data_out = (empty && fifo_en ? data_in : value);
	always @(posedge clk or posedge rst)
		if (rst)
			value <= 1'h0;
		else if (clk_en) begin
			if (~fifo_en || ((valid0 && ready0) && ~((empty && ready1) && valid1)))
				value <= data_in;
		end
	always @(posedge clk or posedge rst)
		if (rst)
			empty_n <= 1'h0;
		else if (clk_en) begin
			if (fifo_en) begin
				if (valid1 && ready1) begin
					if (~(valid0 && ready0))
						empty_n <= 1'h0;
				end
				else if (valid0 && ready0)
					empty_n <= 1'h1;
			end
		end
endmodule
module SliceWrapper_6_1_6 (
	I,
	O
);
	input [5:0] I;
	output wire [4:0] O;
	assign O = I[5:1];
endmodule
module SliceWrapper_6_0_1 (
	I,
	O
);
	input [5:0] I;
	output wire [0:0] O;
	assign O = I[0:0];
endmodule
module SliceWrapper_32_9_10 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[9:9];
endmodule
module SliceWrapper_32_8_9 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[8:8];
endmodule
module SliceWrapper_32_7_8 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[7:7];
endmodule
module SliceWrapper_32_6_7 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[6:6];
endmodule
module SliceWrapper_32_5_6 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[5:5];
endmodule
module SliceWrapper_32_4_5 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[4:4];
endmodule
module SliceWrapper_32_3_4 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[3:3];
endmodule
module SliceWrapper_32_31_32 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[31:31];
endmodule
module SliceWrapper_32_30_31 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[30:30];
endmodule
module SliceWrapper_32_2_3 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[2:2];
endmodule
module SliceWrapper_32_29_30 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[29:29];
endmodule
module SliceWrapper_32_28_31 (
	I,
	O
);
	input [31:0] I;
	output wire [2:0] O;
	assign O = I[30:28];
endmodule
module SliceWrapper_32_28_29 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[28:28];
endmodule
module SliceWrapper_32_27_28 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[27:27];
endmodule
module SliceWrapper_32_26_27 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[26:26];
endmodule
module SliceWrapper_32_25_26 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[25:25];
endmodule
module SliceWrapper_32_24_25 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[24:24];
endmodule
module SliceWrapper_32_23_26 (
	I,
	O
);
	input [31:0] I;
	output wire [2:0] O;
	assign O = I[25:23];
endmodule
module SliceWrapper_32_23_24 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[23:23];
endmodule
module SliceWrapper_32_22_23 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[22:22];
endmodule
module SliceWrapper_32_21_22 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[21:21];
endmodule
module SliceWrapper_32_20_21 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[20:20];
endmodule
module SliceWrapper_32_1_2 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[1:1];
endmodule
module SliceWrapper_32_19_20 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[19:19];
endmodule
module SliceWrapper_32_18_21 (
	I,
	O
);
	input [31:0] I;
	output wire [2:0] O;
	assign O = I[20:18];
endmodule
module SliceWrapper_32_18_19 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[18:18];
endmodule
module SliceWrapper_32_17_18 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[17:17];
endmodule
module SliceWrapper_32_16_17 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[16:16];
endmodule
module SliceWrapper_32_15_16 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[15:15];
endmodule
module SliceWrapper_32_14_15 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[14:14];
endmodule
module SliceWrapper_32_13_14 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[13:13];
endmodule
module SliceWrapper_32_12_13 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[12:12];
endmodule
module SliceWrapper_32_11_12 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[11:11];
endmodule
module SliceWrapper_32_10_11 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[10:10];
endmodule
module SliceWrapper_32_0_32 (
	I,
	O
);
	input [31:0] I;
	output wire [31:0] O;
	assign O = I;
endmodule
module SliceWrapper_32_0_22 (
	I,
	O
);
	input [31:0] I;
	output wire [21:0] O;
	assign O = I[21:0];
endmodule
module SliceWrapper_32_0_1 (
	I,
	O
);
	input [31:0] I;
	output wire [0:0] O;
	assign O = I[0:0];
endmodule
module SliceWrapper_31_9_10 (
	I,
	O
);
	input [30:0] I;
	output wire [0:0] O;
	assign O = I[9:9];
endmodule
module SliceWrapper_31_6_9 (
	I,
	O
);
	input [30:0] I;
	output wire [2:0] O;
	assign O = I[8:6];
endmodule
module SliceWrapper_31_5_6 (
	I,
	O
);
	input [30:0] I;
	output wire [0:0] O;
	assign O = I[5:5];
endmodule
module SliceWrapper_31_4_5 (
	I,
	O
);
	input [30:0] I;
	output wire [0:0] O;
	assign O = I[4:4];
endmodule
module SliceWrapper_31_30_31 (
	I,
	O
);
	input [30:0] I;
	output wire [0:0] O;
	assign O = I[30:30];
endmodule
module SliceWrapper_31_29_30 (
	I,
	O
);
	input [30:0] I;
	output wire [0:0] O;
	assign O = I[29:29];
endmodule
module SliceWrapper_31_26_29 (
	I,
	O
);
	input [30:0] I;
	output wire [2:0] O;
	assign O = I[28:26];
endmodule
module SliceWrapper_31_25_26 (
	I,
	O
);
	input [30:0] I;
	output wire [0:0] O;
	assign O = I[25:25];
endmodule
module SliceWrapper_31_24_25 (
	I,
	O
);
	input [30:0] I;
	output wire [0:0] O;
	assign O = I[24:24];
endmodule
module SliceWrapper_31_21_24 (
	I,
	O
);
	input [30:0] I;
	output wire [2:0] O;
	assign O = I[23:21];
endmodule
module SliceWrapper_31_20_21 (
	I,
	O
);
	input [30:0] I;
	output wire [0:0] O;
	assign O = I[20:20];
endmodule
module SliceWrapper_31_1_4 (
	I,
	O
);
	input [30:0] I;
	output wire [2:0] O;
	assign O = I[3:1];
endmodule
module SliceWrapper_31_19_20 (
	I,
	O
);
	input [30:0] I;
	output wire [0:0] O;
	assign O = I[19:19];
endmodule
module SliceWrapper_31_16_19 (
	I,
	O
);
	input [30:0] I;
	output wire [2:0] O;
	assign O = I[18:16];
endmodule
module SliceWrapper_31_15_16 (
	I,
	O
);
	input [30:0] I;
	output wire [0:0] O;
	assign O = I[15:15];
endmodule
module SliceWrapper_31_14_15 (
	I,
	O
);
	input [30:0] I;
	output wire [0:0] O;
	assign O = I[14:14];
endmodule
module SliceWrapper_31_11_14 (
	I,
	O
);
	input [30:0] I;
	output wire [2:0] O;
	assign O = I[13:11];
endmodule
module SliceWrapper_31_10_11 (
	I,
	O
);
	input [30:0] I;
	output wire [0:0] O;
	assign O = I[10:10];
endmodule
module SliceWrapper_31_0_1 (
	I,
	O
);
	input [30:0] I;
	output wire [0:0] O;
	assign O = I[0:0];
endmodule
module SliceWrapper_30_9_10 (
	I,
	O
);
	input [29:0] I;
	output wire [0:0] O;
	assign O = I[9:9];
endmodule
module SliceWrapper_30_8_9 (
	I,
	O
);
	input [29:0] I;
	output wire [0:0] O;
	assign O = I[8:8];
endmodule
module SliceWrapper_30_5_8 (
	I,
	O
);
	input [29:0] I;
	output wire [2:0] O;
	assign O = I[7:5];
endmodule
module SliceWrapper_30_4_5 (
	I,
	O
);
	input [29:0] I;
	output wire [0:0] O;
	assign O = I[4:4];
endmodule
module SliceWrapper_30_3_4 (
	I,
	O
);
	input [29:0] I;
	output wire [0:0] O;
	assign O = I[3:3];
endmodule
module SliceWrapper_30_29_30 (
	I,
	O
);
	input [29:0] I;
	output wire [0:0] O;
	assign O = I[29:29];
endmodule
module SliceWrapper_30_28_29 (
	I,
	O
);
	input [29:0] I;
	output wire [0:0] O;
	assign O = I[28:28];
endmodule
module SliceWrapper_30_25_28 (
	I,
	O
);
	input [29:0] I;
	output wire [2:0] O;
	assign O = I[27:25];
endmodule
module SliceWrapper_30_24_25 (
	I,
	O
);
	input [29:0] I;
	output wire [0:0] O;
	assign O = I[24:24];
endmodule
module SliceWrapper_30_23_24 (
	I,
	O
);
	input [29:0] I;
	output wire [0:0] O;
	assign O = I[23:23];
endmodule
module SliceWrapper_30_20_23 (
	I,
	O
);
	input [29:0] I;
	output wire [2:0] O;
	assign O = I[22:20];
endmodule
module SliceWrapper_30_19_20 (
	I,
	O
);
	input [29:0] I;
	output wire [0:0] O;
	assign O = I[19:19];
endmodule
module SliceWrapper_30_18_19 (
	I,
	O
);
	input [29:0] I;
	output wire [0:0] O;
	assign O = I[18:18];
endmodule
module SliceWrapper_30_15_18 (
	I,
	O
);
	input [29:0] I;
	output wire [2:0] O;
	assign O = I[17:15];
endmodule
module SliceWrapper_30_14_15 (
	I,
	O
);
	input [29:0] I;
	output wire [0:0] O;
	assign O = I[14:14];
endmodule
module SliceWrapper_30_13_14 (
	I,
	O
);
	input [29:0] I;
	output wire [0:0] O;
	assign O = I[13:13];
endmodule
module SliceWrapper_30_10_13 (
	I,
	O
);
	input [29:0] I;
	output wire [2:0] O;
	assign O = I[12:10];
endmodule
module SliceWrapper_30_0_30 (
	I,
	O
);
	input [29:0] I;
	output wire [29:0] O;
	assign O = I;
endmodule
module SliceWrapper_30_0_3 (
	I,
	O
);
	input [29:0] I;
	output wire [2:0] O;
	assign O = I[2:0];
endmodule
module SliceWrapper_25_9_10 (
	I,
	O
);
	input [24:0] I;
	output wire [0:0] O;
	assign O = I[9:9];
endmodule
module SliceWrapper_25_8_9 (
	I,
	O
);
	input [24:0] I;
	output wire [0:0] O;
	assign O = I[8:8];
endmodule
module SliceWrapper_25_7_8 (
	I,
	O
);
	input [24:0] I;
	output wire [0:0] O;
	assign O = I[7:7];
endmodule
module SliceWrapper_25_6_7 (
	I,
	O
);
	input [24:0] I;
	output wire [0:0] O;
	assign O = I[6:6];
endmodule
module SliceWrapper_25_5_6 (
	I,
	O
);
	input [24:0] I;
	output wire [0:0] O;
	assign O = I[5:5];
endmodule
module SliceWrapper_25_4_5 (
	I,
	O
);
	input [24:0] I;
	output wire [0:0] O;
	assign O = I[4:4];
endmodule
module SliceWrapper_25_3_4 (
	I,
	O
);
	input [24:0] I;
	output wire [0:0] O;
	assign O = I[3:3];
endmodule
module SliceWrapper_25_2_3 (
	I,
	O
);
	input [24:0] I;
	output wire [0:0] O;
	assign O = I[2:2];
endmodule
module SliceWrapper_25_24_25 (
	I,
	O
);
	input [24:0] I;
	output wire [0:0] O;
	assign O = I[24:24];
endmodule
module SliceWrapper_25_23_24 (
	I,
	O
);
	input [24:0] I;
	output wire [0:0] O;
	assign O = I[23:23];
endmodule
module SliceWrapper_25_21_23 (
	I,
	O
);
	input [24:0] I;
	output wire [1:0] O;
	assign O = I[22:21];
endmodule
module SliceWrapper_25_20_21 (
	I,
	O
);
	input [24:0] I;
	output wire [0:0] O;
	assign O = I[20:20];
endmodule
module SliceWrapper_25_1_2 (
	I,
	O
);
	input [24:0] I;
	output wire [0:0] O;
	assign O = I[1:1];
endmodule
module SliceWrapper_25_19_20 (
	I,
	O
);
	input [24:0] I;
	output wire [0:0] O;
	assign O = I[19:19];
endmodule
module SliceWrapper_25_18_19 (
	I,
	O
);
	input [24:0] I;
	output wire [0:0] O;
	assign O = I[18:18];
endmodule
module SliceWrapper_25_17_18 (
	I,
	O
);
	input [24:0] I;
	output wire [0:0] O;
	assign O = I[17:17];
endmodule
module SliceWrapper_25_16_17 (
	I,
	O
);
	input [24:0] I;
	output wire [0:0] O;
	assign O = I[16:16];
endmodule
module SliceWrapper_25_15_16 (
	I,
	O
);
	input [24:0] I;
	output wire [0:0] O;
	assign O = I[15:15];
endmodule
module SliceWrapper_25_14_15 (
	I,
	O
);
	input [24:0] I;
	output wire [0:0] O;
	assign O = I[14:14];
endmodule
module SliceWrapper_25_13_14 (
	I,
	O
);
	input [24:0] I;
	output wire [0:0] O;
	assign O = I[13:13];
endmodule
module SliceWrapper_25_12_13 (
	I,
	O
);
	input [24:0] I;
	output wire [0:0] O;
	assign O = I[12:12];
endmodule
module SliceWrapper_25_11_12 (
	I,
	O
);
	input [24:0] I;
	output wire [0:0] O;
	assign O = I[11:11];
endmodule
module SliceWrapper_25_10_11 (
	I,
	O
);
	input [24:0] I;
	output wire [0:0] O;
	assign O = I[10:10];
endmodule
module SliceWrapper_25_0_1 (
	I,
	O
);
	input [24:0] I;
	output wire [0:0] O;
	assign O = I[0:0];
endmodule
module SliceWrapper_24_9_10 (
	I,
	O
);
	input [23:0] I;
	output wire [0:0] O;
	assign O = I[9:9];
endmodule
module SliceWrapper_24_8_9 (
	I,
	O
);
	input [23:0] I;
	output wire [0:0] O;
	assign O = I[8:8];
endmodule
module SliceWrapper_24_7_8 (
	I,
	O
);
	input [23:0] I;
	output wire [0:0] O;
	assign O = I[7:7];
endmodule
module SliceWrapper_24_6_7 (
	I,
	O
);
	input [23:0] I;
	output wire [0:0] O;
	assign O = I[6:6];
endmodule
module SliceWrapper_24_5_6 (
	I,
	O
);
	input [23:0] I;
	output wire [0:0] O;
	assign O = I[5:5];
endmodule
module SliceWrapper_24_4_5 (
	I,
	O
);
	input [23:0] I;
	output wire [0:0] O;
	assign O = I[4:4];
endmodule
module SliceWrapper_24_3_4 (
	I,
	O
);
	input [23:0] I;
	output wire [0:0] O;
	assign O = I[3:3];
endmodule
module SliceWrapper_24_2_3 (
	I,
	O
);
	input [23:0] I;
	output wire [0:0] O;
	assign O = I[2:2];
endmodule
module SliceWrapper_24_23_24 (
	I,
	O
);
	input [23:0] I;
	output wire [0:0] O;
	assign O = I[23:23];
endmodule
module SliceWrapper_24_22_23 (
	I,
	O
);
	input [23:0] I;
	output wire [0:0] O;
	assign O = I[22:22];
endmodule
module SliceWrapper_24_21_22 (
	I,
	O
);
	input [23:0] I;
	output wire [0:0] O;
	assign O = I[21:21];
endmodule
module SliceWrapper_24_20_21 (
	I,
	O
);
	input [23:0] I;
	output wire [0:0] O;
	assign O = I[20:20];
endmodule
module SliceWrapper_24_1_2 (
	I,
	O
);
	input [23:0] I;
	output wire [0:0] O;
	assign O = I[1:1];
endmodule
module SliceWrapper_24_19_20 (
	I,
	O
);
	input [23:0] I;
	output wire [0:0] O;
	assign O = I[19:19];
endmodule
module SliceWrapper_24_18_19 (
	I,
	O
);
	input [23:0] I;
	output wire [0:0] O;
	assign O = I[18:18];
endmodule
module SliceWrapper_24_17_18 (
	I,
	O
);
	input [23:0] I;
	output wire [0:0] O;
	assign O = I[17:17];
endmodule
module SliceWrapper_24_16_17 (
	I,
	O
);
	input [23:0] I;
	output wire [0:0] O;
	assign O = I[16:16];
endmodule
module SliceWrapper_24_15_16 (
	I,
	O
);
	input [23:0] I;
	output wire [0:0] O;
	assign O = I[15:15];
endmodule
module SliceWrapper_24_14_15 (
	I,
	O
);
	input [23:0] I;
	output wire [0:0] O;
	assign O = I[14:14];
endmodule
module SliceWrapper_24_13_14 (
	I,
	O
);
	input [23:0] I;
	output wire [0:0] O;
	assign O = I[13:13];
endmodule
module SliceWrapper_24_12_13 (
	I,
	O
);
	input [23:0] I;
	output wire [0:0] O;
	assign O = I[12:12];
endmodule
module SliceWrapper_24_11_12 (
	I,
	O
);
	input [23:0] I;
	output wire [0:0] O;
	assign O = I[11:11];
endmodule
module SliceWrapper_24_10_11 (
	I,
	O
);
	input [23:0] I;
	output wire [0:0] O;
	assign O = I[10:10];
endmodule
module SliceWrapper_24_0_1 (
	I,
	O
);
	input [23:0] I;
	output wire [0:0] O;
	assign O = I[0:0];
endmodule
module SliceWrapper_23_9_10 (
	I,
	O
);
	input [22:0] I;
	output wire [0:0] O;
	assign O = I[9:9];
endmodule
module SliceWrapper_23_8_9 (
	I,
	O
);
	input [22:0] I;
	output wire [0:0] O;
	assign O = I[8:8];
endmodule
module SliceWrapper_23_5_8 (
	I,
	O
);
	input [22:0] I;
	output wire [2:0] O;
	assign O = I[7:5];
endmodule
module SliceWrapper_23_4_5 (
	I,
	O
);
	input [22:0] I;
	output wire [0:0] O;
	assign O = I[4:4];
endmodule
module SliceWrapper_23_3_4 (
	I,
	O
);
	input [22:0] I;
	output wire [0:0] O;
	assign O = I[3:3];
endmodule
module SliceWrapper_23_20_23 (
	I,
	O
);
	input [22:0] I;
	output wire [2:0] O;
	assign O = I[22:20];
endmodule
module SliceWrapper_23_19_20 (
	I,
	O
);
	input [22:0] I;
	output wire [0:0] O;
	assign O = I[19:19];
endmodule
module SliceWrapper_23_18_19 (
	I,
	O
);
	input [22:0] I;
	output wire [0:0] O;
	assign O = I[18:18];
endmodule
module SliceWrapper_23_15_18 (
	I,
	O
);
	input [22:0] I;
	output wire [2:0] O;
	assign O = I[17:15];
endmodule
module SliceWrapper_23_14_15 (
	I,
	O
);
	input [22:0] I;
	output wire [0:0] O;
	assign O = I[14:14];
endmodule
module SliceWrapper_23_13_14 (
	I,
	O
);
	input [22:0] I;
	output wire [0:0] O;
	assign O = I[13:13];
endmodule
module SliceWrapper_23_10_13 (
	I,
	O
);
	input [22:0] I;
	output wire [2:0] O;
	assign O = I[12:10];
endmodule
module SliceWrapper_23_0_3 (
	I,
	O
);
	input [22:0] I;
	output wire [2:0] O;
	assign O = I[2:0];
endmodule
module SliceWrapper_20_9_10 (
	I,
	O
);
	input [19:0] I;
	output wire [0:0] O;
	assign O = I[9:9];
endmodule
module SliceWrapper_20_8_9 (
	I,
	O
);
	input [19:0] I;
	output wire [0:0] O;
	assign O = I[8:8];
endmodule
module SliceWrapper_20_7_8 (
	I,
	O
);
	input [19:0] I;
	output wire [0:0] O;
	assign O = I[7:7];
endmodule
module SliceWrapper_20_6_7 (
	I,
	O
);
	input [19:0] I;
	output wire [0:0] O;
	assign O = I[6:6];
endmodule
module SliceWrapper_20_5_6 (
	I,
	O
);
	input [19:0] I;
	output wire [0:0] O;
	assign O = I[5:5];
endmodule
module SliceWrapper_20_4_5 (
	I,
	O
);
	input [19:0] I;
	output wire [0:0] O;
	assign O = I[4:4];
endmodule
module SliceWrapper_20_3_4 (
	I,
	O
);
	input [19:0] I;
	output wire [0:0] O;
	assign O = I[3:3];
endmodule
module SliceWrapper_20_2_3 (
	I,
	O
);
	input [19:0] I;
	output wire [0:0] O;
	assign O = I[2:2];
endmodule
module SliceWrapper_20_1_2 (
	I,
	O
);
	input [19:0] I;
	output wire [0:0] O;
	assign O = I[1:1];
endmodule
module SliceWrapper_20_19_20 (
	I,
	O
);
	input [19:0] I;
	output wire [0:0] O;
	assign O = I[19:19];
endmodule
module SliceWrapper_20_16_19 (
	I,
	O
);
	input [19:0] I;
	output wire [2:0] O;
	assign O = I[18:16];
endmodule
module SliceWrapper_20_15_16 (
	I,
	O
);
	input [19:0] I;
	output wire [0:0] O;
	assign O = I[15:15];
endmodule
module SliceWrapper_20_14_15 (
	I,
	O
);
	input [19:0] I;
	output wire [0:0] O;
	assign O = I[14:14];
endmodule
module SliceWrapper_20_13_14 (
	I,
	O
);
	input [19:0] I;
	output wire [0:0] O;
	assign O = I[13:13];
endmodule
module SliceWrapper_20_12_13 (
	I,
	O
);
	input [19:0] I;
	output wire [0:0] O;
	assign O = I[12:12];
endmodule
module SliceWrapper_20_11_12 (
	I,
	O
);
	input [19:0] I;
	output wire [0:0] O;
	assign O = I[11:11];
endmodule
module SliceWrapper_20_10_11 (
	I,
	O
);
	input [19:0] I;
	output wire [0:0] O;
	assign O = I[10:10];
endmodule
module SliceWrapper_20_0_1 (
	I,
	O
);
	input [19:0] I;
	output wire [0:0] O;
	assign O = I[0:0];
endmodule
module SliceWrapper_1_0_1 (
	I,
	O
);
	input [0:0] I;
	output wire [0:0] O;
	assign O = I;
endmodule
module SliceWrapper_19_0_19 (
	I,
	O
);
	input [18:0] I;
	output wire [18:0] O;
	assign O = I;
endmodule
module SliceWrapper_16_0_16 (
	I,
	O
);
	input [15:0] I;
	output wire [15:0] O;
	assign O = I;
endmodule
module Register_unq9 (
	I,
	O,
	CE,
	CLK,
	ASYNCRESET
);
	input [23:0] I;
	output wire [23:0] O;
	input CE;
	input CLK;
	input ASYNCRESET;
	wire [23:0] reg_PR24_inst0__CE_out;
	regCE_arst #(
		.init(24'h000000),
		.width(24)
	) reg_PR24_inst0__CE(
		.in(I),
		.ce(CE),
		.out(reg_PR24_inst0__CE_out),
		.clk(CLK),
		.arst(ASYNCRESET)
	);
	assign O = reg_PR24_inst0__CE_out;
endmodule
module Register_unq8 (
	I,
	O,
	CE,
	CLK,
	ASYNCRESET
);
	input [24:0] I;
	output wire [24:0] O;
	input CE;
	input CLK;
	input ASYNCRESET;
	wire [24:0] reg_PR25_inst0__CE_out;
	regCE_arst #(
		.init(25'h0000000),
		.width(25)
	) reg_PR25_inst0__CE(
		.in(I),
		.ce(CE),
		.out(reg_PR25_inst0__CE_out),
		.clk(CLK),
		.arst(ASYNCRESET)
	);
	assign O = reg_PR25_inst0__CE_out;
endmodule
module Register_unq7 (
	I,
	O,
	CE,
	CLK,
	ASYNCRESET
);
	input [18:0] I;
	output wire [18:0] O;
	input CE;
	input CLK;
	input ASYNCRESET;
	wire [18:0] reg_PR19_inst0__CE_out;
	regCE_arst #(
		.init(19'h00000),
		.width(19)
	) reg_PR19_inst0__CE(
		.in(I),
		.ce(CE),
		.out(reg_PR19_inst0__CE_out),
		.clk(CLK),
		.arst(ASYNCRESET)
	);
	assign O = reg_PR19_inst0__CE_out;
endmodule
module Register_unq6 (
	I,
	O,
	CE,
	CLK,
	ASYNCRESET
);
	input [22:0] I;
	output wire [22:0] O;
	input CE;
	input CLK;
	input ASYNCRESET;
	wire [22:0] reg_PR23_inst0__CE_out;
	regCE_arst #(
		.init(23'h000000),
		.width(23)
	) reg_PR23_inst0__CE(
		.in(I),
		.ce(CE),
		.out(reg_PR23_inst0__CE_out),
		.clk(CLK),
		.arst(ASYNCRESET)
	);
	assign O = reg_PR23_inst0__CE_out;
endmodule
module Register_unq5 (
	I,
	O,
	CE,
	CLK,
	ASYNCRESET
);
	input [30:0] I;
	output wire [30:0] O;
	input CE;
	input CLK;
	input ASYNCRESET;
	wire [30:0] reg_PR31_inst0__CE_out;
	regCE_arst #(
		.init(31'h00000000),
		.width(31)
	) reg_PR31_inst0__CE(
		.in(I),
		.ce(CE),
		.out(reg_PR31_inst0__CE_out),
		.clk(CLK),
		.arst(ASYNCRESET)
	);
	assign O = reg_PR31_inst0__CE_out;
endmodule
module Register_unq4 (
	I,
	O,
	CE,
	CLK,
	ASYNCRESET
);
	input [0:0] I;
	output wire [0:0] O;
	input CE;
	input CLK;
	input ASYNCRESET;
	wire [0:0] reg_PR1_inst0__CE_out;
	regCE_arst #(
		.init(1'h0),
		.width(1)
	) reg_PR1_inst0__CE(
		.in(I),
		.ce(CE),
		.out(reg_PR1_inst0__CE_out),
		.clk(CLK),
		.arst(ASYNCRESET)
	);
	assign O = reg_PR1_inst0__CE_out;
endmodule
module Register_unq3 (
	I,
	O,
	CE,
	CLK,
	ASYNCRESET
);
	input [29:0] I;
	output wire [29:0] O;
	input CE;
	input CLK;
	input ASYNCRESET;
	wire [29:0] reg_PR30_inst0__CE_out;
	regCE_arst #(
		.init(30'h00000000),
		.width(30)
	) reg_PR30_inst0__CE(
		.in(I),
		.ce(CE),
		.out(reg_PR30_inst0__CE_out),
		.clk(CLK),
		.arst(ASYNCRESET)
	);
	assign O = reg_PR30_inst0__CE_out;
endmodule
module Register_unq2 (
	I,
	O,
	CE,
	CLK,
	ASYNCRESET
);
	input [5:0] I;
	output wire [5:0] O;
	input CE;
	input CLK;
	input ASYNCRESET;
	wire [5:0] reg_PR6_inst0__CE_out;
	regCE_arst #(
		.init(6'h00),
		.width(6)
	) reg_PR6_inst0__CE(
		.in(I),
		.ce(CE),
		.out(reg_PR6_inst0__CE_out),
		.clk(CLK),
		.arst(ASYNCRESET)
	);
	assign O = reg_PR6_inst0__CE_out;
endmodule
module Register_unq1 (
	I,
	O,
	CE,
	CLK,
	ASYNCRESET
);
	input [19:0] I;
	output wire [19:0] O;
	input CE;
	input CLK;
	input ASYNCRESET;
	wire [19:0] reg_PR20_inst0__CE_out;
	regCE_arst #(
		.init(20'h00000),
		.width(20)
	) reg_PR20_inst0__CE(
		.in(I),
		.ce(CE),
		.out(reg_PR20_inst0__CE_out),
		.clk(CLK),
		.arst(ASYNCRESET)
	);
	assign O = reg_PR20_inst0__CE_out;
endmodule
module Register (
	I,
	O,
	CE,
	CLK,
	ASYNCRESET
);
	input [31:0] I;
	output wire [31:0] O;
	input CE;
	input CLK;
	input ASYNCRESET;
	wire [31:0] reg_PR32_inst0__CE_out;
	regCE_arst #(
		.init(32'h00000000),
		.width(32)
	) reg_PR32_inst0__CE(
		.in(I),
		.ce(CE),
		.out(reg_PR32_inst0__CE_out),
		.clk(CLK),
		.arst(ASYNCRESET)
	);
	assign O = reg_PR32_inst0__CE_out;
endmodule
module ReadyValidLoopBack (
	ready_in,
	valid_in,
	valid_out
);
	input wire ready_in;
	input wire valid_in;
	output wire valid_out;
	assign valid_out = ready_in & valid_in;
endmodule
module PowerDomainOR (
	I0,
	I1,
	O,
	I_not
);
	input [31:0] I0;
	input [31:0] I1;
	output wire [31:0] O;
	input [0:0] I_not;
	wire [0:0] Invert1_inst0_out;
	wire [0:0] and1_inst0_out;
	wire [0:0] and1_inst1_out;
	wire [0:0] and1_inst10_out;
	wire [0:0] and1_inst11_out;
	wire [0:0] and1_inst12_out;
	wire [0:0] and1_inst13_out;
	wire [0:0] and1_inst14_out;
	wire [0:0] and1_inst15_out;
	wire [0:0] and1_inst16_out;
	wire [0:0] and1_inst17_out;
	wire [0:0] and1_inst18_out;
	wire [0:0] and1_inst19_out;
	wire [0:0] and1_inst2_out;
	wire [0:0] and1_inst20_out;
	wire [0:0] and1_inst21_out;
	wire [0:0] and1_inst22_out;
	wire [0:0] and1_inst23_out;
	wire [0:0] and1_inst24_out;
	wire [0:0] and1_inst25_out;
	wire [0:0] and1_inst26_out;
	wire [0:0] and1_inst27_out;
	wire [0:0] and1_inst28_out;
	wire [0:0] and1_inst29_out;
	wire [0:0] and1_inst3_out;
	wire [0:0] and1_inst30_out;
	wire [0:0] and1_inst31_out;
	wire [0:0] and1_inst4_out;
	wire [0:0] and1_inst5_out;
	wire [0:0] and1_inst6_out;
	wire [0:0] and1_inst7_out;
	wire [0:0] and1_inst8_out;
	wire [0:0] and1_inst9_out;
	wire [31:0] or32_inst0_out;
	coreir_not #(.width(1)) Invert1_inst0(
		.in(I_not),
		.out(Invert1_inst0_out)
	);
	coreir_and #(.width(1)) and1_inst0(
		.in0(I0[0]),
		.in1(Invert1_inst0_out),
		.out(and1_inst0_out)
	);
	coreir_and #(.width(1)) and1_inst1(
		.in0(I0[1]),
		.in1(Invert1_inst0_out),
		.out(and1_inst1_out)
	);
	coreir_and #(.width(1)) and1_inst10(
		.in0(I0[10]),
		.in1(Invert1_inst0_out),
		.out(and1_inst10_out)
	);
	coreir_and #(.width(1)) and1_inst11(
		.in0(I0[11]),
		.in1(Invert1_inst0_out),
		.out(and1_inst11_out)
	);
	coreir_and #(.width(1)) and1_inst12(
		.in0(I0[12]),
		.in1(Invert1_inst0_out),
		.out(and1_inst12_out)
	);
	coreir_and #(.width(1)) and1_inst13(
		.in0(I0[13]),
		.in1(Invert1_inst0_out),
		.out(and1_inst13_out)
	);
	coreir_and #(.width(1)) and1_inst14(
		.in0(I0[14]),
		.in1(Invert1_inst0_out),
		.out(and1_inst14_out)
	);
	coreir_and #(.width(1)) and1_inst15(
		.in0(I0[15]),
		.in1(Invert1_inst0_out),
		.out(and1_inst15_out)
	);
	coreir_and #(.width(1)) and1_inst16(
		.in0(I0[16]),
		.in1(Invert1_inst0_out),
		.out(and1_inst16_out)
	);
	coreir_and #(.width(1)) and1_inst17(
		.in0(I0[17]),
		.in1(Invert1_inst0_out),
		.out(and1_inst17_out)
	);
	coreir_and #(.width(1)) and1_inst18(
		.in0(I0[18]),
		.in1(Invert1_inst0_out),
		.out(and1_inst18_out)
	);
	coreir_and #(.width(1)) and1_inst19(
		.in0(I0[19]),
		.in1(Invert1_inst0_out),
		.out(and1_inst19_out)
	);
	coreir_and #(.width(1)) and1_inst2(
		.in0(I0[2]),
		.in1(Invert1_inst0_out),
		.out(and1_inst2_out)
	);
	coreir_and #(.width(1)) and1_inst20(
		.in0(I0[20]),
		.in1(Invert1_inst0_out),
		.out(and1_inst20_out)
	);
	coreir_and #(.width(1)) and1_inst21(
		.in0(I0[21]),
		.in1(Invert1_inst0_out),
		.out(and1_inst21_out)
	);
	coreir_and #(.width(1)) and1_inst22(
		.in0(I0[22]),
		.in1(Invert1_inst0_out),
		.out(and1_inst22_out)
	);
	coreir_and #(.width(1)) and1_inst23(
		.in0(I0[23]),
		.in1(Invert1_inst0_out),
		.out(and1_inst23_out)
	);
	coreir_and #(.width(1)) and1_inst24(
		.in0(I0[24]),
		.in1(Invert1_inst0_out),
		.out(and1_inst24_out)
	);
	coreir_and #(.width(1)) and1_inst25(
		.in0(I0[25]),
		.in1(Invert1_inst0_out),
		.out(and1_inst25_out)
	);
	coreir_and #(.width(1)) and1_inst26(
		.in0(I0[26]),
		.in1(Invert1_inst0_out),
		.out(and1_inst26_out)
	);
	coreir_and #(.width(1)) and1_inst27(
		.in0(I0[27]),
		.in1(Invert1_inst0_out),
		.out(and1_inst27_out)
	);
	coreir_and #(.width(1)) and1_inst28(
		.in0(I0[28]),
		.in1(Invert1_inst0_out),
		.out(and1_inst28_out)
	);
	coreir_and #(.width(1)) and1_inst29(
		.in0(I0[29]),
		.in1(Invert1_inst0_out),
		.out(and1_inst29_out)
	);
	coreir_and #(.width(1)) and1_inst3(
		.in0(I0[3]),
		.in1(Invert1_inst0_out),
		.out(and1_inst3_out)
	);
	coreir_and #(.width(1)) and1_inst30(
		.in0(I0[30]),
		.in1(Invert1_inst0_out),
		.out(and1_inst30_out)
	);
	coreir_and #(.width(1)) and1_inst31(
		.in0(I0[31]),
		.in1(Invert1_inst0_out),
		.out(and1_inst31_out)
	);
	coreir_and #(.width(1)) and1_inst4(
		.in0(I0[4]),
		.in1(Invert1_inst0_out),
		.out(and1_inst4_out)
	);
	coreir_and #(.width(1)) and1_inst5(
		.in0(I0[5]),
		.in1(Invert1_inst0_out),
		.out(and1_inst5_out)
	);
	coreir_and #(.width(1)) and1_inst6(
		.in0(I0[6]),
		.in1(Invert1_inst0_out),
		.out(and1_inst6_out)
	);
	coreir_and #(.width(1)) and1_inst7(
		.in0(I0[7]),
		.in1(Invert1_inst0_out),
		.out(and1_inst7_out)
	);
	coreir_and #(.width(1)) and1_inst8(
		.in0(I0[8]),
		.in1(Invert1_inst0_out),
		.out(and1_inst8_out)
	);
	coreir_and #(.width(1)) and1_inst9(
		.in0(I0[9]),
		.in1(Invert1_inst0_out),
		.out(and1_inst9_out)
	);
	wire [31:0] or32_inst0_in0;
	assign or32_inst0_in0 = {and1_inst31_out[0], and1_inst30_out[0], and1_inst29_out[0], and1_inst28_out[0], and1_inst27_out[0], and1_inst26_out[0], and1_inst25_out[0], and1_inst24_out[0], and1_inst23_out[0], and1_inst22_out[0], and1_inst21_out[0], and1_inst20_out[0], and1_inst19_out[0], and1_inst18_out[0], and1_inst17_out[0], and1_inst16_out[0], and1_inst15_out[0], and1_inst14_out[0], and1_inst13_out[0], and1_inst12_out[0], and1_inst11_out[0], and1_inst10_out[0], and1_inst9_out[0], and1_inst8_out[0], and1_inst7_out[0], and1_inst6_out[0], and1_inst5_out[0], and1_inst4_out[0], and1_inst3_out[0], and1_inst2_out[0], and1_inst1_out[0], and1_inst0_out[0]};
	coreir_or #(.width(32)) or32_inst0(
		.in0(or32_inst0_in0),
		.in1(I1),
		.out(or32_inst0_out)
	);
	assign O = or32_inst0_out;
endmodule
module PondTop (
	CONFIG_SPACE_0,
	CONFIG_SPACE_1,
	CONFIG_SPACE_10,
	CONFIG_SPACE_11,
	CONFIG_SPACE_12,
	CONFIG_SPACE_13,
	CONFIG_SPACE_14,
	CONFIG_SPACE_15,
	CONFIG_SPACE_16,
	CONFIG_SPACE_2,
	CONFIG_SPACE_3,
	CONFIG_SPACE_4,
	CONFIG_SPACE_5,
	CONFIG_SPACE_6,
	CONFIG_SPACE_7,
	CONFIG_SPACE_8,
	CONFIG_SPACE_9,
	PondTop_input_width_17_num_0,
	PondTop_input_width_17_num_1,
	clk,
	clk_en,
	config_addr_in,
	config_data_in,
	config_en,
	config_read,
	config_write,
	flush,
	rst_n,
	tile_en,
	PondTop_output_width_17_num_0,
	PondTop_output_width_17_num_1,
	PondTop_output_width_1_num_0,
	PondTop_output_width_1_num_1,
	config_data_out
);
	input wire [31:0] CONFIG_SPACE_0;
	input wire [31:0] CONFIG_SPACE_1;
	input wire [31:0] CONFIG_SPACE_10;
	input wire [31:0] CONFIG_SPACE_11;
	input wire [31:0] CONFIG_SPACE_12;
	input wire [31:0] CONFIG_SPACE_13;
	input wire [31:0] CONFIG_SPACE_14;
	input wire [31:0] CONFIG_SPACE_15;
	input wire [29:0] CONFIG_SPACE_16;
	input wire [31:0] CONFIG_SPACE_2;
	input wire [31:0] CONFIG_SPACE_3;
	input wire [31:0] CONFIG_SPACE_4;
	input wire [31:0] CONFIG_SPACE_5;
	input wire [31:0] CONFIG_SPACE_6;
	input wire [31:0] CONFIG_SPACE_7;
	input wire [31:0] CONFIG_SPACE_8;
	input wire [31:0] CONFIG_SPACE_9;
	input wire [16:0] PondTop_input_width_17_num_0;
	input wire [16:0] PondTop_input_width_17_num_1;
	input wire clk;
	input wire clk_en;
	input wire [7:0] config_addr_in;
	input wire [31:0] config_data_in;
	input wire config_en;
	input wire config_read;
	input wire config_write;
	input wire flush;
	input wire rst_n;
	input wire tile_en;
	output reg [16:0] PondTop_output_width_17_num_0;
	output reg [16:0] PondTop_output_width_17_num_1;
	output reg PondTop_output_width_1_num_0;
	output reg PondTop_output_width_1_num_1;
	output wire [31:0] config_data_out;
	wire [541:0] CONFIG_SPACE;
	wire [15:0] config_data_in_shrt;
	wire [15:0] config_data_out_shrt;
	wire [4:0] config_seq_addr_out;
	wire config_seq_clk_en;
	reg [15:0] config_seq_rd_data_stg;
	wire config_seq_ren_out;
	wire config_seq_wen_out;
	wire [15:0] config_seq_wr_data;
	wire gclk;
	wire mem_ctrl_strg_ub_thin_PondTop_flat_clk;
	wire [16:0] mem_ctrl_strg_ub_thin_PondTop_flat_data_out_f_0;
	wire [16:0] mem_ctrl_strg_ub_thin_PondTop_flat_data_out_f_1;
	reg [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_data_from_strg_lifted;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_data_to_strg_lifted;
	wire [4:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_starting_addr;
	wire [4:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_starting_addr2;
	wire [4:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides2_0;
	wire [4:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides2_1;
	wire [4:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides_0;
	wire [4:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides_1;
	wire [4:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides_2;
	wire [4:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides_3;
	wire [2:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_dimensionality;
	wire [1:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_dimensionality2;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges2_0;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges2_1;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges_0;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges_1;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges_2;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges_3;
	wire mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_enable;
	wire mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_enable2;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_starting_addr;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_starting_addr2;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides2_0;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides2_1;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_0;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_1;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_2;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_3;
	wire [4:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_rd_addr_out_lifted;
	wire [4:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_starting_addr;
	wire [4:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_starting_addr2;
	wire [4:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides2_0;
	wire [4:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides2_1;
	wire [4:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides_0;
	wire [4:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides_1;
	wire [4:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides_2;
	wire [4:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides_3;
	wire [2:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_dimensionality;
	wire [1:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_dimensionality2;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges2_0;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges2_1;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges_0;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges_1;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges_2;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges_3;
	wire mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_enable;
	wire mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_enable2;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_starting_addr;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_starting_addr2;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides2_0;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides2_1;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_0;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_1;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_2;
	wire [15:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_3;
	wire mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_ren_to_strg_lifted;
	wire [4:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_tmp0_rdaddr_lifted;
	wire mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_tmp0_rden_lifted;
	wire mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_wen_to_strg_lifted;
	wire [4:0] mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_wr_addr_out_lifted;
	wire mem_ctrl_strg_ub_thin_PondTop_flat_valid_out_f_b_0;
	wire mem_ctrl_strg_ub_thin_PondTop_flat_valid_out_f_b_1;
	wire memory_0_clk_en;
	reg [15:0] memory_0_data_in_p0;
	wire [15:0] memory_0_data_out_p0;
	wire [15:0] memory_0_data_out_p1;
	reg [4:0] memory_0_read_addr_p0;
	reg [4:0] memory_0_read_addr_p1;
	reg memory_0_read_enable_p0;
	reg memory_0_read_enable_p1;
	reg [4:0] memory_0_write_addr_p0;
	reg memory_0_write_enable_p0;
	wire mode;
	assign mode = 1'h0;
	assign gclk = clk & tile_en;
	assign mem_ctrl_strg_ub_thin_PondTop_flat_clk = gclk;
	always @(*) begin
		PondTop_output_width_17_num_0 = 17'h00000;
		if (1'h0 == mode)
			PondTop_output_width_17_num_0 = mem_ctrl_strg_ub_thin_PondTop_flat_data_out_f_0;
		else
			PondTop_output_width_17_num_0 = 17'h00000;
	end
	always @(*) begin
		PondTop_output_width_17_num_1 = 17'h00000;
		if (1'h0 == mode)
			PondTop_output_width_17_num_1 = mem_ctrl_strg_ub_thin_PondTop_flat_data_out_f_1;
		else
			PondTop_output_width_17_num_1 = 17'h00000;
	end
	always @(*) begin
		PondTop_output_width_1_num_0 = 1'h0;
		if (1'h0 == mode)
			PondTop_output_width_1_num_0 = mem_ctrl_strg_ub_thin_PondTop_flat_valid_out_f_b_0;
		else
			PondTop_output_width_1_num_0 = 1'h0;
	end
	always @(*) begin
		PondTop_output_width_1_num_1 = 1'h0;
		if (1'h0 == mode)
			PondTop_output_width_1_num_1 = mem_ctrl_strg_ub_thin_PondTop_flat_valid_out_f_b_1;
		else
			PondTop_output_width_1_num_1 = 1'h0;
	end
	always @(*) begin
		memory_0_data_in_p0 = 16'h0000;
		memory_0_write_addr_p0 = 5'h00;
		memory_0_write_enable_p0 = 1'h0;
		memory_0_read_addr_p0 = 5'h00;
		memory_0_read_enable_p0 = 1'h0;
		if (|config_en) begin
			memory_0_data_in_p0 = config_seq_wr_data;
			memory_0_write_addr_p0 = config_seq_addr_out;
			memory_0_write_enable_p0 = config_seq_wen_out;
			memory_0_read_addr_p0 = config_seq_addr_out;
			memory_0_read_enable_p0 = config_seq_ren_out;
		end
		else if (1'h0 == mode) begin
			memory_0_data_in_p0 = mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_data_to_strg_lifted;
			memory_0_write_addr_p0 = mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_wr_addr_out_lifted;
			memory_0_write_enable_p0 = mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_wen_to_strg_lifted;
			memory_0_read_addr_p0 = mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_tmp0_rdaddr_lifted;
			memory_0_read_enable_p0 = mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_tmp0_rden_lifted;
		end
	end
	always @(*) config_seq_rd_data_stg = memory_0_data_out_p0;
	always @(*) begin
		memory_0_read_addr_p1 = 5'h00;
		memory_0_read_enable_p1 = 1'h0;
		if (1'h0 == mode) begin
			memory_0_read_addr_p1 = mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_rd_addr_out_lifted;
			memory_0_read_enable_p1 = mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_ren_to_strg_lifted;
		end
	end
	always @(*) mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_data_from_strg_lifted = memory_0_data_out_p1;
	assign config_data_in_shrt = config_data_in[15:0];
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	assign config_data_out[0+:32] = sv2v_cast_32(config_data_out_shrt[0+:16]);
	assign config_seq_clk_en = clk_en | |config_en;
	assign memory_0_clk_en = clk_en | |config_en;
	assign {mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_starting_addr, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_starting_addr2, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides2_0, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides2_1, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides_0, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides_1, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides_2, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides_3, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_dimensionality, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_dimensionality2, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges2_0, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges2_1, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges_0, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges_1, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges_2, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges_3, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_enable, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_enable2, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_starting_addr, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_starting_addr2, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides2_0, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides2_1, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_0, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_1, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_2, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_3, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_starting_addr, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_starting_addr2, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides2_0, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides2_1, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides_0, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides_1, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides_2, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides_3, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_dimensionality, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_dimensionality2, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges2_0, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges2_1, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges_0, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges_1, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges_2, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges_3, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_enable, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_enable2, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_starting_addr, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_starting_addr2, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides2_0, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides2_1, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_0, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_1, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_2, mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_3} = CONFIG_SPACE[541:0];
	assign CONFIG_SPACE[31:0] = CONFIG_SPACE_0;
	assign CONFIG_SPACE[63:32] = CONFIG_SPACE_1;
	assign CONFIG_SPACE[95:64] = CONFIG_SPACE_2;
	assign CONFIG_SPACE[127:96] = CONFIG_SPACE_3;
	assign CONFIG_SPACE[159:128] = CONFIG_SPACE_4;
	assign CONFIG_SPACE[191:160] = CONFIG_SPACE_5;
	assign CONFIG_SPACE[223:192] = CONFIG_SPACE_6;
	assign CONFIG_SPACE[255:224] = CONFIG_SPACE_7;
	assign CONFIG_SPACE[287:256] = CONFIG_SPACE_8;
	assign CONFIG_SPACE[319:288] = CONFIG_SPACE_9;
	assign CONFIG_SPACE[351:320] = CONFIG_SPACE_10;
	assign CONFIG_SPACE[383:352] = CONFIG_SPACE_11;
	assign CONFIG_SPACE[415:384] = CONFIG_SPACE_12;
	assign CONFIG_SPACE[447:416] = CONFIG_SPACE_13;
	assign CONFIG_SPACE[479:448] = CONFIG_SPACE_14;
	assign CONFIG_SPACE[511:480] = CONFIG_SPACE_15;
	assign CONFIG_SPACE[541:512] = CONFIG_SPACE_16;
	strg_ub_thin_PondTop_flat mem_ctrl_strg_ub_thin_PondTop_flat(
		.clk(mem_ctrl_strg_ub_thin_PondTop_flat_clk),
		.clk_en(clk_en),
		.data_in_f_0(PondTop_input_width_17_num_0),
		.data_in_f_1(PondTop_input_width_17_num_1),
		.flush(flush),
		.rst_n(rst_n),
		.strg_ub_thin_PondTop_inst_data_from_strg_lifted(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_data_from_strg_lifted),
		.strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_starting_addr(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_starting_addr),
		.strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_starting_addr2(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_starting_addr2),
		.strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides2_0(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides2_0),
		.strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides2_1(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides2_1),
		.strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides_0(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides_0),
		.strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides_1(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides_1),
		.strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides_2(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides_2),
		.strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides_3(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides_3),
		.strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_dimensionality(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_dimensionality),
		.strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_dimensionality2(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_dimensionality2),
		.strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges2_0(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges2_0),
		.strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges2_1(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges2_1),
		.strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges_0(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges_0),
		.strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges_1(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges_1),
		.strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges_2(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges_2),
		.strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges_3(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges_3),
		.strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_enable(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_enable),
		.strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_enable2(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_enable2),
		.strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_starting_addr),
		.strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_starting_addr2(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_starting_addr2),
		.strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides2_0(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides2_0),
		.strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides2_1(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides2_1),
		.strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_0(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_0),
		.strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_1(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_1),
		.strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_2(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_2),
		.strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_3(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_3),
		.strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_starting_addr(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_starting_addr),
		.strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_starting_addr2(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_starting_addr2),
		.strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides2_0(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides2_0),
		.strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides2_1(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides2_1),
		.strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides_0(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides_0),
		.strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides_1(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides_1),
		.strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides_2(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides_2),
		.strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides_3(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides_3),
		.strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_dimensionality(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_dimensionality),
		.strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_dimensionality2(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_dimensionality2),
		.strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges2_0(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges2_0),
		.strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges2_1(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges2_1),
		.strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges_0(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges_0),
		.strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges_1(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges_1),
		.strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges_2(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges_2),
		.strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges_3(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges_3),
		.strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_enable(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_enable),
		.strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_enable2(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_enable2),
		.strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_starting_addr),
		.strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_starting_addr2(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_starting_addr2),
		.strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides2_0(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides2_0),
		.strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides2_1(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides2_1),
		.strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_0(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_0),
		.strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_1(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_1),
		.strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_2(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_2),
		.strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_3(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_3),
		.data_out_f_0(mem_ctrl_strg_ub_thin_PondTop_flat_data_out_f_0),
		.data_out_f_1(mem_ctrl_strg_ub_thin_PondTop_flat_data_out_f_1),
		.strg_ub_thin_PondTop_inst_data_to_strg_lifted(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_data_to_strg_lifted),
		.strg_ub_thin_PondTop_inst_rd_addr_out_lifted(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_rd_addr_out_lifted),
		.strg_ub_thin_PondTop_inst_ren_to_strg_lifted(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_ren_to_strg_lifted),
		.strg_ub_thin_PondTop_inst_tmp0_rdaddr_lifted(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_tmp0_rdaddr_lifted),
		.strg_ub_thin_PondTop_inst_tmp0_rden_lifted(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_tmp0_rden_lifted),
		.strg_ub_thin_PondTop_inst_wen_to_strg_lifted(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_wen_to_strg_lifted),
		.strg_ub_thin_PondTop_inst_wr_addr_out_lifted(mem_ctrl_strg_ub_thin_PondTop_flat_strg_ub_thin_PondTop_inst_wr_addr_out_lifted),
		.valid_out_f_b_0(mem_ctrl_strg_ub_thin_PondTop_flat_valid_out_f_b_0),
		.valid_out_f_b_1(mem_ctrl_strg_ub_thin_PondTop_flat_valid_out_f_b_1)
	);
	sram_dp__0 memory_0(
		.clk(gclk),
		.clk_en(memory_0_clk_en),
		.data_in_p0(memory_0_data_in_p0),
		.flush(flush),
		.read_addr_p0(memory_0_read_addr_p0),
		.read_addr_p1(memory_0_read_addr_p1),
		.read_enable_p0(memory_0_read_enable_p0),
		.read_enable_p1(memory_0_read_enable_p1),
		.write_addr_p0(memory_0_write_addr_p0),
		.write_enable_p0(memory_0_write_enable_p0),
		.data_out_p0(memory_0_data_out_p0),
		.data_out_p1(memory_0_data_out_p1)
	);
	storage_config_seq_1_16_16 config_seq(
		.clk(gclk),
		.clk_en(config_seq_clk_en),
		.config_addr_in(config_addr_in),
		.config_data_in(config_data_in_shrt),
		.config_en(config_en),
		.config_rd(config_read),
		.config_wr(config_write),
		.flush(flush),
		.rd_data_stg(config_seq_rd_data_stg),
		.rst_n(rst_n),
		.addr_out(config_seq_addr_out),
		.rd_data_out(config_data_out_shrt),
		.ren_out(config_seq_ren_out),
		.wen_out(config_seq_wen_out),
		.wr_data(config_seq_wr_data)
	);
endmodule
module PondTop_W (
	CONFIG_SPACE_0,
	CONFIG_SPACE_1,
	CONFIG_SPACE_10,
	CONFIG_SPACE_11,
	CONFIG_SPACE_12,
	CONFIG_SPACE_13,
	CONFIG_SPACE_14,
	CONFIG_SPACE_15,
	CONFIG_SPACE_16,
	CONFIG_SPACE_2,
	CONFIG_SPACE_3,
	CONFIG_SPACE_4,
	CONFIG_SPACE_5,
	CONFIG_SPACE_6,
	CONFIG_SPACE_7,
	CONFIG_SPACE_8,
	CONFIG_SPACE_9,
	PondTop_input_width_17_num_0,
	PondTop_input_width_17_num_1,
	clk,
	clk_en,
	config_addr_in,
	config_data_in,
	config_en,
	config_read,
	config_write,
	flush,
	rst_n,
	tile_en,
	PondTop_output_width_17_num_0,
	PondTop_output_width_17_num_1,
	PondTop_output_width_1_num_0,
	PondTop_output_width_1_num_1,
	config_data_out
);
	input wire [31:0] CONFIG_SPACE_0;
	input wire [31:0] CONFIG_SPACE_1;
	input wire [31:0] CONFIG_SPACE_10;
	input wire [31:0] CONFIG_SPACE_11;
	input wire [31:0] CONFIG_SPACE_12;
	input wire [31:0] CONFIG_SPACE_13;
	input wire [31:0] CONFIG_SPACE_14;
	input wire [31:0] CONFIG_SPACE_15;
	input wire [29:0] CONFIG_SPACE_16;
	input wire [31:0] CONFIG_SPACE_2;
	input wire [31:0] CONFIG_SPACE_3;
	input wire [31:0] CONFIG_SPACE_4;
	input wire [31:0] CONFIG_SPACE_5;
	input wire [31:0] CONFIG_SPACE_6;
	input wire [31:0] CONFIG_SPACE_7;
	input wire [31:0] CONFIG_SPACE_8;
	input wire [31:0] CONFIG_SPACE_9;
	input wire [16:0] PondTop_input_width_17_num_0;
	input wire [16:0] PondTop_input_width_17_num_1;
	input wire clk;
	input wire clk_en;
	input wire [7:0] config_addr_in;
	input wire [31:0] config_data_in;
	input wire config_en;
	input wire config_read;
	input wire config_write;
	input wire flush;
	input wire rst_n;
	input wire tile_en;
	output wire [16:0] PondTop_output_width_17_num_0;
	output wire [16:0] PondTop_output_width_17_num_1;
	output wire PondTop_output_width_1_num_0;
	output wire PondTop_output_width_1_num_1;
	output wire [31:0] config_data_out;
	PondTop PondTop(
		.CONFIG_SPACE_0(CONFIG_SPACE_0),
		.CONFIG_SPACE_1(CONFIG_SPACE_1),
		.CONFIG_SPACE_10(CONFIG_SPACE_10),
		.CONFIG_SPACE_11(CONFIG_SPACE_11),
		.CONFIG_SPACE_12(CONFIG_SPACE_12),
		.CONFIG_SPACE_13(CONFIG_SPACE_13),
		.CONFIG_SPACE_14(CONFIG_SPACE_14),
		.CONFIG_SPACE_15(CONFIG_SPACE_15),
		.CONFIG_SPACE_16(CONFIG_SPACE_16),
		.CONFIG_SPACE_2(CONFIG_SPACE_2),
		.CONFIG_SPACE_3(CONFIG_SPACE_3),
		.CONFIG_SPACE_4(CONFIG_SPACE_4),
		.CONFIG_SPACE_5(CONFIG_SPACE_5),
		.CONFIG_SPACE_6(CONFIG_SPACE_6),
		.CONFIG_SPACE_7(CONFIG_SPACE_7),
		.CONFIG_SPACE_8(CONFIG_SPACE_8),
		.CONFIG_SPACE_9(CONFIG_SPACE_9),
		.PondTop_input_width_17_num_0(PondTop_input_width_17_num_0),
		.PondTop_input_width_17_num_1(PondTop_input_width_17_num_1),
		.clk(clk),
		.clk_en(clk_en),
		.config_addr_in(config_addr_in),
		.config_data_in(config_data_in),
		.config_en(config_en),
		.config_read(config_read),
		.config_write(config_write),
		.flush(flush),
		.rst_n(rst_n),
		.tile_en(tile_en),
		.PondTop_output_width_17_num_0(PondTop_output_width_17_num_0),
		.PondTop_output_width_17_num_1(PondTop_output_width_17_num_1),
		.PondTop_output_width_1_num_0(PondTop_output_width_1_num_0),
		.PondTop_output_width_1_num_1(PondTop_output_width_1_num_1),
		.config_data_out(config_data_out)
	);
endmodule
module addr_gen_4_16_dual_config_2 (
	clk,
	clk_en,
	flush,
	mux_sel,
	mux_sel_msb_init,
	restart,
	rst_n,
	starting_addr,
	starting_addr2,
	step,
	strides,
	strides2,
	addr_out,
	starting_addr_comp
);
	input wire clk;
	input wire clk_en;
	input wire flush;
	input wire [2:0] mux_sel;
	input wire mux_sel_msb_init;
	input wire restart;
	input wire rst_n;
	input wire [15:0] starting_addr;
	input wire [15:0] starting_addr2;
	input wire step;
	input wire [63:0] strides;
	input wire [31:0] strides2;
	output wire [15:0] addr_out;
	output wire starting_addr_comp;
	wire [15:0] calc_addr;
	wire [15:0] cur_stride;
	reg [15:0] current_addr;
	wire [15:0] flush_addr;
	wire [1:0] mux_sel_iter1;
	wire mux_sel_iter2;
	wire mux_sel_msb;
	wire [15:0] restart_addr;
	wire [15:0] strt_addr;
	assign starting_addr_comp = starting_addr2 < starting_addr;
	assign mux_sel_iter1 = mux_sel[1:0];
	assign mux_sel_iter2 = mux_sel[0];
	assign mux_sel_msb = mux_sel[2];
	assign flush_addr = (mux_sel_msb_init ? starting_addr2 : starting_addr);
	assign strt_addr = (mux_sel_msb ? starting_addr2 : starting_addr);
	assign restart_addr = (~mux_sel_msb ? starting_addr2 : starting_addr);
	assign cur_stride = (mux_sel_msb ? strides2[mux_sel_iter2 * 16+:16] : strides[mux_sel_iter1 * 16+:16]);
	assign addr_out = calc_addr;
	assign calc_addr = current_addr;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			current_addr <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				current_addr <= flush_addr;
			else if (step) begin
				if (restart)
					current_addr <= restart_addr;
				else
					current_addr <= current_addr + cur_stride;
			end
		end
endmodule
module addr_gen_4_5_dual_config_2 (
	clk,
	clk_en,
	flush,
	mux_sel,
	mux_sel_msb_init,
	restart,
	rst_n,
	starting_addr,
	starting_addr2,
	step,
	strides,
	strides2,
	addr_out,
	starting_addr_comp
);
	input wire clk;
	input wire clk_en;
	input wire flush;
	input wire [2:0] mux_sel;
	input wire mux_sel_msb_init;
	input wire restart;
	input wire rst_n;
	input wire [4:0] starting_addr;
	input wire [4:0] starting_addr2;
	input wire step;
	input wire [19:0] strides;
	input wire [9:0] strides2;
	output wire [4:0] addr_out;
	output wire starting_addr_comp;
	wire [4:0] calc_addr;
	wire [4:0] cur_stride;
	reg [4:0] current_addr;
	wire [4:0] flush_addr;
	wire [1:0] mux_sel_iter1;
	wire mux_sel_iter2;
	wire mux_sel_msb;
	wire [4:0] restart_addr;
	wire [4:0] strt_addr;
	assign starting_addr_comp = starting_addr2 < starting_addr;
	assign mux_sel_iter1 = mux_sel[1:0];
	assign mux_sel_iter2 = mux_sel[0];
	assign mux_sel_msb = mux_sel[2];
	assign flush_addr = (mux_sel_msb_init ? starting_addr2 : starting_addr);
	assign strt_addr = (mux_sel_msb ? starting_addr2 : starting_addr);
	assign restart_addr = (~mux_sel_msb ? starting_addr2 : starting_addr);
	assign cur_stride = (mux_sel_msb ? strides2[mux_sel_iter2 * 5+:5] : strides[mux_sel_iter1 * 5+:5]);
	assign addr_out = calc_addr;
	assign calc_addr = current_addr;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			current_addr <= 5'h00;
		else if (clk_en) begin
			if (flush)
				current_addr <= flush_addr;
			else if (step) begin
				if (restart)
					current_addr <= restart_addr;
				else
					current_addr <= current_addr + cur_stride;
			end
		end
endmodule
module for_loop_dual_config_4_2_16 (
	clk,
	clk_en,
	dimensionality,
	dimensionality2,
	flush,
	mux_sel_msb_init,
	ranges,
	ranges2,
	rst_n,
	step,
	mux_sel_out,
	restart
);
	parameter CONFIG_WIDTH = 5'h10;
	parameter ITERATOR_SUPPORT = 3'h4;
	parameter ITERATOR_SUPPORT2 = 2'h2;
	input wire clk;
	input wire clk_en;
	input wire [2:0] dimensionality;
	input wire [1:0] dimensionality2;
	input wire flush;
	input wire mux_sel_msb_init;
	input wire [63:0] ranges;
	input wire [31:0] ranges2;
	input wire rst_n;
	input wire step;
	output wire [2:0] mux_sel_out;
	output wire restart;
	reg [3:0] clear;
	wire [2:0] cur_dimensionality;
	wire [15:0] cur_range;
	reg [63:0] dim_counter;
	reg done;
	reg [3:0] inc;
	wire [15:0] inced_cnt;
	reg [3:0] max_value;
	wire maxed_value;
	reg [1:0] mux_sel;
	wire [1:0] mux_sel_iter1;
	wire mux_sel_iter2;
	wire mux_sel_msb;
	reg mux_sel_msb_r;
	assign mux_sel_msb = mux_sel_msb_r;
	function automatic [2:0] sv2v_cast_3;
		input reg [2:0] inp;
		sv2v_cast_3 = inp;
	endfunction
	assign cur_dimensionality = (mux_sel_msb ? sv2v_cast_3(dimensionality2) : dimensionality);
	assign mux_sel_iter1 = mux_sel[1:0];
	assign mux_sel_iter2 = mux_sel[0];
	assign mux_sel_out = {mux_sel_msb, mux_sel};
	assign inced_cnt = dim_counter[mux_sel * 16+:16] + 16'h0001;
	assign cur_range = (mux_sel_msb ? ranges2[mux_sel_iter2 * 16+:16] : ranges[mux_sel_iter1 * 16+:16]);
	assign maxed_value = (dim_counter[mux_sel * 16+:16] == cur_range) & inc[mux_sel];
	always @(*) begin
		mux_sel = 2'h0;
		done = 1'h0;
		if (~done) begin
			if (~max_value[0] & (cur_dimensionality > 3'h0)) begin
				mux_sel = 2'h0;
				done = 1'h1;
			end
		end
		if (~done) begin
			if (~max_value[1] & (cur_dimensionality > 3'h1)) begin
				mux_sel = 2'h1;
				done = 1'h1;
			end
		end
		if (~done) begin
			if (~max_value[2] & (cur_dimensionality > 3'h2)) begin
				mux_sel = 2'h2;
				done = 1'h1;
			end
		end
		if (~done) begin
			if (~max_value[3] & (cur_dimensionality > 3'h3)) begin
				mux_sel = 2'h3;
				done = 1'h1;
			end
		end
	end
	always @(*) begin
		clear[0] = 1'h0;
		if (((mux_sel > 2'h0) | ~done) & step)
			clear[0] = 1'h1;
	end
	always @(*) begin
		inc[0] = 1'h0;
		if ((1'd1 & step) & (cur_dimensionality > 3'h0))
			inc[0] = 1'h1;
		else if (((mux_sel == 2'h0) & step) & (cur_dimensionality > 3'h0))
			inc[0] = 1'h1;
	end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			dim_counter[0+:16] <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				dim_counter[0+:16] <= 16'h0000;
			else if (clear[0])
				dim_counter[0+:16] <= 16'h0000;
			else if (inc[0])
				dim_counter[0+:16] <= inced_cnt;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			max_value[0] <= 1'h0;
		else if (clk_en) begin
			if (flush)
				max_value[0] <= 1'h0;
			else if (clear[0])
				max_value[0] <= 1'h0;
			else if (inc[0])
				max_value[0] <= maxed_value;
		end
	always @(*) begin
		clear[1] = 1'h0;
		if (((mux_sel > 2'h1) | ~done) & step)
			clear[1] = 1'h1;
	end
	always @(*) begin
		inc[1] = 1'h0;
		if ((1'd0 & step) & (cur_dimensionality > 3'h1))
			inc[1] = 1'h1;
		else if (((mux_sel == 2'h1) & step) & (cur_dimensionality > 3'h1))
			inc[1] = 1'h1;
	end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			dim_counter[16+:16] <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				dim_counter[16+:16] <= 16'h0000;
			else if (clear[1])
				dim_counter[16+:16] <= 16'h0000;
			else if (inc[1])
				dim_counter[16+:16] <= inced_cnt;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			max_value[1] <= 1'h0;
		else if (clk_en) begin
			if (flush)
				max_value[1] <= 1'h0;
			else if (clear[1])
				max_value[1] <= 1'h0;
			else if (inc[1])
				max_value[1] <= maxed_value;
		end
	always @(*) begin
		clear[2] = 1'h0;
		if (((mux_sel > 2'h2) | ~done) & step)
			clear[2] = 1'h1;
	end
	always @(*) begin
		inc[2] = 1'h0;
		if ((1'd0 & step) & (cur_dimensionality > 3'h2))
			inc[2] = 1'h1;
		else if (((mux_sel == 2'h2) & step) & (cur_dimensionality > 3'h2))
			inc[2] = 1'h1;
	end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			dim_counter[32+:16] <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				dim_counter[32+:16] <= 16'h0000;
			else if (clear[2])
				dim_counter[32+:16] <= 16'h0000;
			else if (inc[2])
				dim_counter[32+:16] <= inced_cnt;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			max_value[2] <= 1'h0;
		else if (clk_en) begin
			if (flush)
				max_value[2] <= 1'h0;
			else if (clear[2])
				max_value[2] <= 1'h0;
			else if (inc[2])
				max_value[2] <= maxed_value;
		end
	always @(*) begin
		clear[3] = 1'h0;
		if (((mux_sel > 2'h3) | ~done) & step)
			clear[3] = 1'h1;
	end
	always @(*) begin
		inc[3] = 1'h0;
		if ((1'd0 & step) & (cur_dimensionality > 3'h3))
			inc[3] = 1'h1;
		else if (((mux_sel == 2'h3) & step) & (cur_dimensionality > 3'h3))
			inc[3] = 1'h1;
	end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			dim_counter[48+:16] <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				dim_counter[48+:16] <= 16'h0000;
			else if (clear[3])
				dim_counter[48+:16] <= 16'h0000;
			else if (inc[3])
				dim_counter[48+:16] <= inced_cnt;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			max_value[3] <= 1'h0;
		else if (clk_en) begin
			if (flush)
				max_value[3] <= 1'h0;
			else if (clear[3])
				max_value[3] <= 1'h0;
			else if (inc[3])
				max_value[3] <= maxed_value;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			mux_sel_msb_r <= 1'h0;
		else if (clk_en) begin
			if (flush)
				mux_sel_msb_r <= mux_sel_msb_init;
			else if (restart)
				mux_sel_msb_r <= ~mux_sel_msb_r;
		end
	assign restart = step & ~done;
endmodule
module sched_gen_4_16_dual_config_2 (
	clk,
	clk_en,
	cycle_count,
	enable,
	enable2,
	finished,
	flush,
	mux_sel,
	rst_n,
	sched_addr_gen_starting_addr,
	sched_addr_gen_starting_addr2,
	sched_addr_gen_strides2_0,
	sched_addr_gen_strides2_1,
	sched_addr_gen_strides_0,
	sched_addr_gen_strides_1,
	sched_addr_gen_strides_2,
	sched_addr_gen_strides_3,
	mux_sel_msb_init,
	valid_output
);
	input wire clk;
	input wire clk_en;
	input wire [15:0] cycle_count;
	input wire enable;
	input wire enable2;
	input wire finished;
	input wire flush;
	input wire [2:0] mux_sel;
	input wire rst_n;
	input wire [15:0] sched_addr_gen_starting_addr;
	input wire [15:0] sched_addr_gen_starting_addr2;
	input wire [15:0] sched_addr_gen_strides2_0;
	input wire [15:0] sched_addr_gen_strides2_1;
	input wire [15:0] sched_addr_gen_strides_0;
	input wire [15:0] sched_addr_gen_strides_1;
	input wire [15:0] sched_addr_gen_strides_2;
	input wire [15:0] sched_addr_gen_strides_3;
	output wire mux_sel_msb_init;
	output reg valid_output;
	wire [15:0] addr_out;
	wire cur_enable;
	wire cur_valid_gate;
	reg mux_sel_msb_init_w;
	wire sched_addr_gen_starting_addr_comp;
	wire [63:0] sched_addr_gen_strides;
	wire [31:0] sched_addr_gen_strides2;
	wire [1:0] valid_gate;
	reg [1:0] valid_gate_inv;
	reg valid_out;
	assign cur_valid_gate = valid_gate[mux_sel[2]];
	assign valid_gate = ~valid_gate_inv;
	assign cur_enable = (mux_sel[2] ? enable2 : enable);
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			valid_gate_inv <= 2'h0;
		else if (clk_en) begin
			if (flush)
				valid_gate_inv <= 2'h0;
			else if (finished)
				valid_gate_inv[mux_sel[2]] <= 1'h1;
		end
	always @(*)
		if (enable & enable2)
			mux_sel_msb_init_w = sched_addr_gen_starting_addr_comp;
		else if (enable & ~enable2)
			mux_sel_msb_init_w = 1'h0;
		else if (~enable & enable2)
			mux_sel_msb_init_w = 1'h1;
		else
			mux_sel_msb_init_w = 1'h0;
	assign mux_sel_msb_init = mux_sel_msb_init_w;
	always @(*) valid_out = ((cycle_count == addr_out) & cur_valid_gate) & cur_enable;
	always @(*) valid_output = valid_out;
	assign sched_addr_gen_strides2[0+:16] = sched_addr_gen_strides2_0;
	assign sched_addr_gen_strides2[16+:16] = sched_addr_gen_strides2_1;
	assign sched_addr_gen_strides[0+:16] = sched_addr_gen_strides_0;
	assign sched_addr_gen_strides[16+:16] = sched_addr_gen_strides_1;
	assign sched_addr_gen_strides[32+:16] = sched_addr_gen_strides_2;
	assign sched_addr_gen_strides[48+:16] = sched_addr_gen_strides_3;
	addr_gen_4_16_dual_config_2 sched_addr_gen(
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.mux_sel(mux_sel),
		.mux_sel_msb_init(mux_sel_msb_init_w),
		.restart(finished),
		.rst_n(rst_n),
		.starting_addr(sched_addr_gen_starting_addr),
		.starting_addr2(sched_addr_gen_starting_addr2),
		.step(valid_out),
		.strides(sched_addr_gen_strides),
		.strides2(sched_addr_gen_strides2),
		.addr_out(addr_out),
		.starting_addr_comp(sched_addr_gen_starting_addr_comp)
	);
endmodule
module sram_dp__0 (
	clk,
	clk_en,
	data_in_p0,
	flush,
	read_addr_p0,
	read_addr_p1,
	read_enable_p0,
	read_enable_p1,
	write_addr_p0,
	write_enable_p0,
	data_out_p0,
	data_out_p1
);
	input wire clk;
	input wire clk_en;
	input wire [15:0] data_in_p0;
	input wire flush;
	input wire [4:0] read_addr_p0;
	input wire [4:0] read_addr_p1;
	input wire read_enable_p0;
	input wire read_enable_p1;
	input wire [4:0] write_addr_p0;
	input wire write_enable_p0;
	output wire [15:0] data_out_p0;
	output reg [15:0] data_out_p1;
	reg [15:0] data_array [31:0];
	always @(posedge clk)
		if (clk_en) begin
			if (write_enable_p0 == 1'h1)
				data_array[write_addr_p0] <= data_in_p0;
		end
	assign data_out_p0 = data_array[read_addr_p0];
	always @(*) data_out_p1 = data_array[read_addr_p1];
endmodule
module storage_config_seq_1_16_16 (
	clk,
	clk_en,
	config_addr_in,
	config_data_in,
	config_en,
	config_rd,
	config_wr,
	flush,
	rd_data_stg,
	rst_n,
	addr_out,
	rd_data_out,
	ren_out,
	wen_out,
	wr_data
);
	input wire clk;
	input wire clk_en;
	input wire [7:0] config_addr_in;
	input wire [15:0] config_data_in;
	input wire config_en;
	input wire config_rd;
	input wire config_wr;
	input wire flush;
	input wire [15:0] rd_data_stg;
	input wire rst_n;
	output wire [4:0] addr_out;
	output wire [15:0] rd_data_out;
	output wire ren_out;
	output wire wen_out;
	output wire [15:0] wr_data;
	assign addr_out = config_addr_in[4:0];
	assign wr_data[0+:16] = config_data_in;
	assign rd_data_out[0+:16] = rd_data_stg[0+:16];
	assign wen_out = config_wr;
	assign ren_out = config_rd;
endmodule
module strg_ub_thin_PondTop (
	clk,
	clk_en,
	data_from_strg,
	data_in,
	flush,
	in2regfile_0_addr_gen_starting_addr,
	in2regfile_0_addr_gen_starting_addr2,
	in2regfile_0_addr_gen_strides2_0,
	in2regfile_0_addr_gen_strides2_1,
	in2regfile_0_addr_gen_strides_0,
	in2regfile_0_addr_gen_strides_1,
	in2regfile_0_addr_gen_strides_2,
	in2regfile_0_addr_gen_strides_3,
	in2regfile_0_for_loop_dimensionality,
	in2regfile_0_for_loop_dimensionality2,
	in2regfile_0_for_loop_ranges2_0,
	in2regfile_0_for_loop_ranges2_1,
	in2regfile_0_for_loop_ranges_0,
	in2regfile_0_for_loop_ranges_1,
	in2regfile_0_for_loop_ranges_2,
	in2regfile_0_for_loop_ranges_3,
	in2regfile_0_sched_gen_enable,
	in2regfile_0_sched_gen_enable2,
	in2regfile_0_sched_gen_sched_addr_gen_starting_addr,
	in2regfile_0_sched_gen_sched_addr_gen_starting_addr2,
	in2regfile_0_sched_gen_sched_addr_gen_strides2_0,
	in2regfile_0_sched_gen_sched_addr_gen_strides2_1,
	in2regfile_0_sched_gen_sched_addr_gen_strides_0,
	in2regfile_0_sched_gen_sched_addr_gen_strides_1,
	in2regfile_0_sched_gen_sched_addr_gen_strides_2,
	in2regfile_0_sched_gen_sched_addr_gen_strides_3,
	regfile2out_0_addr_gen_starting_addr,
	regfile2out_0_addr_gen_starting_addr2,
	regfile2out_0_addr_gen_strides2_0,
	regfile2out_0_addr_gen_strides2_1,
	regfile2out_0_addr_gen_strides_0,
	regfile2out_0_addr_gen_strides_1,
	regfile2out_0_addr_gen_strides_2,
	regfile2out_0_addr_gen_strides_3,
	regfile2out_0_for_loop_dimensionality,
	regfile2out_0_for_loop_dimensionality2,
	regfile2out_0_for_loop_ranges2_0,
	regfile2out_0_for_loop_ranges2_1,
	regfile2out_0_for_loop_ranges_0,
	regfile2out_0_for_loop_ranges_1,
	regfile2out_0_for_loop_ranges_2,
	regfile2out_0_for_loop_ranges_3,
	regfile2out_0_sched_gen_enable,
	regfile2out_0_sched_gen_enable2,
	regfile2out_0_sched_gen_sched_addr_gen_starting_addr,
	regfile2out_0_sched_gen_sched_addr_gen_starting_addr2,
	regfile2out_0_sched_gen_sched_addr_gen_strides2_0,
	regfile2out_0_sched_gen_sched_addr_gen_strides2_1,
	regfile2out_0_sched_gen_sched_addr_gen_strides_0,
	regfile2out_0_sched_gen_sched_addr_gen_strides_1,
	regfile2out_0_sched_gen_sched_addr_gen_strides_2,
	regfile2out_0_sched_gen_sched_addr_gen_strides_3,
	rst_n,
	data_out,
	data_to_strg,
	rd_addr_out,
	ren_to_strg,
	tmp0_rdaddr,
	tmp0_rden,
	valid_out,
	wen_to_strg,
	wr_addr_out
);
	input wire clk;
	input wire clk_en;
	input wire [15:0] data_from_strg;
	input wire [33:0] data_in;
	input wire flush;
	input wire [4:0] in2regfile_0_addr_gen_starting_addr;
	input wire [4:0] in2regfile_0_addr_gen_starting_addr2;
	input wire [4:0] in2regfile_0_addr_gen_strides2_0;
	input wire [4:0] in2regfile_0_addr_gen_strides2_1;
	input wire [4:0] in2regfile_0_addr_gen_strides_0;
	input wire [4:0] in2regfile_0_addr_gen_strides_1;
	input wire [4:0] in2regfile_0_addr_gen_strides_2;
	input wire [4:0] in2regfile_0_addr_gen_strides_3;
	input wire [2:0] in2regfile_0_for_loop_dimensionality;
	input wire [1:0] in2regfile_0_for_loop_dimensionality2;
	input wire [15:0] in2regfile_0_for_loop_ranges2_0;
	input wire [15:0] in2regfile_0_for_loop_ranges2_1;
	input wire [15:0] in2regfile_0_for_loop_ranges_0;
	input wire [15:0] in2regfile_0_for_loop_ranges_1;
	input wire [15:0] in2regfile_0_for_loop_ranges_2;
	input wire [15:0] in2regfile_0_for_loop_ranges_3;
	input wire in2regfile_0_sched_gen_enable;
	input wire in2regfile_0_sched_gen_enable2;
	input wire [15:0] in2regfile_0_sched_gen_sched_addr_gen_starting_addr;
	input wire [15:0] in2regfile_0_sched_gen_sched_addr_gen_starting_addr2;
	input wire [15:0] in2regfile_0_sched_gen_sched_addr_gen_strides2_0;
	input wire [15:0] in2regfile_0_sched_gen_sched_addr_gen_strides2_1;
	input wire [15:0] in2regfile_0_sched_gen_sched_addr_gen_strides_0;
	input wire [15:0] in2regfile_0_sched_gen_sched_addr_gen_strides_1;
	input wire [15:0] in2regfile_0_sched_gen_sched_addr_gen_strides_2;
	input wire [15:0] in2regfile_0_sched_gen_sched_addr_gen_strides_3;
	input wire [4:0] regfile2out_0_addr_gen_starting_addr;
	input wire [4:0] regfile2out_0_addr_gen_starting_addr2;
	input wire [4:0] regfile2out_0_addr_gen_strides2_0;
	input wire [4:0] regfile2out_0_addr_gen_strides2_1;
	input wire [4:0] regfile2out_0_addr_gen_strides_0;
	input wire [4:0] regfile2out_0_addr_gen_strides_1;
	input wire [4:0] regfile2out_0_addr_gen_strides_2;
	input wire [4:0] regfile2out_0_addr_gen_strides_3;
	input wire [2:0] regfile2out_0_for_loop_dimensionality;
	input wire [1:0] regfile2out_0_for_loop_dimensionality2;
	input wire [15:0] regfile2out_0_for_loop_ranges2_0;
	input wire [15:0] regfile2out_0_for_loop_ranges2_1;
	input wire [15:0] regfile2out_0_for_loop_ranges_0;
	input wire [15:0] regfile2out_0_for_loop_ranges_1;
	input wire [15:0] regfile2out_0_for_loop_ranges_2;
	input wire [15:0] regfile2out_0_for_loop_ranges_3;
	input wire regfile2out_0_sched_gen_enable;
	input wire regfile2out_0_sched_gen_enable2;
	input wire [15:0] regfile2out_0_sched_gen_sched_addr_gen_starting_addr;
	input wire [15:0] regfile2out_0_sched_gen_sched_addr_gen_starting_addr2;
	input wire [15:0] regfile2out_0_sched_gen_sched_addr_gen_strides2_0;
	input wire [15:0] regfile2out_0_sched_gen_sched_addr_gen_strides2_1;
	input wire [15:0] regfile2out_0_sched_gen_sched_addr_gen_strides_0;
	input wire [15:0] regfile2out_0_sched_gen_sched_addr_gen_strides_1;
	input wire [15:0] regfile2out_0_sched_gen_sched_addr_gen_strides_2;
	input wire [15:0] regfile2out_0_sched_gen_sched_addr_gen_strides_3;
	input wire rst_n;
	output wire [33:0] data_out;
	output wire [15:0] data_to_strg;
	output wire [4:0] rd_addr_out;
	output wire ren_to_strg;
	output wire [4:0] tmp0_rdaddr;
	output wire tmp0_rden;
	output wire [1:0] valid_out;
	output wire wen_to_strg;
	output wire [4:0] wr_addr_out;
	reg [15:0] cycle_count;
	wire [31:0] data_in_thin;
	wire [31:0] data_out_int;
	wire [31:0] data_out_int_thin;
	wire in2regfile_0_addr_gen_mux_sel_msb_init;
	wire [19:0] in2regfile_0_addr_gen_strides;
	wire [9:0] in2regfile_0_addr_gen_strides2;
	wire in2regfile_0_for_loop_mux_sel_msb_init;
	wire [2:0] in2regfile_0_for_loop_mux_sel_out;
	wire [63:0] in2regfile_0_for_loop_ranges;
	wire [31:0] in2regfile_0_for_loop_ranges2;
	wire in2regfile_0_for_loop_restart;
	wire in2regfile_0_sched_gen_mux_sel_msb_init;
	wire in2regfile_0_sched_gen_valid_output;
	wire read;
	wire [4:0] read_addr;
	wire read_mux_sel_msb;
	wire regfile2out_0_addr_gen_mux_sel_msb_init;
	wire [19:0] regfile2out_0_addr_gen_strides;
	wire [9:0] regfile2out_0_addr_gen_strides2;
	wire regfile2out_0_for_loop_mux_sel_msb_init;
	wire [2:0] regfile2out_0_for_loop_mux_sel_out;
	wire [63:0] regfile2out_0_for_loop_ranges;
	wire [31:0] regfile2out_0_for_loop_ranges2;
	wire regfile2out_0_for_loop_restart;
	wire regfile2out_0_sched_gen_mux_sel_msb_init;
	wire regfile2out_0_sched_gen_valid_output;
	wire [1:0] valid_out_int;
	wire write;
	wire [4:0] write_addr;
	wire write_mux_sel_msb;
	assign data_in_thin[0+:16] = data_in[15-:16];
	assign data_in_thin[16+:16] = data_in[32-:16];
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			cycle_count <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				cycle_count <= 16'h0000;
			else
				cycle_count <= cycle_count + 16'h0001;
		end
	assign valid_out_int[0] = read & ~read_mux_sel_msb;
	assign valid_out_int[1] = read & read_mux_sel_msb;
	assign data_out_int_thin = data_out_int;
	assign data_out[15-:16] = data_out_int_thin[0+:16];
	assign data_out[16] = 1'h0;
	assign data_out[32-:16] = data_out_int_thin[16+:16];
	assign data_out[33] = 1'h0;
	assign valid_out = valid_out_int;
	assign write = in2regfile_0_sched_gen_valid_output;
	assign in2regfile_0_for_loop_mux_sel_msb_init = in2regfile_0_sched_gen_mux_sel_msb_init;
	assign in2regfile_0_addr_gen_mux_sel_msb_init = in2regfile_0_sched_gen_mux_sel_msb_init;
	assign write_mux_sel_msb = in2regfile_0_for_loop_mux_sel_out[2];
	assign read = regfile2out_0_sched_gen_valid_output;
	assign regfile2out_0_for_loop_mux_sel_msb_init = regfile2out_0_sched_gen_mux_sel_msb_init;
	assign regfile2out_0_addr_gen_mux_sel_msb_init = regfile2out_0_sched_gen_mux_sel_msb_init;
	assign read_mux_sel_msb = regfile2out_0_for_loop_mux_sel_out[2];
	assign wen_to_strg = |write;
	assign ren_to_strg = |read;
	assign data_out_int[0+:16] = data_from_strg;
	assign data_out_int[16+:16] = data_from_strg;
	assign wr_addr_out = write_addr[4:0];
	assign data_to_strg = data_in_thin[write_mux_sel_msb * 16+:16];
	assign rd_addr_out = read_addr[4:0];
	assign tmp0_rdaddr = 5'h00;
	assign tmp0_rden = 1'h0;
	assign in2regfile_0_for_loop_ranges2[0+:16] = in2regfile_0_for_loop_ranges2_0;
	assign in2regfile_0_for_loop_ranges2[16+:16] = in2regfile_0_for_loop_ranges2_1;
	assign in2regfile_0_for_loop_ranges[0+:16] = in2regfile_0_for_loop_ranges_0;
	assign in2regfile_0_for_loop_ranges[16+:16] = in2regfile_0_for_loop_ranges_1;
	assign in2regfile_0_for_loop_ranges[32+:16] = in2regfile_0_for_loop_ranges_2;
	assign in2regfile_0_for_loop_ranges[48+:16] = in2regfile_0_for_loop_ranges_3;
	assign in2regfile_0_addr_gen_strides2[0+:5] = in2regfile_0_addr_gen_strides2_0;
	assign in2regfile_0_addr_gen_strides2[5+:5] = in2regfile_0_addr_gen_strides2_1;
	assign in2regfile_0_addr_gen_strides[0+:5] = in2regfile_0_addr_gen_strides_0;
	assign in2regfile_0_addr_gen_strides[5+:5] = in2regfile_0_addr_gen_strides_1;
	assign in2regfile_0_addr_gen_strides[10+:5] = in2regfile_0_addr_gen_strides_2;
	assign in2regfile_0_addr_gen_strides[15+:5] = in2regfile_0_addr_gen_strides_3;
	assign regfile2out_0_for_loop_ranges2[0+:16] = regfile2out_0_for_loop_ranges2_0;
	assign regfile2out_0_for_loop_ranges2[16+:16] = regfile2out_0_for_loop_ranges2_1;
	assign regfile2out_0_for_loop_ranges[0+:16] = regfile2out_0_for_loop_ranges_0;
	assign regfile2out_0_for_loop_ranges[16+:16] = regfile2out_0_for_loop_ranges_1;
	assign regfile2out_0_for_loop_ranges[32+:16] = regfile2out_0_for_loop_ranges_2;
	assign regfile2out_0_for_loop_ranges[48+:16] = regfile2out_0_for_loop_ranges_3;
	assign regfile2out_0_addr_gen_strides2[0+:5] = regfile2out_0_addr_gen_strides2_0;
	assign regfile2out_0_addr_gen_strides2[5+:5] = regfile2out_0_addr_gen_strides2_1;
	assign regfile2out_0_addr_gen_strides[0+:5] = regfile2out_0_addr_gen_strides_0;
	assign regfile2out_0_addr_gen_strides[5+:5] = regfile2out_0_addr_gen_strides_1;
	assign regfile2out_0_addr_gen_strides[10+:5] = regfile2out_0_addr_gen_strides_2;
	assign regfile2out_0_addr_gen_strides[15+:5] = regfile2out_0_addr_gen_strides_3;
	for_loop_dual_config_4_2_16 in2regfile_0_for_loop(
		.clk(clk),
		.clk_en(clk_en),
		.dimensionality(in2regfile_0_for_loop_dimensionality),
		.dimensionality2(in2regfile_0_for_loop_dimensionality2),
		.flush(flush),
		.mux_sel_msb_init(in2regfile_0_for_loop_mux_sel_msb_init),
		.ranges(in2regfile_0_for_loop_ranges),
		.ranges2(in2regfile_0_for_loop_ranges2),
		.rst_n(rst_n),
		.step(write),
		.mux_sel_out(in2regfile_0_for_loop_mux_sel_out),
		.restart(in2regfile_0_for_loop_restart)
	);
	addr_gen_4_5_dual_config_2 in2regfile_0_addr_gen(
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.mux_sel(in2regfile_0_for_loop_mux_sel_out),
		.mux_sel_msb_init(in2regfile_0_addr_gen_mux_sel_msb_init),
		.restart(in2regfile_0_for_loop_restart),
		.rst_n(rst_n),
		.starting_addr(in2regfile_0_addr_gen_starting_addr),
		.starting_addr2(in2regfile_0_addr_gen_starting_addr2),
		.step(write),
		.strides(in2regfile_0_addr_gen_strides),
		.strides2(in2regfile_0_addr_gen_strides2),
		.addr_out(write_addr)
	);
	sched_gen_4_16_dual_config_2 in2regfile_0_sched_gen(
		.clk(clk),
		.clk_en(clk_en),
		.cycle_count(cycle_count),
		.enable(in2regfile_0_sched_gen_enable),
		.enable2(in2regfile_0_sched_gen_enable2),
		.finished(in2regfile_0_for_loop_restart),
		.flush(flush),
		.mux_sel(in2regfile_0_for_loop_mux_sel_out),
		.rst_n(rst_n),
		.sched_addr_gen_starting_addr(in2regfile_0_sched_gen_sched_addr_gen_starting_addr),
		.sched_addr_gen_starting_addr2(in2regfile_0_sched_gen_sched_addr_gen_starting_addr2),
		.sched_addr_gen_strides2_0(in2regfile_0_sched_gen_sched_addr_gen_strides2_0),
		.sched_addr_gen_strides2_1(in2regfile_0_sched_gen_sched_addr_gen_strides2_1),
		.sched_addr_gen_strides_0(in2regfile_0_sched_gen_sched_addr_gen_strides_0),
		.sched_addr_gen_strides_1(in2regfile_0_sched_gen_sched_addr_gen_strides_1),
		.sched_addr_gen_strides_2(in2regfile_0_sched_gen_sched_addr_gen_strides_2),
		.sched_addr_gen_strides_3(in2regfile_0_sched_gen_sched_addr_gen_strides_3),
		.mux_sel_msb_init(in2regfile_0_sched_gen_mux_sel_msb_init),
		.valid_output(in2regfile_0_sched_gen_valid_output)
	);
	for_loop_dual_config_4_2_16 regfile2out_0_for_loop(
		.clk(clk),
		.clk_en(clk_en),
		.dimensionality(regfile2out_0_for_loop_dimensionality),
		.dimensionality2(regfile2out_0_for_loop_dimensionality2),
		.flush(flush),
		.mux_sel_msb_init(regfile2out_0_for_loop_mux_sel_msb_init),
		.ranges(regfile2out_0_for_loop_ranges),
		.ranges2(regfile2out_0_for_loop_ranges2),
		.rst_n(rst_n),
		.step(read),
		.mux_sel_out(regfile2out_0_for_loop_mux_sel_out),
		.restart(regfile2out_0_for_loop_restart)
	);
	addr_gen_4_5_dual_config_2 regfile2out_0_addr_gen(
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.mux_sel(regfile2out_0_for_loop_mux_sel_out),
		.mux_sel_msb_init(regfile2out_0_addr_gen_mux_sel_msb_init),
		.restart(regfile2out_0_for_loop_restart),
		.rst_n(rst_n),
		.starting_addr(regfile2out_0_addr_gen_starting_addr),
		.starting_addr2(regfile2out_0_addr_gen_starting_addr2),
		.step(read),
		.strides(regfile2out_0_addr_gen_strides),
		.strides2(regfile2out_0_addr_gen_strides2),
		.addr_out(read_addr)
	);
	sched_gen_4_16_dual_config_2 regfile2out_0_sched_gen(
		.clk(clk),
		.clk_en(clk_en),
		.cycle_count(cycle_count),
		.enable(regfile2out_0_sched_gen_enable),
		.enable2(regfile2out_0_sched_gen_enable2),
		.finished(regfile2out_0_for_loop_restart),
		.flush(flush),
		.mux_sel(regfile2out_0_for_loop_mux_sel_out),
		.rst_n(rst_n),
		.sched_addr_gen_starting_addr(regfile2out_0_sched_gen_sched_addr_gen_starting_addr),
		.sched_addr_gen_starting_addr2(regfile2out_0_sched_gen_sched_addr_gen_starting_addr2),
		.sched_addr_gen_strides2_0(regfile2out_0_sched_gen_sched_addr_gen_strides2_0),
		.sched_addr_gen_strides2_1(regfile2out_0_sched_gen_sched_addr_gen_strides2_1),
		.sched_addr_gen_strides_0(regfile2out_0_sched_gen_sched_addr_gen_strides_0),
		.sched_addr_gen_strides_1(regfile2out_0_sched_gen_sched_addr_gen_strides_1),
		.sched_addr_gen_strides_2(regfile2out_0_sched_gen_sched_addr_gen_strides_2),
		.sched_addr_gen_strides_3(regfile2out_0_sched_gen_sched_addr_gen_strides_3),
		.mux_sel_msb_init(regfile2out_0_sched_gen_mux_sel_msb_init),
		.valid_output(regfile2out_0_sched_gen_valid_output)
	);
endmodule
module strg_ub_thin_PondTop_flat (
	clk,
	clk_en,
	data_in_f_0,
	data_in_f_1,
	flush,
	rst_n,
	strg_ub_thin_PondTop_inst_data_from_strg_lifted,
	strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_starting_addr,
	strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_starting_addr2,
	strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides2_0,
	strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides2_1,
	strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides_0,
	strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides_1,
	strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides_2,
	strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides_3,
	strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_dimensionality,
	strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_dimensionality2,
	strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges2_0,
	strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges2_1,
	strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges_0,
	strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges_1,
	strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges_2,
	strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges_3,
	strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_enable,
	strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_enable2,
	strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_starting_addr,
	strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_starting_addr2,
	strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides2_0,
	strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides2_1,
	strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_0,
	strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_1,
	strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_2,
	strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_3,
	strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_starting_addr,
	strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_starting_addr2,
	strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides2_0,
	strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides2_1,
	strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides_0,
	strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides_1,
	strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides_2,
	strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides_3,
	strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_dimensionality,
	strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_dimensionality2,
	strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges2_0,
	strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges2_1,
	strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges_0,
	strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges_1,
	strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges_2,
	strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges_3,
	strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_enable,
	strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_enable2,
	strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_starting_addr,
	strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_starting_addr2,
	strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides2_0,
	strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides2_1,
	strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_0,
	strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_1,
	strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_2,
	strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_3,
	data_out_f_0,
	data_out_f_1,
	strg_ub_thin_PondTop_inst_data_to_strg_lifted,
	strg_ub_thin_PondTop_inst_rd_addr_out_lifted,
	strg_ub_thin_PondTop_inst_ren_to_strg_lifted,
	strg_ub_thin_PondTop_inst_tmp0_rdaddr_lifted,
	strg_ub_thin_PondTop_inst_tmp0_rden_lifted,
	strg_ub_thin_PondTop_inst_wen_to_strg_lifted,
	strg_ub_thin_PondTop_inst_wr_addr_out_lifted,
	valid_out_f_b_0,
	valid_out_f_b_1
);
	input wire clk;
	input wire clk_en;
	input wire [16:0] data_in_f_0;
	input wire [16:0] data_in_f_1;
	input wire flush;
	input wire rst_n;
	input wire [15:0] strg_ub_thin_PondTop_inst_data_from_strg_lifted;
	input wire [4:0] strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_starting_addr;
	input wire [4:0] strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_starting_addr2;
	input wire [4:0] strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides2_0;
	input wire [4:0] strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides2_1;
	input wire [4:0] strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides_0;
	input wire [4:0] strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides_1;
	input wire [4:0] strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides_2;
	input wire [4:0] strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides_3;
	input wire [2:0] strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_dimensionality;
	input wire [1:0] strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_dimensionality2;
	input wire [15:0] strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges2_0;
	input wire [15:0] strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges2_1;
	input wire [15:0] strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges_0;
	input wire [15:0] strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges_1;
	input wire [15:0] strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges_2;
	input wire [15:0] strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges_3;
	input wire strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_enable;
	input wire strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_enable2;
	input wire [15:0] strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_starting_addr;
	input wire [15:0] strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_starting_addr2;
	input wire [15:0] strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides2_0;
	input wire [15:0] strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides2_1;
	input wire [15:0] strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_0;
	input wire [15:0] strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_1;
	input wire [15:0] strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_2;
	input wire [15:0] strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_3;
	input wire [4:0] strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_starting_addr;
	input wire [4:0] strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_starting_addr2;
	input wire [4:0] strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides2_0;
	input wire [4:0] strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides2_1;
	input wire [4:0] strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides_0;
	input wire [4:0] strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides_1;
	input wire [4:0] strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides_2;
	input wire [4:0] strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides_3;
	input wire [2:0] strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_dimensionality;
	input wire [1:0] strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_dimensionality2;
	input wire [15:0] strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges2_0;
	input wire [15:0] strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges2_1;
	input wire [15:0] strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges_0;
	input wire [15:0] strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges_1;
	input wire [15:0] strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges_2;
	input wire [15:0] strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges_3;
	input wire strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_enable;
	input wire strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_enable2;
	input wire [15:0] strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_starting_addr;
	input wire [15:0] strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_starting_addr2;
	input wire [15:0] strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides2_0;
	input wire [15:0] strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides2_1;
	input wire [15:0] strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_0;
	input wire [15:0] strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_1;
	input wire [15:0] strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_2;
	input wire [15:0] strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_3;
	output wire [16:0] data_out_f_0;
	output wire [16:0] data_out_f_1;
	output wire [15:0] strg_ub_thin_PondTop_inst_data_to_strg_lifted;
	output wire [4:0] strg_ub_thin_PondTop_inst_rd_addr_out_lifted;
	output wire strg_ub_thin_PondTop_inst_ren_to_strg_lifted;
	output wire [4:0] strg_ub_thin_PondTop_inst_tmp0_rdaddr_lifted;
	output wire strg_ub_thin_PondTop_inst_tmp0_rden_lifted;
	output wire strg_ub_thin_PondTop_inst_wen_to_strg_lifted;
	output wire [4:0] strg_ub_thin_PondTop_inst_wr_addr_out_lifted;
	output wire valid_out_f_b_0;
	output wire valid_out_f_b_1;
	wire [33:0] strg_ub_thin_PondTop_inst_data_in;
	wire [33:0] strg_ub_thin_PondTop_inst_data_out;
	wire [1:0] strg_ub_thin_PondTop_inst_valid_out;
	assign strg_ub_thin_PondTop_inst_data_in[0+:17] = data_in_f_0;
	assign strg_ub_thin_PondTop_inst_data_in[17+:17] = data_in_f_1;
	assign valid_out_f_b_0 = strg_ub_thin_PondTop_inst_valid_out[0];
	assign valid_out_f_b_1 = strg_ub_thin_PondTop_inst_valid_out[1];
	assign data_out_f_0 = strg_ub_thin_PondTop_inst_data_out[0+:17];
	assign data_out_f_1 = strg_ub_thin_PondTop_inst_data_out[17+:17];
	strg_ub_thin_PondTop strg_ub_thin_PondTop_inst(
		.clk(clk),
		.clk_en(clk_en),
		.data_from_strg(strg_ub_thin_PondTop_inst_data_from_strg_lifted),
		.data_in(strg_ub_thin_PondTop_inst_data_in),
		.flush(flush),
		.in2regfile_0_addr_gen_starting_addr(strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_starting_addr),
		.in2regfile_0_addr_gen_starting_addr2(strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_starting_addr2),
		.in2regfile_0_addr_gen_strides2_0(strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides2_0),
		.in2regfile_0_addr_gen_strides2_1(strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides2_1),
		.in2regfile_0_addr_gen_strides_0(strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides_0),
		.in2regfile_0_addr_gen_strides_1(strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides_1),
		.in2regfile_0_addr_gen_strides_2(strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides_2),
		.in2regfile_0_addr_gen_strides_3(strg_ub_thin_PondTop_inst_in2regfile_0_addr_gen_strides_3),
		.in2regfile_0_for_loop_dimensionality(strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_dimensionality),
		.in2regfile_0_for_loop_dimensionality2(strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_dimensionality2),
		.in2regfile_0_for_loop_ranges2_0(strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges2_0),
		.in2regfile_0_for_loop_ranges2_1(strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges2_1),
		.in2regfile_0_for_loop_ranges_0(strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges_0),
		.in2regfile_0_for_loop_ranges_1(strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges_1),
		.in2regfile_0_for_loop_ranges_2(strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges_2),
		.in2regfile_0_for_loop_ranges_3(strg_ub_thin_PondTop_inst_in2regfile_0_for_loop_ranges_3),
		.in2regfile_0_sched_gen_enable(strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_enable),
		.in2regfile_0_sched_gen_enable2(strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_enable2),
		.in2regfile_0_sched_gen_sched_addr_gen_starting_addr(strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_starting_addr),
		.in2regfile_0_sched_gen_sched_addr_gen_starting_addr2(strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_starting_addr2),
		.in2regfile_0_sched_gen_sched_addr_gen_strides2_0(strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides2_0),
		.in2regfile_0_sched_gen_sched_addr_gen_strides2_1(strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides2_1),
		.in2regfile_0_sched_gen_sched_addr_gen_strides_0(strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_0),
		.in2regfile_0_sched_gen_sched_addr_gen_strides_1(strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_1),
		.in2regfile_0_sched_gen_sched_addr_gen_strides_2(strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_2),
		.in2regfile_0_sched_gen_sched_addr_gen_strides_3(strg_ub_thin_PondTop_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_3),
		.regfile2out_0_addr_gen_starting_addr(strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_starting_addr),
		.regfile2out_0_addr_gen_starting_addr2(strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_starting_addr2),
		.regfile2out_0_addr_gen_strides2_0(strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides2_0),
		.regfile2out_0_addr_gen_strides2_1(strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides2_1),
		.regfile2out_0_addr_gen_strides_0(strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides_0),
		.regfile2out_0_addr_gen_strides_1(strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides_1),
		.regfile2out_0_addr_gen_strides_2(strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides_2),
		.regfile2out_0_addr_gen_strides_3(strg_ub_thin_PondTop_inst_regfile2out_0_addr_gen_strides_3),
		.regfile2out_0_for_loop_dimensionality(strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_dimensionality),
		.regfile2out_0_for_loop_dimensionality2(strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_dimensionality2),
		.regfile2out_0_for_loop_ranges2_0(strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges2_0),
		.regfile2out_0_for_loop_ranges2_1(strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges2_1),
		.regfile2out_0_for_loop_ranges_0(strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges_0),
		.regfile2out_0_for_loop_ranges_1(strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges_1),
		.regfile2out_0_for_loop_ranges_2(strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges_2),
		.regfile2out_0_for_loop_ranges_3(strg_ub_thin_PondTop_inst_regfile2out_0_for_loop_ranges_3),
		.regfile2out_0_sched_gen_enable(strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_enable),
		.regfile2out_0_sched_gen_enable2(strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_enable2),
		.regfile2out_0_sched_gen_sched_addr_gen_starting_addr(strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_starting_addr),
		.regfile2out_0_sched_gen_sched_addr_gen_starting_addr2(strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_starting_addr2),
		.regfile2out_0_sched_gen_sched_addr_gen_strides2_0(strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides2_0),
		.regfile2out_0_sched_gen_sched_addr_gen_strides2_1(strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides2_1),
		.regfile2out_0_sched_gen_sched_addr_gen_strides_0(strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_0),
		.regfile2out_0_sched_gen_sched_addr_gen_strides_1(strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_1),
		.regfile2out_0_sched_gen_sched_addr_gen_strides_2(strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_2),
		.regfile2out_0_sched_gen_sched_addr_gen_strides_3(strg_ub_thin_PondTop_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_3),
		.rst_n(rst_n),
		.data_out(strg_ub_thin_PondTop_inst_data_out),
		.data_to_strg(strg_ub_thin_PondTop_inst_data_to_strg_lifted),
		.rd_addr_out(strg_ub_thin_PondTop_inst_rd_addr_out_lifted),
		.ren_to_strg(strg_ub_thin_PondTop_inst_ren_to_strg_lifted),
		.tmp0_rdaddr(strg_ub_thin_PondTop_inst_tmp0_rdaddr_lifted),
		.tmp0_rden(strg_ub_thin_PondTop_inst_tmp0_rden_lifted),
		.valid_out(strg_ub_thin_PondTop_inst_valid_out),
		.wen_to_strg(strg_ub_thin_PondTop_inst_wen_to_strg_lifted),
		.wr_addr_out(strg_ub_thin_PondTop_inst_wr_addr_out_lifted)
	);
endmodule
module PE_inner (
	CONFIG_SPACE_0,
	CONFIG_SPACE_1,
	CONFIG_SPACE_2,
	PE_input_width_17_num_0,
	PE_input_width_17_num_0_dense,
	PE_input_width_17_num_0_valid,
	PE_input_width_17_num_1,
	PE_input_width_17_num_1_dense,
	PE_input_width_17_num_1_valid,
	PE_input_width_17_num_2,
	PE_input_width_17_num_2_valid,
	PE_input_width_17_num_3,
	PE_input_width_17_num_3_valid,
	PE_input_width_1_num_0,
	PE_input_width_1_num_1,
	PE_input_width_1_num_2,
	PE_output_width_17_num_0_dense,
	PE_output_width_17_num_0_ready,
	PE_output_width_17_num_1_ready,
	PE_output_width_17_num_2_ready,
	clk,
	clk_en,
	flush,
	mode,
	rst_n,
	tile_en,
	PE_input_width_17_num_0_ready,
	PE_input_width_17_num_1_ready,
	PE_input_width_17_num_2_ready,
	PE_input_width_17_num_3_ready,
	PE_onyx_inst_onyxpeintf_O2,
	PE_onyx_inst_onyxpeintf_O3,
	PE_onyx_inst_onyxpeintf_O4,
	PE_output_width_17_num_0,
	PE_output_width_17_num_0_valid,
	PE_output_width_17_num_1,
	PE_output_width_17_num_1_valid,
	PE_output_width_17_num_2,
	PE_output_width_17_num_2_valid,
	PE_output_width_1_num_0
);
	input wire [31:0] CONFIG_SPACE_0;
	input wire [31:0] CONFIG_SPACE_1;
	input wire [21:0] CONFIG_SPACE_2;
	input wire [16:0] PE_input_width_17_num_0;
	input wire PE_input_width_17_num_0_dense;
	input wire PE_input_width_17_num_0_valid;
	input wire [16:0] PE_input_width_17_num_1;
	input wire PE_input_width_17_num_1_dense;
	input wire PE_input_width_17_num_1_valid;
	input wire [16:0] PE_input_width_17_num_2;
	input wire PE_input_width_17_num_2_valid;
	input wire [16:0] PE_input_width_17_num_3;
	input wire PE_input_width_17_num_3_valid;
	input wire PE_input_width_1_num_0;
	input wire PE_input_width_1_num_1;
	input wire PE_input_width_1_num_2;
	input wire PE_output_width_17_num_0_dense;
	input wire PE_output_width_17_num_0_ready;
	input wire PE_output_width_17_num_1_ready;
	input wire PE_output_width_17_num_2_ready;
	input wire clk;
	input wire clk_en;
	input wire flush;
	input wire [2:0] mode;
	input wire rst_n;
	input wire tile_en;
	output reg PE_input_width_17_num_0_ready;
	output reg PE_input_width_17_num_1_ready;
	output reg PE_input_width_17_num_2_ready;
	output reg PE_input_width_17_num_3_ready;
	output wire [15:0] PE_onyx_inst_onyxpeintf_O2;
	output wire [15:0] PE_onyx_inst_onyxpeintf_O3;
	output wire [15:0] PE_onyx_inst_onyxpeintf_O4;
	output reg [16:0] PE_output_width_17_num_0;
	output reg PE_output_width_17_num_0_valid;
	output reg [16:0] PE_output_width_17_num_1;
	output reg PE_output_width_17_num_1_valid;
	output reg [16:0] PE_output_width_17_num_2;
	output reg PE_output_width_17_num_2_valid;
	output reg PE_output_width_1_num_0;
	wire [85:0] CONFIG_SPACE;
	wire gclk;
	wire [16:0] input_width_17_num_0_fifo_out;
	reg input_width_17_num_0_fifo_out_ready;
	wire input_width_17_num_0_fifo_out_valid;
	wire input_width_17_num_0_input_fifo_empty;
	wire input_width_17_num_0_input_fifo_full;
	wire [16:0] input_width_17_num_1_fifo_out;
	reg input_width_17_num_1_fifo_out_ready;
	wire input_width_17_num_1_fifo_out_valid;
	wire input_width_17_num_1_input_fifo_empty;
	wire input_width_17_num_1_input_fifo_full;
	wire [16:0] input_width_17_num_2_fifo_out;
	reg input_width_17_num_2_fifo_out_ready;
	wire input_width_17_num_2_fifo_out_valid;
	wire input_width_17_num_2_input_fifo_empty;
	wire input_width_17_num_2_input_fifo_full;
	wire [16:0] input_width_17_num_3_fifo_out;
	reg input_width_17_num_3_fifo_out_ready;
	wire input_width_17_num_3_fifo_out_valid;
	wire input_width_17_num_3_input_fifo_empty;
	wire input_width_17_num_3_input_fifo_full;
	wire mem_ctrl_PE_onyx_flat_PE_onyx_inst_dense_mode;
	wire [83:0] mem_ctrl_PE_onyx_flat_PE_onyx_inst_onyxpeintf_inst;
	wire mem_ctrl_PE_onyx_flat_PE_onyx_inst_tile_en;
	wire mem_ctrl_PE_onyx_flat_clk;
	wire [16:0] mem_ctrl_PE_onyx_flat_data0_f_;
	wire mem_ctrl_PE_onyx_flat_data0_ready_f_;
	wire mem_ctrl_PE_onyx_flat_data0_valid_f_;
	wire [16:0] mem_ctrl_PE_onyx_flat_data1_f_;
	wire mem_ctrl_PE_onyx_flat_data1_ready_f_;
	wire mem_ctrl_PE_onyx_flat_data1_valid_f_;
	wire [16:0] mem_ctrl_PE_onyx_flat_res_f_;
	wire mem_ctrl_PE_onyx_flat_res_p_f_;
	wire mem_ctrl_PE_onyx_flat_res_ready_f_;
	wire mem_ctrl_PE_onyx_flat_res_valid_f_;
	wire [15:0] mem_ctrl_RepeatSignalGenerator_flat_RepeatSignalGenerator_inst_stop_lvl;
	wire mem_ctrl_RepeatSignalGenerator_flat_RepeatSignalGenerator_inst_tile_en;
	wire mem_ctrl_RepeatSignalGenerator_flat_base_data_in_ready_f_;
	wire mem_ctrl_RepeatSignalGenerator_flat_clk;
	wire [16:0] mem_ctrl_RepeatSignalGenerator_flat_repsig_data_out_f_;
	wire mem_ctrl_RepeatSignalGenerator_flat_repsig_data_out_valid_f_;
	wire mem_ctrl_Repeat_flat_Repeat_inst_root;
	wire mem_ctrl_Repeat_flat_Repeat_inst_spacc_mode;
	wire [15:0] mem_ctrl_Repeat_flat_Repeat_inst_stop_lvl;
	wire mem_ctrl_Repeat_flat_Repeat_inst_tile_en;
	wire mem_ctrl_Repeat_flat_clk;
	wire mem_ctrl_Repeat_flat_proc_data_in_ready_f_;
	wire [16:0] mem_ctrl_Repeat_flat_ref_data_out_f_;
	wire mem_ctrl_Repeat_flat_ref_data_out_valid_f_;
	wire mem_ctrl_Repeat_flat_repsig_data_in_ready_f_;
	wire mem_ctrl_crddrop_flat_clk;
	wire mem_ctrl_crddrop_flat_cmrg_coord_in_0_ready_f_;
	wire mem_ctrl_crddrop_flat_cmrg_coord_in_1_ready_f_;
	wire [16:0] mem_ctrl_crddrop_flat_cmrg_coord_out_0_f_;
	wire mem_ctrl_crddrop_flat_cmrg_coord_out_0_valid_f_;
	wire [16:0] mem_ctrl_crddrop_flat_cmrg_coord_out_1_f_;
	wire mem_ctrl_crddrop_flat_cmrg_coord_out_1_valid_f_;
	wire mem_ctrl_crddrop_flat_crddrop_inst_cmrg_enable;
	wire [15:0] mem_ctrl_crddrop_flat_crddrop_inst_cmrg_stop_lvl;
	wire mem_ctrl_crddrop_flat_crddrop_inst_tile_en;
	wire mem_ctrl_crdhold_flat_clk;
	wire mem_ctrl_crdhold_flat_cmrg_coord_in_0_ready_f_;
	wire mem_ctrl_crdhold_flat_cmrg_coord_in_1_ready_f_;
	wire [16:0] mem_ctrl_crdhold_flat_cmrg_coord_out_0_f_;
	wire mem_ctrl_crdhold_flat_cmrg_coord_out_0_valid_f_;
	wire [16:0] mem_ctrl_crdhold_flat_cmrg_coord_out_1_f_;
	wire mem_ctrl_crdhold_flat_cmrg_coord_out_1_valid_f_;
	wire mem_ctrl_crdhold_flat_crdhold_inst_cmrg_enable;
	wire [15:0] mem_ctrl_crdhold_flat_crdhold_inst_cmrg_stop_lvl;
	wire mem_ctrl_crdhold_flat_crdhold_inst_tile_en;
	wire mem_ctrl_intersect_unit_flat_clk;
	wire mem_ctrl_intersect_unit_flat_coord_in_0_ready_f_;
	wire mem_ctrl_intersect_unit_flat_coord_in_1_ready_f_;
	wire [16:0] mem_ctrl_intersect_unit_flat_coord_out_f_;
	wire mem_ctrl_intersect_unit_flat_coord_out_valid_f_;
	wire mem_ctrl_intersect_unit_flat_intersect_unit_inst_joiner_op;
	wire mem_ctrl_intersect_unit_flat_intersect_unit_inst_tile_en;
	wire mem_ctrl_intersect_unit_flat_pos_in_0_ready_f_;
	wire mem_ctrl_intersect_unit_flat_pos_in_1_ready_f_;
	wire [16:0] mem_ctrl_intersect_unit_flat_pos_out_0_f_;
	wire mem_ctrl_intersect_unit_flat_pos_out_0_valid_f_;
	wire [16:0] mem_ctrl_intersect_unit_flat_pos_out_1_f_;
	wire mem_ctrl_intersect_unit_flat_pos_out_1_valid_f_;
	wire mem_ctrl_reg_cr_flat_clk;
	wire mem_ctrl_reg_cr_flat_data_in_ready_f_;
	wire [16:0] mem_ctrl_reg_cr_flat_data_out_f_;
	wire mem_ctrl_reg_cr_flat_data_out_valid_f_;
	wire [15:0] mem_ctrl_reg_cr_flat_reg_cr_inst_default_value;
	wire [15:0] mem_ctrl_reg_cr_flat_reg_cr_inst_stop_lvl;
	wire mem_ctrl_reg_cr_flat_reg_cr_inst_tile_en;
	reg [16:0] output_width_17_num_0_fifo_in;
	wire output_width_17_num_0_fifo_in_ready;
	reg output_width_17_num_0_fifo_in_valid;
	wire [16:0] output_width_17_num_0_output_fifo_data_out;
	wire output_width_17_num_0_output_fifo_empty;
	wire output_width_17_num_0_output_fifo_full;
	reg [16:0] output_width_17_num_1_fifo_in;
	wire output_width_17_num_1_fifo_in_ready;
	reg output_width_17_num_1_fifo_in_valid;
	wire [16:0] output_width_17_num_1_output_fifo_data_out;
	wire output_width_17_num_1_output_fifo_empty;
	wire output_width_17_num_1_output_fifo_full;
	reg [16:0] output_width_17_num_2_fifo_in;
	wire output_width_17_num_2_fifo_in_ready;
	reg output_width_17_num_2_fifo_in_valid;
	wire [16:0] output_width_17_num_2_output_fifo_data_out;
	wire output_width_17_num_2_output_fifo_empty;
	wire output_width_17_num_2_output_fifo_full;
	assign gclk = clk & tile_en;
	assign mem_ctrl_intersect_unit_flat_clk = gclk & (mode == 3'h0);
	assign mem_ctrl_crddrop_flat_clk = gclk & (mode == 3'h1);
	assign mem_ctrl_crdhold_flat_clk = gclk & (mode == 3'h2);
	assign mem_ctrl_PE_onyx_flat_clk = gclk & (mode == 3'h3);
	assign mem_ctrl_Repeat_flat_clk = gclk & (mode == 3'h4);
	assign mem_ctrl_RepeatSignalGenerator_flat_clk = gclk & (mode == 3'h5);
	assign mem_ctrl_reg_cr_flat_clk = gclk & (mode == 3'h6);
	assign input_width_17_num_0_fifo_out_valid = ~input_width_17_num_0_input_fifo_empty;
	always @(*) begin
		input_width_17_num_0_fifo_out_ready = 1'h1;
		if (mode == 3'h0)
			input_width_17_num_0_fifo_out_ready = mem_ctrl_intersect_unit_flat_coord_in_0_ready_f_;
		else if (mode == 3'h1)
			input_width_17_num_0_fifo_out_ready = mem_ctrl_crddrop_flat_cmrg_coord_in_0_ready_f_;
		else if (mode == 3'h2)
			input_width_17_num_0_fifo_out_ready = mem_ctrl_crdhold_flat_cmrg_coord_in_0_ready_f_;
		else if (mode == 3'h3)
			input_width_17_num_0_fifo_out_ready = mem_ctrl_PE_onyx_flat_data0_ready_f_;
		else if (mode == 3'h4)
			input_width_17_num_0_fifo_out_ready = mem_ctrl_Repeat_flat_proc_data_in_ready_f_;
		else if (mode == 3'h5)
			input_width_17_num_0_fifo_out_ready = mem_ctrl_RepeatSignalGenerator_flat_base_data_in_ready_f_;
		else if (mode == 3'h6)
			input_width_17_num_0_fifo_out_ready = mem_ctrl_reg_cr_flat_data_in_ready_f_;
	end
	assign mem_ctrl_PE_onyx_flat_data0_f_ = (PE_input_width_17_num_0_dense ? PE_input_width_17_num_0 : input_width_17_num_0_fifo_out);
	assign mem_ctrl_PE_onyx_flat_data0_valid_f_ = (PE_input_width_17_num_0_dense ? 1'h1 : input_width_17_num_0_fifo_out_valid);
	always @(*) begin
		PE_input_width_17_num_0_ready = 1'h1;
		if (mode == 3'h0)
			PE_input_width_17_num_0_ready = ~input_width_17_num_0_input_fifo_full;
		else if (mode == 3'h1)
			PE_input_width_17_num_0_ready = ~input_width_17_num_0_input_fifo_full;
		else if (mode == 3'h2)
			PE_input_width_17_num_0_ready = ~input_width_17_num_0_input_fifo_full;
		else if (mode == 3'h3)
			PE_input_width_17_num_0_ready = (PE_input_width_17_num_0_dense ? 1'h1 : ~input_width_17_num_0_input_fifo_full);
		else if (mode == 3'h4)
			PE_input_width_17_num_0_ready = ~input_width_17_num_0_input_fifo_full;
		else if (mode == 3'h5)
			PE_input_width_17_num_0_ready = ~input_width_17_num_0_input_fifo_full;
		else if (mode == 3'h6)
			PE_input_width_17_num_0_ready = ~input_width_17_num_0_input_fifo_full;
	end
	assign input_width_17_num_1_fifo_out_valid = ~input_width_17_num_1_input_fifo_empty;
	always @(*) begin
		input_width_17_num_1_fifo_out_ready = 1'h1;
		if (mode == 3'h0)
			input_width_17_num_1_fifo_out_ready = mem_ctrl_intersect_unit_flat_coord_in_1_ready_f_;
		else if (mode == 3'h1)
			input_width_17_num_1_fifo_out_ready = mem_ctrl_crddrop_flat_cmrg_coord_in_1_ready_f_;
		else if (mode == 3'h2)
			input_width_17_num_1_fifo_out_ready = mem_ctrl_crdhold_flat_cmrg_coord_in_1_ready_f_;
		else if (mode == 3'h3)
			input_width_17_num_1_fifo_out_ready = mem_ctrl_PE_onyx_flat_data1_ready_f_;
		else if (mode == 3'h4)
			input_width_17_num_1_fifo_out_ready = mem_ctrl_Repeat_flat_repsig_data_in_ready_f_;
	end
	assign mem_ctrl_PE_onyx_flat_data1_f_ = (PE_input_width_17_num_1_dense ? PE_input_width_17_num_1 : input_width_17_num_1_fifo_out);
	assign mem_ctrl_PE_onyx_flat_data1_valid_f_ = (PE_input_width_17_num_1_dense ? 1'h1 : input_width_17_num_1_fifo_out_valid);
	always @(*) begin
		PE_input_width_17_num_1_ready = 1'h1;
		if (mode == 3'h0)
			PE_input_width_17_num_1_ready = ~input_width_17_num_1_input_fifo_full;
		else if (mode == 3'h1)
			PE_input_width_17_num_1_ready = ~input_width_17_num_1_input_fifo_full;
		else if (mode == 3'h2)
			PE_input_width_17_num_1_ready = ~input_width_17_num_1_input_fifo_full;
		else if (mode == 3'h3)
			PE_input_width_17_num_1_ready = (PE_input_width_17_num_1_dense ? 1'h1 : ~input_width_17_num_1_input_fifo_full);
		else if (mode == 3'h4)
			PE_input_width_17_num_1_ready = ~input_width_17_num_1_input_fifo_full;
	end
	assign input_width_17_num_2_fifo_out_valid = ~input_width_17_num_2_input_fifo_empty;
	always @(*) begin
		input_width_17_num_2_fifo_out_ready = 1'h1;
		if (mode == 3'h0)
			input_width_17_num_2_fifo_out_ready = mem_ctrl_intersect_unit_flat_pos_in_0_ready_f_;
		else
			input_width_17_num_2_fifo_out_ready = 1'h1;
	end
	always @(*) begin
		PE_input_width_17_num_2_ready = 1'h1;
		if (mode == 3'h0)
			PE_input_width_17_num_2_ready = ~input_width_17_num_2_input_fifo_full;
		else if (mode == 3'h3)
			PE_input_width_17_num_2_ready = 1'h1;
	end
	assign input_width_17_num_3_fifo_out_valid = ~input_width_17_num_3_input_fifo_empty;
	always @(*) begin
		input_width_17_num_3_fifo_out_ready = 1'h1;
		if (mode == 3'h0)
			input_width_17_num_3_fifo_out_ready = mem_ctrl_intersect_unit_flat_pos_in_1_ready_f_;
		else
			input_width_17_num_3_fifo_out_ready = 1'h1;
	end
	always @(*) begin
		PE_input_width_17_num_3_ready = 1'h1;
		if (mode == 3'h0)
			PE_input_width_17_num_3_ready = ~input_width_17_num_3_input_fifo_full;
		else
			PE_input_width_17_num_3_ready = 1'h1;
	end
	assign output_width_17_num_0_fifo_in_ready = ~output_width_17_num_0_output_fifo_full;
	always @(*) begin
		output_width_17_num_0_fifo_in = 17'h00000;
		output_width_17_num_0_fifo_in_valid = 1'h0;
		if (mode == 3'h0) begin
			output_width_17_num_0_fifo_in = mem_ctrl_intersect_unit_flat_coord_out_f_;
			output_width_17_num_0_fifo_in_valid = mem_ctrl_intersect_unit_flat_coord_out_valid_f_;
		end
		else if (mode == 3'h1) begin
			output_width_17_num_0_fifo_in = mem_ctrl_crddrop_flat_cmrg_coord_out_0_f_;
			output_width_17_num_0_fifo_in_valid = mem_ctrl_crddrop_flat_cmrg_coord_out_0_valid_f_;
		end
		else if (mode == 3'h2) begin
			output_width_17_num_0_fifo_in = mem_ctrl_crdhold_flat_cmrg_coord_out_0_f_;
			output_width_17_num_0_fifo_in_valid = mem_ctrl_crdhold_flat_cmrg_coord_out_0_valid_f_;
		end
		else if (mode == 3'h3) begin
			output_width_17_num_0_fifo_in = mem_ctrl_PE_onyx_flat_res_f_;
			output_width_17_num_0_fifo_in_valid = mem_ctrl_PE_onyx_flat_res_valid_f_;
		end
		else if (mode == 3'h4) begin
			output_width_17_num_0_fifo_in = mem_ctrl_Repeat_flat_ref_data_out_f_;
			output_width_17_num_0_fifo_in_valid = mem_ctrl_Repeat_flat_ref_data_out_valid_f_;
		end
		else if (mode == 3'h5) begin
			output_width_17_num_0_fifo_in = mem_ctrl_RepeatSignalGenerator_flat_repsig_data_out_f_;
			output_width_17_num_0_fifo_in_valid = mem_ctrl_RepeatSignalGenerator_flat_repsig_data_out_valid_f_;
		end
		else if (mode == 3'h6) begin
			output_width_17_num_0_fifo_in = mem_ctrl_reg_cr_flat_data_out_f_;
			output_width_17_num_0_fifo_in_valid = mem_ctrl_reg_cr_flat_data_out_valid_f_;
		end
	end
	assign mem_ctrl_PE_onyx_flat_res_ready_f_ = (PE_output_width_17_num_0_dense ? 1'h1 : output_width_17_num_0_fifo_in_ready);
	always @(*) begin
		PE_output_width_17_num_0 = 17'h00000;
		if (mode == 3'h0)
			PE_output_width_17_num_0 = output_width_17_num_0_output_fifo_data_out;
		else if (mode == 3'h1)
			PE_output_width_17_num_0 = output_width_17_num_0_output_fifo_data_out;
		else if (mode == 3'h2)
			PE_output_width_17_num_0 = output_width_17_num_0_output_fifo_data_out;
		else if (mode == 3'h3)
			PE_output_width_17_num_0 = (PE_output_width_17_num_0_dense ? mem_ctrl_PE_onyx_flat_res_f_ : output_width_17_num_0_output_fifo_data_out);
		else if (mode == 3'h4)
			PE_output_width_17_num_0 = output_width_17_num_0_output_fifo_data_out;
		else if (mode == 3'h5)
			PE_output_width_17_num_0 = output_width_17_num_0_output_fifo_data_out;
		else if (mode == 3'h6)
			PE_output_width_17_num_0 = output_width_17_num_0_output_fifo_data_out;
	end
	always @(*) begin
		PE_output_width_17_num_0_valid = 1'h0;
		if (mode == 3'h0)
			PE_output_width_17_num_0_valid = ~output_width_17_num_0_output_fifo_empty;
		else if (mode == 3'h1)
			PE_output_width_17_num_0_valid = ~output_width_17_num_0_output_fifo_empty;
		else if (mode == 3'h2)
			PE_output_width_17_num_0_valid = ~output_width_17_num_0_output_fifo_empty;
		else if (mode == 3'h3)
			PE_output_width_17_num_0_valid = (PE_output_width_17_num_0_dense ? 1'h1 : ~output_width_17_num_0_output_fifo_empty);
		else if (mode == 3'h4)
			PE_output_width_17_num_0_valid = ~output_width_17_num_0_output_fifo_empty;
		else if (mode == 3'h5)
			PE_output_width_17_num_0_valid = ~output_width_17_num_0_output_fifo_empty;
		else if (mode == 3'h6)
			PE_output_width_17_num_0_valid = ~output_width_17_num_0_output_fifo_empty;
	end
	assign output_width_17_num_1_fifo_in_ready = ~output_width_17_num_1_output_fifo_full;
	always @(*) begin
		output_width_17_num_1_fifo_in = 17'h00000;
		output_width_17_num_1_fifo_in_valid = 1'h0;
		if (mode == 3'h0) begin
			output_width_17_num_1_fifo_in = mem_ctrl_intersect_unit_flat_pos_out_0_f_;
			output_width_17_num_1_fifo_in_valid = mem_ctrl_intersect_unit_flat_pos_out_0_valid_f_;
		end
		else if (mode == 3'h1) begin
			output_width_17_num_1_fifo_in = mem_ctrl_crddrop_flat_cmrg_coord_out_1_f_;
			output_width_17_num_1_fifo_in_valid = mem_ctrl_crddrop_flat_cmrg_coord_out_1_valid_f_;
		end
		else if (mode == 3'h2) begin
			output_width_17_num_1_fifo_in = mem_ctrl_crdhold_flat_cmrg_coord_out_1_f_;
			output_width_17_num_1_fifo_in_valid = mem_ctrl_crdhold_flat_cmrg_coord_out_1_valid_f_;
		end
	end
	always @(*) begin
		PE_output_width_17_num_1 = 17'h00000;
		if (mode == 3'h0)
			PE_output_width_17_num_1 = output_width_17_num_1_output_fifo_data_out;
		else if (mode == 3'h1)
			PE_output_width_17_num_1 = output_width_17_num_1_output_fifo_data_out;
		else if (mode == 3'h2)
			PE_output_width_17_num_1 = output_width_17_num_1_output_fifo_data_out;
	end
	always @(*) begin
		PE_output_width_17_num_1_valid = 1'h0;
		if (mode == 3'h0)
			PE_output_width_17_num_1_valid = ~output_width_17_num_1_output_fifo_empty;
		else if (mode == 3'h1)
			PE_output_width_17_num_1_valid = ~output_width_17_num_1_output_fifo_empty;
		else if (mode == 3'h2)
			PE_output_width_17_num_1_valid = ~output_width_17_num_1_output_fifo_empty;
	end
	assign output_width_17_num_2_fifo_in_ready = ~output_width_17_num_2_output_fifo_full;
	always @(*) begin
		output_width_17_num_2_fifo_in = 17'h00000;
		output_width_17_num_2_fifo_in_valid = 1'h0;
		output_width_17_num_2_fifo_in = mem_ctrl_intersect_unit_flat_pos_out_1_f_;
		output_width_17_num_2_fifo_in_valid = mem_ctrl_intersect_unit_flat_pos_out_1_valid_f_;
	end
	always @(*) begin
		PE_output_width_17_num_2 = 17'h00000;
		if (mode == 3'h0)
			PE_output_width_17_num_2 = output_width_17_num_2_output_fifo_data_out;
		else
			PE_output_width_17_num_2 = 17'h00000;
	end
	always @(*) begin
		PE_output_width_17_num_2_valid = 1'h0;
		if (mode == 3'h0)
			PE_output_width_17_num_2_valid = ~output_width_17_num_2_output_fifo_empty;
		else
			PE_output_width_17_num_2_valid = 1'h0;
	end
	always @(*) begin
		PE_output_width_1_num_0 = 1'h0;
		if (mode == 3'h3)
			PE_output_width_1_num_0 = mem_ctrl_PE_onyx_flat_res_p_f_;
		else
			PE_output_width_1_num_0 = 1'h0;
	end
	assign {mem_ctrl_intersect_unit_flat_intersect_unit_inst_joiner_op, mem_ctrl_intersect_unit_flat_intersect_unit_inst_tile_en} = CONFIG_SPACE[1:0];
	assign {mem_ctrl_crddrop_flat_crddrop_inst_cmrg_enable, mem_ctrl_crddrop_flat_crddrop_inst_cmrg_stop_lvl, mem_ctrl_crddrop_flat_crddrop_inst_tile_en} = CONFIG_SPACE[17:0];
	assign {mem_ctrl_crdhold_flat_crdhold_inst_cmrg_enable, mem_ctrl_crdhold_flat_crdhold_inst_cmrg_stop_lvl, mem_ctrl_crdhold_flat_crdhold_inst_tile_en} = CONFIG_SPACE[17:0];
	assign {mem_ctrl_PE_onyx_flat_PE_onyx_inst_dense_mode, mem_ctrl_PE_onyx_flat_PE_onyx_inst_onyxpeintf_inst, mem_ctrl_PE_onyx_flat_PE_onyx_inst_tile_en} = CONFIG_SPACE[85:0];
	assign {mem_ctrl_Repeat_flat_Repeat_inst_root, mem_ctrl_Repeat_flat_Repeat_inst_spacc_mode, mem_ctrl_Repeat_flat_Repeat_inst_stop_lvl, mem_ctrl_Repeat_flat_Repeat_inst_tile_en} = CONFIG_SPACE[18:0];
	assign {mem_ctrl_RepeatSignalGenerator_flat_RepeatSignalGenerator_inst_stop_lvl, mem_ctrl_RepeatSignalGenerator_flat_RepeatSignalGenerator_inst_tile_en} = CONFIG_SPACE[16:0];
	assign {mem_ctrl_reg_cr_flat_reg_cr_inst_default_value, mem_ctrl_reg_cr_flat_reg_cr_inst_stop_lvl, mem_ctrl_reg_cr_flat_reg_cr_inst_tile_en} = CONFIG_SPACE[32:0];
	assign CONFIG_SPACE[31:0] = CONFIG_SPACE_0;
	assign CONFIG_SPACE[63:32] = CONFIG_SPACE_1;
	assign CONFIG_SPACE[85:64] = CONFIG_SPACE_2;
	intersect_unit_flat mem_ctrl_intersect_unit_flat(
		.clk(mem_ctrl_intersect_unit_flat_clk),
		.clk_en(clk_en),
		.coord_in_0_f_(input_width_17_num_0_fifo_out),
		.coord_in_0_valid_f_(input_width_17_num_0_fifo_out_valid),
		.coord_in_1_f_(input_width_17_num_1_fifo_out),
		.coord_in_1_valid_f_(input_width_17_num_1_fifo_out_valid),
		.coord_out_ready_f_(output_width_17_num_0_fifo_in_ready),
		.flush(flush),
		.intersect_unit_inst_joiner_op(mem_ctrl_intersect_unit_flat_intersect_unit_inst_joiner_op),
		.intersect_unit_inst_tile_en(mem_ctrl_intersect_unit_flat_intersect_unit_inst_tile_en),
		.pos_in_0_f_(input_width_17_num_2_fifo_out),
		.pos_in_0_valid_f_(input_width_17_num_2_fifo_out_valid),
		.pos_in_1_f_(input_width_17_num_3_fifo_out),
		.pos_in_1_valid_f_(input_width_17_num_3_fifo_out_valid),
		.pos_out_0_ready_f_(output_width_17_num_1_fifo_in_ready),
		.pos_out_1_ready_f_(output_width_17_num_2_fifo_in_ready),
		.rst_n(rst_n),
		.coord_in_0_ready_f_(mem_ctrl_intersect_unit_flat_coord_in_0_ready_f_),
		.coord_in_1_ready_f_(mem_ctrl_intersect_unit_flat_coord_in_1_ready_f_),
		.coord_out_f_(mem_ctrl_intersect_unit_flat_coord_out_f_),
		.coord_out_valid_f_(mem_ctrl_intersect_unit_flat_coord_out_valid_f_),
		.pos_in_0_ready_f_(mem_ctrl_intersect_unit_flat_pos_in_0_ready_f_),
		.pos_in_1_ready_f_(mem_ctrl_intersect_unit_flat_pos_in_1_ready_f_),
		.pos_out_0_f_(mem_ctrl_intersect_unit_flat_pos_out_0_f_),
		.pos_out_0_valid_f_(mem_ctrl_intersect_unit_flat_pos_out_0_valid_f_),
		.pos_out_1_f_(mem_ctrl_intersect_unit_flat_pos_out_1_f_),
		.pos_out_1_valid_f_(mem_ctrl_intersect_unit_flat_pos_out_1_valid_f_)
	);
	crddrop_flat mem_ctrl_crddrop_flat(
		.clk(mem_ctrl_crddrop_flat_clk),
		.clk_en(clk_en),
		.cmrg_coord_in_0_f_(input_width_17_num_0_fifo_out),
		.cmrg_coord_in_0_valid_f_(input_width_17_num_0_fifo_out_valid),
		.cmrg_coord_in_1_f_(input_width_17_num_1_fifo_out),
		.cmrg_coord_in_1_valid_f_(input_width_17_num_1_fifo_out_valid),
		.cmrg_coord_out_0_ready_f_(output_width_17_num_0_fifo_in_ready),
		.cmrg_coord_out_1_ready_f_(output_width_17_num_1_fifo_in_ready),
		.crddrop_inst_cmrg_enable(mem_ctrl_crddrop_flat_crddrop_inst_cmrg_enable),
		.crddrop_inst_cmrg_stop_lvl(mem_ctrl_crddrop_flat_crddrop_inst_cmrg_stop_lvl),
		.crddrop_inst_tile_en(mem_ctrl_crddrop_flat_crddrop_inst_tile_en),
		.flush(flush),
		.rst_n(rst_n),
		.cmrg_coord_in_0_ready_f_(mem_ctrl_crddrop_flat_cmrg_coord_in_0_ready_f_),
		.cmrg_coord_in_1_ready_f_(mem_ctrl_crddrop_flat_cmrg_coord_in_1_ready_f_),
		.cmrg_coord_out_0_f_(mem_ctrl_crddrop_flat_cmrg_coord_out_0_f_),
		.cmrg_coord_out_0_valid_f_(mem_ctrl_crddrop_flat_cmrg_coord_out_0_valid_f_),
		.cmrg_coord_out_1_f_(mem_ctrl_crddrop_flat_cmrg_coord_out_1_f_),
		.cmrg_coord_out_1_valid_f_(mem_ctrl_crddrop_flat_cmrg_coord_out_1_valid_f_)
	);
	crdhold_flat mem_ctrl_crdhold_flat(
		.clk(mem_ctrl_crdhold_flat_clk),
		.clk_en(clk_en),
		.cmrg_coord_in_0_f_(input_width_17_num_0_fifo_out),
		.cmrg_coord_in_0_valid_f_(input_width_17_num_0_fifo_out_valid),
		.cmrg_coord_in_1_f_(input_width_17_num_1_fifo_out),
		.cmrg_coord_in_1_valid_f_(input_width_17_num_1_fifo_out_valid),
		.cmrg_coord_out_0_ready_f_(output_width_17_num_0_fifo_in_ready),
		.cmrg_coord_out_1_ready_f_(output_width_17_num_1_fifo_in_ready),
		.crdhold_inst_cmrg_enable(mem_ctrl_crdhold_flat_crdhold_inst_cmrg_enable),
		.crdhold_inst_cmrg_stop_lvl(mem_ctrl_crdhold_flat_crdhold_inst_cmrg_stop_lvl),
		.crdhold_inst_tile_en(mem_ctrl_crdhold_flat_crdhold_inst_tile_en),
		.flush(flush),
		.rst_n(rst_n),
		.cmrg_coord_in_0_ready_f_(mem_ctrl_crdhold_flat_cmrg_coord_in_0_ready_f_),
		.cmrg_coord_in_1_ready_f_(mem_ctrl_crdhold_flat_cmrg_coord_in_1_ready_f_),
		.cmrg_coord_out_0_f_(mem_ctrl_crdhold_flat_cmrg_coord_out_0_f_),
		.cmrg_coord_out_0_valid_f_(mem_ctrl_crdhold_flat_cmrg_coord_out_0_valid_f_),
		.cmrg_coord_out_1_f_(mem_ctrl_crdhold_flat_cmrg_coord_out_1_f_),
		.cmrg_coord_out_1_valid_f_(mem_ctrl_crdhold_flat_cmrg_coord_out_1_valid_f_)
	);
	PE_onyx_flat mem_ctrl_PE_onyx_flat(
		.PE_onyx_inst_dense_mode(mem_ctrl_PE_onyx_flat_PE_onyx_inst_dense_mode),
		.PE_onyx_inst_onyxpeintf_inst(mem_ctrl_PE_onyx_flat_PE_onyx_inst_onyxpeintf_inst),
		.PE_onyx_inst_tile_en(mem_ctrl_PE_onyx_flat_PE_onyx_inst_tile_en),
		.bit0_f_(PE_input_width_1_num_0),
		.bit1_f_(PE_input_width_1_num_1),
		.bit2_f_(PE_input_width_1_num_2),
		.clk(mem_ctrl_PE_onyx_flat_clk),
		.clk_en(clk_en),
		.data0_f_(mem_ctrl_PE_onyx_flat_data0_f_),
		.data0_valid_f_(mem_ctrl_PE_onyx_flat_data0_valid_f_),
		.data1_f_(mem_ctrl_PE_onyx_flat_data1_f_),
		.data1_valid_f_(mem_ctrl_PE_onyx_flat_data1_valid_f_),
		.data2_f_(PE_input_width_17_num_2),
		.flush(flush),
		.res_ready_f_(mem_ctrl_PE_onyx_flat_res_ready_f_),
		.rst_n(rst_n),
		.PE_onyx_inst_onyxpeintf_O2(PE_onyx_inst_onyxpeintf_O2),
		.PE_onyx_inst_onyxpeintf_O3(PE_onyx_inst_onyxpeintf_O3),
		.PE_onyx_inst_onyxpeintf_O4(PE_onyx_inst_onyxpeintf_O4),
		.data0_ready_f_(mem_ctrl_PE_onyx_flat_data0_ready_f_),
		.data1_ready_f_(mem_ctrl_PE_onyx_flat_data1_ready_f_),
		.res_f_(mem_ctrl_PE_onyx_flat_res_f_),
		.res_p_f_(mem_ctrl_PE_onyx_flat_res_p_f_),
		.res_valid_f_(mem_ctrl_PE_onyx_flat_res_valid_f_)
	);
	Repeat_flat mem_ctrl_Repeat_flat(
		.Repeat_inst_root(mem_ctrl_Repeat_flat_Repeat_inst_root),
		.Repeat_inst_spacc_mode(mem_ctrl_Repeat_flat_Repeat_inst_spacc_mode),
		.Repeat_inst_stop_lvl(mem_ctrl_Repeat_flat_Repeat_inst_stop_lvl),
		.Repeat_inst_tile_en(mem_ctrl_Repeat_flat_Repeat_inst_tile_en),
		.clk(mem_ctrl_Repeat_flat_clk),
		.clk_en(clk_en),
		.flush(flush),
		.proc_data_in_f_(input_width_17_num_0_fifo_out),
		.proc_data_in_valid_f_(input_width_17_num_0_fifo_out_valid),
		.ref_data_out_ready_f_(output_width_17_num_0_fifo_in_ready),
		.repsig_data_in_f_(input_width_17_num_1_fifo_out),
		.repsig_data_in_valid_f_(input_width_17_num_1_fifo_out_valid),
		.rst_n(rst_n),
		.proc_data_in_ready_f_(mem_ctrl_Repeat_flat_proc_data_in_ready_f_),
		.ref_data_out_f_(mem_ctrl_Repeat_flat_ref_data_out_f_),
		.ref_data_out_valid_f_(mem_ctrl_Repeat_flat_ref_data_out_valid_f_),
		.repsig_data_in_ready_f_(mem_ctrl_Repeat_flat_repsig_data_in_ready_f_)
	);
	RepeatSignalGenerator_flat mem_ctrl_RepeatSignalGenerator_flat(
		.RepeatSignalGenerator_inst_stop_lvl(mem_ctrl_RepeatSignalGenerator_flat_RepeatSignalGenerator_inst_stop_lvl),
		.RepeatSignalGenerator_inst_tile_en(mem_ctrl_RepeatSignalGenerator_flat_RepeatSignalGenerator_inst_tile_en),
		.base_data_in_f_(input_width_17_num_0_fifo_out),
		.base_data_in_valid_f_(input_width_17_num_0_fifo_out_valid),
		.clk(mem_ctrl_RepeatSignalGenerator_flat_clk),
		.clk_en(clk_en),
		.flush(flush),
		.repsig_data_out_ready_f_(output_width_17_num_0_fifo_in_ready),
		.rst_n(rst_n),
		.base_data_in_ready_f_(mem_ctrl_RepeatSignalGenerator_flat_base_data_in_ready_f_),
		.repsig_data_out_f_(mem_ctrl_RepeatSignalGenerator_flat_repsig_data_out_f_),
		.repsig_data_out_valid_f_(mem_ctrl_RepeatSignalGenerator_flat_repsig_data_out_valid_f_)
	);
	reg_cr_flat mem_ctrl_reg_cr_flat(
		.clk(mem_ctrl_reg_cr_flat_clk),
		.clk_en(clk_en),
		.data_in_f_(input_width_17_num_0_fifo_out),
		.data_in_valid_f_(input_width_17_num_0_fifo_out_valid),
		.data_out_ready_f_(output_width_17_num_0_fifo_in_ready),
		.flush(flush),
		.reg_cr_inst_default_value(mem_ctrl_reg_cr_flat_reg_cr_inst_default_value),
		.reg_cr_inst_stop_lvl(mem_ctrl_reg_cr_flat_reg_cr_inst_stop_lvl),
		.reg_cr_inst_tile_en(mem_ctrl_reg_cr_flat_reg_cr_inst_tile_en),
		.rst_n(rst_n),
		.data_in_ready_f_(mem_ctrl_reg_cr_flat_data_in_ready_f_),
		.data_out_f_(mem_ctrl_reg_cr_flat_data_out_f_),
		.data_out_valid_f_(mem_ctrl_reg_cr_flat_data_out_valid_f_)
	);
	reg_fifo_depth_2_w_17_afd_2 input_width_17_num_0_input_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(PE_input_width_17_num_0),
		.flush(flush),
		.pop(input_width_17_num_0_fifo_out_ready),
		.push(PE_input_width_17_num_0_valid),
		.rst_n(rst_n),
		.data_out(input_width_17_num_0_fifo_out),
		.empty(input_width_17_num_0_input_fifo_empty),
		.full(input_width_17_num_0_input_fifo_full)
	);
	reg_fifo_depth_2_w_17_afd_2 input_width_17_num_1_input_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(PE_input_width_17_num_1),
		.flush(flush),
		.pop(input_width_17_num_1_fifo_out_ready),
		.push(PE_input_width_17_num_1_valid),
		.rst_n(rst_n),
		.data_out(input_width_17_num_1_fifo_out),
		.empty(input_width_17_num_1_input_fifo_empty),
		.full(input_width_17_num_1_input_fifo_full)
	);
	reg_fifo_depth_2_w_17_afd_2 input_width_17_num_2_input_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(PE_input_width_17_num_2),
		.flush(flush),
		.pop(input_width_17_num_2_fifo_out_ready),
		.push(PE_input_width_17_num_2_valid),
		.rst_n(rst_n),
		.data_out(input_width_17_num_2_fifo_out),
		.empty(input_width_17_num_2_input_fifo_empty),
		.full(input_width_17_num_2_input_fifo_full)
	);
	reg_fifo_depth_2_w_17_afd_2 input_width_17_num_3_input_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(PE_input_width_17_num_3),
		.flush(flush),
		.pop(input_width_17_num_3_fifo_out_ready),
		.push(PE_input_width_17_num_3_valid),
		.rst_n(rst_n),
		.data_out(input_width_17_num_3_fifo_out),
		.empty(input_width_17_num_3_input_fifo_empty),
		.full(input_width_17_num_3_input_fifo_full)
	);
	reg_fifo_depth_2_w_17_afd_2 output_width_17_num_0_output_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(output_width_17_num_0_fifo_in),
		.flush(flush),
		.pop(PE_output_width_17_num_0_ready),
		.push(output_width_17_num_0_fifo_in_valid),
		.rst_n(rst_n),
		.data_out(output_width_17_num_0_output_fifo_data_out),
		.empty(output_width_17_num_0_output_fifo_empty),
		.full(output_width_17_num_0_output_fifo_full)
	);
	reg_fifo_depth_2_w_17_afd_2 output_width_17_num_1_output_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(output_width_17_num_1_fifo_in),
		.flush(flush),
		.pop(PE_output_width_17_num_1_ready),
		.push(output_width_17_num_1_fifo_in_valid),
		.rst_n(rst_n),
		.data_out(output_width_17_num_1_output_fifo_data_out),
		.empty(output_width_17_num_1_output_fifo_empty),
		.full(output_width_17_num_1_output_fifo_full)
	);
	reg_fifo_depth_2_w_17_afd_2 output_width_17_num_2_output_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(output_width_17_num_2_fifo_in),
		.flush(flush),
		.pop(PE_output_width_17_num_2_ready),
		.push(output_width_17_num_2_fifo_in_valid),
		.rst_n(rst_n),
		.data_out(output_width_17_num_2_output_fifo_data_out),
		.empty(output_width_17_num_2_output_fifo_empty),
		.full(output_width_17_num_2_output_fifo_full)
	);
endmodule
module PE_inner_W (
	CONFIG_SPACE_0,
	CONFIG_SPACE_1,
	CONFIG_SPACE_2,
	PE_input_width_17_num_0,
	PE_input_width_17_num_0_dense,
	PE_input_width_17_num_0_valid,
	PE_input_width_17_num_1,
	PE_input_width_17_num_1_dense,
	PE_input_width_17_num_1_valid,
	PE_input_width_17_num_2,
	PE_input_width_17_num_2_valid,
	PE_input_width_17_num_3,
	PE_input_width_17_num_3_valid,
	PE_input_width_1_num_0,
	PE_input_width_1_num_1,
	PE_input_width_1_num_2,
	PE_output_width_17_num_0_dense,
	PE_output_width_17_num_0_ready,
	PE_output_width_17_num_1_ready,
	PE_output_width_17_num_2_ready,
	clk,
	clk_en,
	flush,
	mode,
	rst_n,
	tile_en,
	PE_input_width_17_num_0_ready,
	PE_input_width_17_num_1_ready,
	PE_input_width_17_num_2_ready,
	PE_input_width_17_num_3_ready,
	PE_onyx_inst_onyxpeintf_O2,
	PE_onyx_inst_onyxpeintf_O3,
	PE_onyx_inst_onyxpeintf_O4,
	PE_output_width_17_num_0,
	PE_output_width_17_num_0_valid,
	PE_output_width_17_num_1,
	PE_output_width_17_num_1_valid,
	PE_output_width_17_num_2,
	PE_output_width_17_num_2_valid,
	PE_output_width_1_num_0
);
	input wire [31:0] CONFIG_SPACE_0;
	input wire [31:0] CONFIG_SPACE_1;
	input wire [21:0] CONFIG_SPACE_2;
	input wire [16:0] PE_input_width_17_num_0;
	input wire PE_input_width_17_num_0_dense;
	input wire PE_input_width_17_num_0_valid;
	input wire [16:0] PE_input_width_17_num_1;
	input wire PE_input_width_17_num_1_dense;
	input wire PE_input_width_17_num_1_valid;
	input wire [16:0] PE_input_width_17_num_2;
	input wire PE_input_width_17_num_2_valid;
	input wire [16:0] PE_input_width_17_num_3;
	input wire PE_input_width_17_num_3_valid;
	input wire PE_input_width_1_num_0;
	input wire PE_input_width_1_num_1;
	input wire PE_input_width_1_num_2;
	input wire PE_output_width_17_num_0_dense;
	input wire PE_output_width_17_num_0_ready;
	input wire PE_output_width_17_num_1_ready;
	input wire PE_output_width_17_num_2_ready;
	input wire clk;
	input wire clk_en;
	input wire flush;
	input wire [2:0] mode;
	input wire rst_n;
	input wire tile_en;
	output wire PE_input_width_17_num_0_ready;
	output wire PE_input_width_17_num_1_ready;
	output wire PE_input_width_17_num_2_ready;
	output wire PE_input_width_17_num_3_ready;
	output wire [15:0] PE_onyx_inst_onyxpeintf_O2;
	output wire [15:0] PE_onyx_inst_onyxpeintf_O3;
	output wire [15:0] PE_onyx_inst_onyxpeintf_O4;
	output wire [16:0] PE_output_width_17_num_0;
	output wire PE_output_width_17_num_0_valid;
	output wire [16:0] PE_output_width_17_num_1;
	output wire PE_output_width_17_num_1_valid;
	output wire [16:0] PE_output_width_17_num_2;
	output wire PE_output_width_17_num_2_valid;
	output wire PE_output_width_1_num_0;
	PE_inner PE_inner(
		.CONFIG_SPACE_0(CONFIG_SPACE_0),
		.CONFIG_SPACE_1(CONFIG_SPACE_1),
		.CONFIG_SPACE_2(CONFIG_SPACE_2),
		.PE_input_width_17_num_0(PE_input_width_17_num_0),
		.PE_input_width_17_num_0_dense(PE_input_width_17_num_0_dense),
		.PE_input_width_17_num_0_valid(PE_input_width_17_num_0_valid),
		.PE_input_width_17_num_1(PE_input_width_17_num_1),
		.PE_input_width_17_num_1_dense(PE_input_width_17_num_1_dense),
		.PE_input_width_17_num_1_valid(PE_input_width_17_num_1_valid),
		.PE_input_width_17_num_2(PE_input_width_17_num_2),
		.PE_input_width_17_num_2_valid(PE_input_width_17_num_2_valid),
		.PE_input_width_17_num_3(PE_input_width_17_num_3),
		.PE_input_width_17_num_3_valid(PE_input_width_17_num_3_valid),
		.PE_input_width_1_num_0(PE_input_width_1_num_0),
		.PE_input_width_1_num_1(PE_input_width_1_num_1),
		.PE_input_width_1_num_2(PE_input_width_1_num_2),
		.PE_output_width_17_num_0_dense(PE_output_width_17_num_0_dense),
		.PE_output_width_17_num_0_ready(PE_output_width_17_num_0_ready),
		.PE_output_width_17_num_1_ready(PE_output_width_17_num_1_ready),
		.PE_output_width_17_num_2_ready(PE_output_width_17_num_2_ready),
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.mode(mode),
		.rst_n(rst_n),
		.tile_en(tile_en),
		.PE_input_width_17_num_0_ready(PE_input_width_17_num_0_ready),
		.PE_input_width_17_num_1_ready(PE_input_width_17_num_1_ready),
		.PE_input_width_17_num_2_ready(PE_input_width_17_num_2_ready),
		.PE_input_width_17_num_3_ready(PE_input_width_17_num_3_ready),
		.PE_onyx_inst_onyxpeintf_O2(PE_onyx_inst_onyxpeintf_O2),
		.PE_onyx_inst_onyxpeintf_O3(PE_onyx_inst_onyxpeintf_O3),
		.PE_onyx_inst_onyxpeintf_O4(PE_onyx_inst_onyxpeintf_O4),
		.PE_output_width_17_num_0(PE_output_width_17_num_0),
		.PE_output_width_17_num_0_valid(PE_output_width_17_num_0_valid),
		.PE_output_width_17_num_1(PE_output_width_17_num_1),
		.PE_output_width_17_num_1_valid(PE_output_width_17_num_1_valid),
		.PE_output_width_17_num_2(PE_output_width_17_num_2),
		.PE_output_width_17_num_2_valid(PE_output_width_17_num_2_valid),
		.PE_output_width_1_num_0(PE_output_width_1_num_0)
	);
endmodule
module PE_onyx (
	bit0,
	bit1,
	bit2,
	clk,
	clk_en,
	data0,
	data0_valid,
	data1,
	data1_valid,
	data2,
	dense_mode,
	flush,
	onyxpeintf_inst,
	res_ready,
	rst_n,
	tile_en,
	data0_ready,
	data1_ready,
	onyxpeintf_O2,
	onyxpeintf_O3,
	onyxpeintf_O4,
	res,
	res_p,
	res_valid
);
	input wire bit0;
	input wire bit1;
	input wire bit2;
	input wire clk;
	input wire clk_en;
	input wire [16:0] data0;
	input wire data0_valid;
	input wire [16:0] data1;
	input wire data1_valid;
	input wire [16:0] data2;
	input wire dense_mode;
	input wire flush;
	input wire [83:0] onyxpeintf_inst;
	input wire res_ready;
	input wire rst_n;
	input wire tile_en;
	output wire data0_ready;
	output wire data1_ready;
	output wire [15:0] onyxpeintf_O2;
	output wire [15:0] onyxpeintf_O3;
	output wire [15:0] onyxpeintf_O4;
	output wire [16:0] res;
	output wire res_p;
	output wire res_valid;
	reg [15:0] data_to_fifo;
	wire gclk;
	wire [33:0] infifo_in_packed;
	wire [31:0] infifo_out_data;
	wire [1:0] infifo_out_eos;
	wire infifo_out_maybe_0;
	wire infifo_out_maybe_1;
	wire [33:0] infifo_out_packed;
	wire [1:0] infifo_out_valid;
	reg [1:0] infifo_pop;
	wire infifo_push_0;
	wire infifo_push_1;
	wire [16:0] input_fifo_0_data_out;
	wire input_fifo_0_empty;
	wire input_fifo_0_full;
	wire [16:0] input_fifo_1_data_out;
	wire input_fifo_1_empty;
	wire input_fifo_1_full;
	wire onyxpeintf_ASYNCRESET;
	wire [15:0] onyxpeintf_data0;
	wire [15:0] onyxpeintf_data1;
	wire outfifo_full;
	reg outfifo_in_eos;
	wire [16:0] outfifo_in_packed;
	wire [16:0] outfifo_out_packed;
	wire outfifo_pop;
	reg outfifo_push;
	wire output_fifo_empty;
	wire [15:0] pe_output;
	assign gclk = clk & tile_en;
	assign data0_ready = (dense_mode ? 1'h1 : ~input_fifo_0_full);
	assign data1_ready = (dense_mode ? 1'h1 : ~input_fifo_1_full);
	assign infifo_in_packed[0+:17] = data0;
	assign infifo_out_eos[0] = infifo_out_packed[16];
	assign infifo_out_data[0+:16] = infifo_out_packed[15-:16];
	assign infifo_in_packed[17+:17] = data1;
	assign infifo_out_eos[1] = infifo_out_packed[33];
	assign infifo_out_data[16+:16] = infifo_out_packed[32-:16];
	assign infifo_push_0 = data0_valid;
	assign infifo_push_1 = data1_valid;
	assign infifo_out_packed[0+:17] = input_fifo_0_data_out;
	assign infifo_out_packed[17+:17] = input_fifo_1_data_out;
	assign infifo_out_valid[0] = ~input_fifo_0_empty;
	assign infifo_out_valid[1] = ~input_fifo_1_empty;
	assign outfifo_in_packed[16] = outfifo_in_eos;
	assign outfifo_in_packed[15:0] = data_to_fifo;
	function automatic [16:0] sv2v_cast_17;
		input reg [16:0] inp;
		sv2v_cast_17 = inp;
	endfunction
	assign res = (dense_mode ? sv2v_cast_17(pe_output) : outfifo_out_packed);
	assign res_valid = (dense_mode ? 1'h1 : ~output_fifo_empty);
	assign outfifo_pop = res_ready;
	assign infifo_out_maybe_0 = (infifo_out_eos[0] & infifo_out_valid[0]) & (infifo_out_data[9-:2] == 2'h2);
	assign infifo_out_maybe_1 = (infifo_out_eos[1] & infifo_out_valid[1]) & (infifo_out_data[25-:2] == 2'h2);
	assign onyxpeintf_ASYNCRESET = ~rst_n;
	assign onyxpeintf_data0 = (dense_mode ? data0[15:0] : (infifo_out_maybe_0 ? 16'h0000 : infifo_out_data[0+:16]));
	assign onyxpeintf_data1 = (dense_mode ? data1[15:0] : (infifo_out_maybe_1 ? 16'h0000 : infifo_out_data[16+:16]));
	always @(*) begin
		outfifo_push = 1'h0;
		outfifo_in_eos = 1'h0;
		data_to_fifo = 16'h0000;
		infifo_pop[0] = 1'h0;
		infifo_pop[1] = 1'h0;
		if ((&infifo_out_valid & ~outfifo_full) & ~dense_mode) begin
			if (~(&infifo_out_eos)) begin
				outfifo_push = 1'h1;
				outfifo_in_eos = 1'h0;
				data_to_fifo = pe_output;
				infifo_pop[0] = 1'h1;
				infifo_pop[1] = 1'h1;
			end
			else begin
				outfifo_push = 1'h1;
				outfifo_in_eos = 1'h1;
				data_to_fifo = infifo_out_data[0+:16];
				infifo_pop[0] = 1'h1;
				infifo_pop[1] = 1'h1;
			end
		end
	end
	reg_fifo_depth_0_w_17_afd_2 input_fifo_0(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(infifo_in_packed[0+:17]),
		.flush(flush),
		.pop(infifo_pop[0]),
		.push(infifo_push_0),
		.rst_n(rst_n),
		.data_out(input_fifo_0_data_out),
		.empty(input_fifo_0_empty),
		.full(input_fifo_0_full)
	);
	reg_fifo_depth_0_w_17_afd_2 input_fifo_1(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(infifo_in_packed[17+:17]),
		.flush(flush),
		.pop(infifo_pop[1]),
		.push(infifo_push_1),
		.rst_n(rst_n),
		.data_out(input_fifo_1_data_out),
		.empty(input_fifo_1_empty),
		.full(input_fifo_1_full)
	);
	reg_fifo_depth_2_w_17_afd_2 output_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(outfifo_in_packed),
		.flush(flush),
		.pop(outfifo_pop),
		.push(outfifo_push),
		.rst_n(rst_n),
		.data_out(outfifo_out_packed),
		.empty(output_fifo_empty),
		.full(outfifo_full)
	);
	PEGEN_PE onyxpeintf(
		.ASYNCRESET(onyxpeintf_ASYNCRESET),
		.CLK(gclk),
		.bit0(bit0),
		.bit1(bit1),
		.bit2(bit2),
		.clk_en(clk_en),
		.data0(onyxpeintf_data0),
		.data1(onyxpeintf_data1),
		.data2(data2[15:0]),
		.inst(onyxpeintf_inst),
		.O0(pe_output),
		.O1(res_p),
		.O2(onyxpeintf_O2),
		.O3(onyxpeintf_O3),
		.O4(onyxpeintf_O4)
	);
endmodule
module PE_onyx_flat (
	PE_onyx_inst_dense_mode,
	PE_onyx_inst_onyxpeintf_inst,
	PE_onyx_inst_tile_en,
	bit0_f_,
	bit1_f_,
	bit2_f_,
	clk,
	clk_en,
	data0_f_,
	data0_valid_f_,
	data1_f_,
	data1_valid_f_,
	data2_f_,
	flush,
	res_ready_f_,
	rst_n,
	PE_onyx_inst_onyxpeintf_O2,
	PE_onyx_inst_onyxpeintf_O3,
	PE_onyx_inst_onyxpeintf_O4,
	data0_ready_f_,
	data1_ready_f_,
	res_f_,
	res_p_f_,
	res_valid_f_
);
	input wire PE_onyx_inst_dense_mode;
	input wire [83:0] PE_onyx_inst_onyxpeintf_inst;
	input wire PE_onyx_inst_tile_en;
	input wire bit0_f_;
	input wire bit1_f_;
	input wire bit2_f_;
	input wire clk;
	input wire clk_en;
	input wire [16:0] data0_f_;
	input wire data0_valid_f_;
	input wire [16:0] data1_f_;
	input wire data1_valid_f_;
	input wire [16:0] data2_f_;
	input wire flush;
	input wire res_ready_f_;
	input wire rst_n;
	output wire [15:0] PE_onyx_inst_onyxpeintf_O2;
	output wire [15:0] PE_onyx_inst_onyxpeintf_O3;
	output wire [15:0] PE_onyx_inst_onyxpeintf_O4;
	output wire data0_ready_f_;
	output wire data1_ready_f_;
	output wire [16:0] res_f_;
	output wire res_p_f_;
	output wire res_valid_f_;
	PE_onyx PE_onyx_inst(
		.bit0(bit0_f_),
		.bit1(bit1_f_),
		.bit2(bit2_f_),
		.clk(clk),
		.clk_en(clk_en),
		.data0(data0_f_),
		.data0_valid(data0_valid_f_),
		.data1(data1_f_),
		.data1_valid(data1_valid_f_),
		.data2(data2_f_),
		.dense_mode(PE_onyx_inst_dense_mode),
		.flush(flush),
		.onyxpeintf_inst(PE_onyx_inst_onyxpeintf_inst),
		.res_ready(res_ready_f_),
		.rst_n(rst_n),
		.tile_en(PE_onyx_inst_tile_en),
		.data0_ready(data0_ready_f_),
		.data1_ready(data1_ready_f_),
		.onyxpeintf_O2(PE_onyx_inst_onyxpeintf_O2),
		.onyxpeintf_O3(PE_onyx_inst_onyxpeintf_O3),
		.onyxpeintf_O4(PE_onyx_inst_onyxpeintf_O4),
		.res(res_f_),
		.res_p(res_p_f_),
		.res_valid(res_valid_f_)
	);
endmodule
module Repeat (
	clk,
	clk_en,
	flush,
	proc_data_in,
	proc_data_in_valid,
	ref_data_out_ready,
	repsig_data_in,
	repsig_data_in_valid,
	root,
	rst_n,
	spacc_mode,
	stop_lvl,
	tile_en,
	proc_data_in_ready,
	ref_data_out,
	ref_data_out_valid,
	repsig_data_in_ready
);
	input wire clk;
	input wire clk_en;
	input wire flush;
	input wire [16:0] proc_data_in;
	input wire proc_data_in_valid;
	input wire ref_data_out_ready;
	input wire [16:0] repsig_data_in;
	input wire repsig_data_in_valid;
	input wire root;
	input wire rst_n;
	input wire spacc_mode;
	input wire [15:0] stop_lvl;
	input wire tile_en;
	output wire proc_data_in_ready;
	output wire [16:0] ref_data_out;
	output wire ref_data_out_valid;
	output wire repsig_data_in_ready;
	wire clr_last_pushed_data;
	wire gclk;
	wire proc_done;
	wire proc_fifo_full;
	reg [15:0] proc_fifo_inject_data;
	reg proc_fifo_inject_eos;
	reg proc_fifo_inject_push;
	wire [15:0] proc_fifo_out_data;
	wire proc_fifo_out_eos;
	reg proc_fifo_pop;
	wire proc_fifo_push;
	wire proc_fifo_valid;
	wire [16:0] proc_in_fifo_data_in;
	wire [16:0] proc_in_fifo_data_out;
	wire proc_in_fifo_empty;
	wire proc_in_fifo_full;
	wire proc_stop;
	wire ref_fifo_full;
	reg [15:0] ref_fifo_in_data;
	reg ref_fifo_in_eos;
	reg ref_fifo_push;
	wire ref_maybe;
	wire [16:0] ref_out_fifo_data_in;
	wire ref_out_fifo_empty;
	reg [2:0] repeat_fsm_current_state;
	reg [2:0] repeat_fsm_next_state;
	wire repsig_done;
	wire [15:0] repsig_fifo_out_data;
	wire repsig_fifo_out_eos;
	reg repsig_fifo_pop;
	wire repsig_fifo_valid;
	wire [16:0] repsig_in_fifo_data_out;
	wire repsig_in_fifo_empty;
	wire repsig_in_fifo_full;
	wire repsig_stop;
	wire seen_root_eos_sticky;
	reg seen_root_eos_was_high;
	wire set_last_pushed_data;
	wire set_last_pushed_data_sticky;
	reg set_last_pushed_data_was_high;
	assign gclk = clk & tile_en;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			set_last_pushed_data_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				set_last_pushed_data_was_high <= 1'h0;
			else if (clr_last_pushed_data)
				set_last_pushed_data_was_high <= 1'h0;
			else if (set_last_pushed_data)
				set_last_pushed_data_was_high <= 1'h1;
		end
	assign set_last_pushed_data_sticky = set_last_pushed_data_was_high;
	assign {repsig_fifo_out_eos, repsig_fifo_out_data} = repsig_in_fifo_data_out;
	assign repsig_data_in_ready = ~repsig_in_fifo_full;
	assign repsig_fifo_valid = ~repsig_in_fifo_empty;
	assign proc_fifo_push = (root ? proc_fifo_inject_push : proc_data_in_valid);
	assign proc_in_fifo_data_in = (root ? {proc_fifo_inject_eos, proc_fifo_inject_data} : proc_data_in);
	assign {proc_fifo_out_eos, proc_fifo_out_data} = proc_in_fifo_data_out;
	assign proc_data_in_ready = ~proc_in_fifo_full;
	assign proc_fifo_full = proc_in_fifo_full;
	assign proc_fifo_valid = ~proc_in_fifo_empty;
	assign ref_out_fifo_data_in = {ref_fifo_in_eos, ref_fifo_in_data};
	assign ref_data_out_valid = ~ref_out_fifo_empty;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			seen_root_eos_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				seen_root_eos_was_high <= 1'h0;
			else if (((proc_fifo_out_data == 16'h0000) & proc_fifo_out_eos) & proc_fifo_valid)
				seen_root_eos_was_high <= 1'h1;
		end
	assign seen_root_eos_sticky = (((proc_fifo_out_data == 16'h0000) & proc_fifo_out_eos) & proc_fifo_valid) | seen_root_eos_was_high;
	assign proc_stop = ((proc_fifo_out_data[9:8] == 2'h0) & proc_fifo_out_eos) & proc_fifo_valid;
	assign proc_done = ((proc_fifo_out_data[9:8] == 2'h1) & proc_fifo_out_eos) & proc_fifo_valid;
	assign repsig_stop = ((repsig_fifo_out_data[9:8] == 2'h0) & repsig_fifo_out_eos) & repsig_fifo_valid;
	assign repsig_done = ((repsig_fifo_out_data[9:8] == 2'h1) & repsig_fifo_out_eos) & repsig_fifo_valid;
	assign ref_maybe = (proc_fifo_valid & proc_fifo_out_eos) & (proc_fifo_out_data[9:8] == 2'h2);
	always @(posedge clk or negedge rst_n)
		if (!rst_n)
			repeat_fsm_current_state <= 3'h5;
		else if (clk_en) begin
			if (flush)
				repeat_fsm_current_state <= 3'h5;
			else
				repeat_fsm_current_state <= repeat_fsm_next_state;
		end
	always @(*) begin
		repeat_fsm_next_state = repeat_fsm_current_state;
		case (repeat_fsm_current_state)
			3'h0:
				if ((~ref_fifo_full & proc_done) & repsig_done)
					repeat_fsm_next_state = 3'h5;
			3'h1:
				if (~proc_fifo_full)
					repeat_fsm_next_state = 3'h2;
				else
					repeat_fsm_next_state = 3'h1;
			3'h2:
				if (~proc_fifo_full)
					repeat_fsm_next_state = 3'h3;
				else
					repeat_fsm_next_state = 3'h2;
			3'h3:
				if (proc_done)
					repeat_fsm_next_state = 3'h0;
				else if ((repsig_fifo_out_eos & repsig_fifo_valid) & (repsig_fifo_out_data[9:8] == 2'h0))
					repeat_fsm_next_state = 3'h4;
				else
					repeat_fsm_next_state = 3'h3;
			3'h4:
				if ((proc_fifo_valid & ~proc_stop) & ~ref_fifo_full)
					repeat_fsm_next_state = 3'h3;
				else
					repeat_fsm_next_state = 3'h4;
			3'h5:
				if (root & tile_en)
					repeat_fsm_next_state = 3'h1;
				else if (~root & tile_en)
					repeat_fsm_next_state = 3'h3;
				else
					repeat_fsm_next_state = 3'h5;
			default: repeat_fsm_next_state = repeat_fsm_current_state;
		endcase
	end
	always @(*)
		case (repeat_fsm_current_state)
			3'h0: begin : repeat_fsm_DONE_Output
				ref_fifo_in_data = proc_fifo_out_data;
				ref_fifo_in_eos = 1'h1;
				ref_fifo_push = (~ref_fifo_full & proc_done) & repsig_done;
				proc_fifo_pop = (~ref_fifo_full & proc_done) & repsig_done;
				repsig_fifo_pop = (~ref_fifo_full & proc_done) & repsig_done;
				proc_fifo_inject_push = 1'h0;
				proc_fifo_inject_data = 16'h0000;
				proc_fifo_inject_eos = 1'h0;
			end
			3'h1: begin : repeat_fsm_INJECT0_Output
				ref_fifo_in_data = 16'h0000;
				ref_fifo_in_eos = 1'h0;
				ref_fifo_push = 1'h0;
				proc_fifo_pop = 1'h0;
				repsig_fifo_pop = 1'h0;
				proc_fifo_inject_push = 1'h1;
				proc_fifo_inject_data = 16'h0000;
				proc_fifo_inject_eos = 1'h0;
			end
			3'h2: begin : repeat_fsm_INJECT1_Output
				ref_fifo_in_data = 16'h0000;
				ref_fifo_in_eos = 1'h0;
				ref_fifo_push = 1'h0;
				proc_fifo_pop = 1'h0;
				repsig_fifo_pop = 1'h0;
				proc_fifo_inject_push = 1'h1;
				proc_fifo_inject_data = 16'h0100;
				proc_fifo_inject_eos = 1'h1;
			end
			3'h3: begin : repeat_fsm_PASS_REPEAT_Output
				ref_fifo_in_data = proc_fifo_out_data;
				ref_fifo_in_eos = ref_maybe;
				ref_fifo_push = (((repsig_fifo_valid & proc_fifo_valid) & ~repsig_fifo_out_eos) & ~proc_done) & ~ref_fifo_full;
				proc_fifo_pop = (((repsig_fifo_valid & repsig_fifo_out_eos) & ~spacc_mode) | (spacc_mode & repsig_done)) & ~proc_done;
				repsig_fifo_pop = (((~ref_fifo_full & repsig_fifo_valid) & ~repsig_fifo_out_eos) & proc_fifo_valid) & ~proc_done;
				proc_fifo_inject_push = 1'h0;
				proc_fifo_inject_data = 16'h0000;
				proc_fifo_inject_eos = 1'h0;
			end
			3'h4: begin : repeat_fsm_PASS_STOP_Output
				ref_fifo_in_data = repsig_fifo_out_data;
				ref_fifo_in_eos = 1'h1;
				ref_fifo_push = (repsig_stop & proc_fifo_valid) & ~ref_fifo_full;
				proc_fifo_pop = (repsig_fifo_valid & proc_stop) & ~ref_fifo_full;
				repsig_fifo_pop = (repsig_stop & proc_fifo_valid) & ~ref_fifo_full;
				proc_fifo_inject_push = 1'h0;
				proc_fifo_inject_data = 16'h0000;
				proc_fifo_inject_eos = 1'h0;
			end
			3'h5: begin : repeat_fsm_START_Output
				ref_fifo_in_data = 16'h0000;
				ref_fifo_in_eos = 1'h0;
				ref_fifo_push = 1'h0;
				proc_fifo_pop = 1'h0;
				repsig_fifo_pop = 1'h0;
				proc_fifo_inject_push = 1'h0;
				proc_fifo_inject_data = 16'h0000;
				proc_fifo_inject_eos = 1'h0;
			end
			default: begin : repeat_fsm_default_Output
				ref_fifo_in_data = 16'h0000;
				ref_fifo_in_eos = 1'h0;
				ref_fifo_push = 1'h0;
				proc_fifo_pop = 1'h0;
				repsig_fifo_pop = 1'h0;
				proc_fifo_inject_push = 1'h0;
				proc_fifo_inject_data = 16'h0000;
				proc_fifo_inject_eos = 1'h0;
			end
		endcase
	reg_fifo_depth_0_w_17_afd_2 repsig_in_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(repsig_data_in),
		.flush(flush),
		.pop(repsig_fifo_pop),
		.push(repsig_data_in_valid),
		.rst_n(rst_n),
		.data_out(repsig_in_fifo_data_out),
		.empty(repsig_in_fifo_empty),
		.full(repsig_in_fifo_full)
	);
	reg_fifo_depth_2_w_17_afd_2 proc_in_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(proc_in_fifo_data_in),
		.flush(flush),
		.pop(proc_fifo_pop),
		.push(proc_fifo_push),
		.rst_n(rst_n),
		.data_out(proc_in_fifo_data_out),
		.empty(proc_in_fifo_empty),
		.full(proc_in_fifo_full)
	);
	reg_fifo_depth_0_w_17_afd_2 ref_out_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(ref_out_fifo_data_in),
		.flush(flush),
		.pop(ref_data_out_ready),
		.push(ref_fifo_push),
		.rst_n(rst_n),
		.data_out(ref_data_out),
		.empty(ref_out_fifo_empty),
		.full(ref_fifo_full)
	);
endmodule
module RepeatSignalGenerator (
	base_data_in,
	base_data_in_valid,
	clk,
	clk_en,
	flush,
	repsig_data_out_ready,
	rst_n,
	stop_lvl,
	tile_en,
	base_data_in_ready,
	repsig_data_out,
	repsig_data_out_valid
);
	input wire [16:0] base_data_in;
	input wire base_data_in_valid;
	input wire clk;
	input wire clk_en;
	input wire flush;
	input wire repsig_data_out_ready;
	input wire rst_n;
	input wire [15:0] stop_lvl;
	input wire tile_en;
	output wire base_data_in_ready;
	output wire [16:0] repsig_data_out;
	output wire repsig_data_out_valid;
	wire already_pushed_repsig_eos_sticky;
	reg already_pushed_repsig_eos_was_high;
	wire [15:0] base_fifo_out_data;
	wire base_fifo_out_eos;
	reg base_fifo_pop;
	wire base_fifo_valid;
	wire [16:0] base_in_fifo_data_out;
	wire base_in_fifo_empty;
	wire base_in_fifo_full;
	reg clr_already_pushed_repsig_eos;
	wire gclk;
	wire repsig_fifo_full;
	reg [15:0] repsig_fifo_in_data;
	reg repsig_fifo_in_eos;
	reg repsig_fifo_push;
	wire [16:0] repsig_out_fifo_data_in;
	wire repsig_out_fifo_empty;
	reg [1:0] rsg_fsm_current_state;
	reg [1:0] rsg_fsm_next_state;
	wire seen_root_eos_sticky;
	reg seen_root_eos_was_high;
	assign gclk = clk & tile_en;
	assign {base_fifo_out_eos, base_fifo_out_data} = base_in_fifo_data_out;
	assign base_data_in_ready = ~base_in_fifo_full;
	assign base_fifo_valid = ~base_in_fifo_empty;
	assign repsig_out_fifo_data_in = {repsig_fifo_in_eos, repsig_fifo_in_data};
	assign repsig_data_out_valid = ~repsig_out_fifo_empty;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			seen_root_eos_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				seen_root_eos_was_high <= 1'h0;
			else if (((base_fifo_out_data[9:8] == 2'h1) & base_fifo_out_eos) & base_fifo_valid)
				seen_root_eos_was_high <= 1'h1;
		end
	assign seen_root_eos_sticky = (((base_fifo_out_data[9:8] == 2'h1) & base_fifo_out_eos) & base_fifo_valid) | seen_root_eos_was_high;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			already_pushed_repsig_eos_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				already_pushed_repsig_eos_was_high <= 1'h0;
			else if (clr_already_pushed_repsig_eos)
				already_pushed_repsig_eos_was_high <= 1'h0;
			else if (repsig_fifo_push & ~repsig_fifo_full)
				already_pushed_repsig_eos_was_high <= 1'h1;
		end
	assign already_pushed_repsig_eos_sticky = already_pushed_repsig_eos_was_high;
	always @(posedge clk or negedge rst_n)
		if (!rst_n)
			rsg_fsm_current_state <= 2'h3;
		else if (clk_en) begin
			if (flush)
				rsg_fsm_current_state <= 2'h3;
			else
				rsg_fsm_current_state <= rsg_fsm_next_state;
		end
	always @(*) begin
		rsg_fsm_next_state = rsg_fsm_current_state;
		case (rsg_fsm_current_state)
			2'h0: rsg_fsm_next_state = 2'h3;
			2'h1:
				if (base_fifo_out_eos & base_fifo_valid)
					rsg_fsm_next_state = 2'h2;
				else
					rsg_fsm_next_state = 2'h1;
			2'h2:
				if (((base_fifo_valid & base_fifo_out_eos) & (base_fifo_out_data[9:8] == 2'h1)) & ~repsig_fifo_full)
					rsg_fsm_next_state = 2'h0;
				else if (base_fifo_valid & ~base_fifo_out_eos)
					rsg_fsm_next_state = 2'h1;
				else
					rsg_fsm_next_state = 2'h2;
			2'h3:
				if (tile_en)
					rsg_fsm_next_state = 2'h1;
				else
					rsg_fsm_next_state = 2'h3;
			default:
				;
		endcase
	end
	always @(*)
		case (rsg_fsm_current_state)
			2'h0: begin : rsg_fsm_DONE_Output
				repsig_fifo_in_data = 16'h0000;
				repsig_fifo_in_eos = 1'h0;
				repsig_fifo_push = 1'h0;
				base_fifo_pop = 1'h0;
				clr_already_pushed_repsig_eos = 1'h0;
			end
			2'h1: begin : rsg_fsm_PASS_REPEAT_Output
				repsig_fifo_in_data = 16'h0001;
				repsig_fifo_in_eos = 1'h0;
				repsig_fifo_push = ~base_fifo_out_eos & base_fifo_valid;
				clr_already_pushed_repsig_eos = 1'h1;
				base_fifo_pop = (~base_fifo_out_eos & base_fifo_valid) & ~repsig_fifo_full;
			end
			2'h2: begin : rsg_fsm_PASS_STOP_Output
				repsig_fifo_in_data = (base_fifo_out_data[9:8] == 2'h1 ? base_fifo_out_data : base_fifo_out_data);
				repsig_fifo_in_eos = 1'h1;
				repsig_fifo_push = base_fifo_out_eos & base_fifo_valid;
				clr_already_pushed_repsig_eos = 1'h0;
				base_fifo_pop = (base_fifo_out_eos & base_fifo_valid) & ~repsig_fifo_full;
			end
			2'h3: begin : rsg_fsm_START_Output
				repsig_fifo_in_data = 16'h0000;
				repsig_fifo_in_eos = 1'h0;
				repsig_fifo_push = 1'h0;
				base_fifo_pop = 1'h0;
				clr_already_pushed_repsig_eos = 1'h0;
			end
			default:
				;
		endcase
	reg_fifo_depth_0_w_17_afd_2 base_in_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(base_data_in),
		.flush(flush),
		.pop(base_fifo_pop),
		.push(base_data_in_valid),
		.rst_n(rst_n),
		.data_out(base_in_fifo_data_out),
		.empty(base_in_fifo_empty),
		.full(base_in_fifo_full)
	);
	reg_fifo_depth_0_w_17_afd_2 repsig_out_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(repsig_out_fifo_data_in),
		.flush(flush),
		.pop(repsig_data_out_ready),
		.push(repsig_fifo_push),
		.rst_n(rst_n),
		.data_out(repsig_data_out),
		.empty(repsig_out_fifo_empty),
		.full(repsig_fifo_full)
	);
endmodule
module RepeatSignalGenerator_flat (
	RepeatSignalGenerator_inst_stop_lvl,
	RepeatSignalGenerator_inst_tile_en,
	base_data_in_f_,
	base_data_in_valid_f_,
	clk,
	clk_en,
	flush,
	repsig_data_out_ready_f_,
	rst_n,
	base_data_in_ready_f_,
	repsig_data_out_f_,
	repsig_data_out_valid_f_
);
	input wire [15:0] RepeatSignalGenerator_inst_stop_lvl;
	input wire RepeatSignalGenerator_inst_tile_en;
	input wire [16:0] base_data_in_f_;
	input wire base_data_in_valid_f_;
	input wire clk;
	input wire clk_en;
	input wire flush;
	input wire repsig_data_out_ready_f_;
	input wire rst_n;
	output wire base_data_in_ready_f_;
	output wire [16:0] repsig_data_out_f_;
	output wire repsig_data_out_valid_f_;
	RepeatSignalGenerator RepeatSignalGenerator_inst(
		.base_data_in(base_data_in_f_),
		.base_data_in_valid(base_data_in_valid_f_),
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.repsig_data_out_ready(repsig_data_out_ready_f_),
		.rst_n(rst_n),
		.stop_lvl(RepeatSignalGenerator_inst_stop_lvl),
		.tile_en(RepeatSignalGenerator_inst_tile_en),
		.base_data_in_ready(base_data_in_ready_f_),
		.repsig_data_out(repsig_data_out_f_),
		.repsig_data_out_valid(repsig_data_out_valid_f_)
	);
endmodule
module Repeat_flat (
	Repeat_inst_root,
	Repeat_inst_spacc_mode,
	Repeat_inst_stop_lvl,
	Repeat_inst_tile_en,
	clk,
	clk_en,
	flush,
	proc_data_in_f_,
	proc_data_in_valid_f_,
	ref_data_out_ready_f_,
	repsig_data_in_f_,
	repsig_data_in_valid_f_,
	rst_n,
	proc_data_in_ready_f_,
	ref_data_out_f_,
	ref_data_out_valid_f_,
	repsig_data_in_ready_f_
);
	input wire Repeat_inst_root;
	input wire Repeat_inst_spacc_mode;
	input wire [15:0] Repeat_inst_stop_lvl;
	input wire Repeat_inst_tile_en;
	input wire clk;
	input wire clk_en;
	input wire flush;
	input wire [16:0] proc_data_in_f_;
	input wire proc_data_in_valid_f_;
	input wire ref_data_out_ready_f_;
	input wire [16:0] repsig_data_in_f_;
	input wire repsig_data_in_valid_f_;
	input wire rst_n;
	output wire proc_data_in_ready_f_;
	output wire [16:0] ref_data_out_f_;
	output wire ref_data_out_valid_f_;
	output wire repsig_data_in_ready_f_;
	Repeat Repeat_inst(
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.proc_data_in(proc_data_in_f_),
		.proc_data_in_valid(proc_data_in_valid_f_),
		.ref_data_out_ready(ref_data_out_ready_f_),
		.repsig_data_in(repsig_data_in_f_),
		.repsig_data_in_valid(repsig_data_in_valid_f_),
		.root(Repeat_inst_root),
		.rst_n(rst_n),
		.spacc_mode(Repeat_inst_spacc_mode),
		.stop_lvl(Repeat_inst_stop_lvl),
		.tile_en(Repeat_inst_tile_en),
		.proc_data_in_ready(proc_data_in_ready_f_),
		.ref_data_out(ref_data_out_f_),
		.ref_data_out_valid(ref_data_out_valid_f_),
		.repsig_data_in_ready(repsig_data_in_ready_f_)
	);
endmodule
module crddrop (
	clk,
	clk_en,
	cmrg_coord_in_0,
	cmrg_coord_in_0_valid,
	cmrg_coord_in_1,
	cmrg_coord_in_1_valid,
	cmrg_coord_out_0_ready,
	cmrg_coord_out_1_ready,
	cmrg_enable,
	cmrg_stop_lvl,
	flush,
	rst_n,
	tile_en,
	cmrg_coord_in_0_ready,
	cmrg_coord_in_1_ready,
	cmrg_coord_out_0,
	cmrg_coord_out_0_valid,
	cmrg_coord_out_1,
	cmrg_coord_out_1_valid
);
	input wire clk;
	input wire clk_en;
	input wire [16:0] cmrg_coord_in_0;
	input wire cmrg_coord_in_0_valid;
	input wire [16:0] cmrg_coord_in_1;
	input wire cmrg_coord_in_1_valid;
	input wire cmrg_coord_out_0_ready;
	input wire cmrg_coord_out_1_ready;
	input wire cmrg_enable;
	input wire [15:0] cmrg_stop_lvl;
	input wire flush;
	input wire rst_n;
	input wire tile_en;
	output wire cmrg_coord_in_0_ready;
	output wire cmrg_coord_in_1_ready;
	output wire [16:0] cmrg_coord_out_0;
	output wire cmrg_coord_out_0_valid;
	output wire [16:0] cmrg_coord_out_1;
	output wire cmrg_coord_out_1_valid;
	wire base_data_seen;
	wire base_done;
	wire base_done_seen;
	wire base_eos_seen;
	wire base_infifo_empty;
	wire base_infifo_full;
	wire [15:0] base_infifo_in_data;
	wire base_infifo_in_eos;
	wire [16:0] base_infifo_in_packed;
	wire base_infifo_in_valid;
	wire [16:0] base_infifo_out_packed;
	wire base_outfifo_empty;
	wire base_outfifo_full;
	wire [16:0] base_outfifo_in_packed;
	wire [16:0] base_outfifo_out_packed;
	wire both_done;
	reg clr_pushed_data_lower;
	reg clr_pushed_proc;
	reg clr_pushed_stop_lvl;
	wire cmrg_coord_in_0_eos;
	wire cmrg_coord_in_1_eos;
	reg [1:0] cmrg_fifo_pop;
	reg [1:0] cmrg_fifo_push;
	wire gclk;
	wire proc_data_seen;
	wire proc_done;
	wire proc_infifo_empty;
	wire proc_infifo_full;
	wire [15:0] proc_infifo_in_data;
	wire proc_infifo_in_eos;
	wire [16:0] proc_infifo_in_packed;
	wire proc_infifo_in_valid;
	wire [16:0] proc_infifo_out_packed;
	wire proc_outfifo_empty;
	wire proc_outfifo_full;
	wire [16:0] proc_outfifo_in_packed;
	wire [16:0] proc_outfifo_out_packed;
	reg proc_seq_current_state;
	reg proc_seq_next_state;
	wire pushed_data_sticky_sticky;
	reg pushed_data_sticky_was_high;
	wire pushed_proc_sticky;
	reg pushed_proc_was_high;
	wire pushed_stop_lvl_sticky;
	reg pushed_stop_lvl_was_high;
	wire pushing_done;
	reg set_pushed_data_lower;
	assign gclk = clk & tile_en;
	assign cmrg_coord_in_0_eos = cmrg_coord_in_0[16];
	assign cmrg_coord_in_1_eos = cmrg_coord_in_1[16];
	assign base_infifo_in_packed[16] = cmrg_coord_in_0_eos;
	assign base_infifo_in_packed[15:0] = cmrg_coord_in_0[15:0];
	assign base_infifo_in_eos = base_infifo_out_packed[16];
	assign base_infifo_in_data = base_infifo_out_packed[15:0];
	assign base_infifo_in_valid = ~base_infifo_empty;
	assign cmrg_coord_in_0_ready = ~base_infifo_full;
	assign proc_infifo_in_packed[16] = cmrg_coord_in_1_eos;
	assign proc_infifo_in_packed[15:0] = cmrg_coord_in_1[15:0];
	assign proc_infifo_in_eos = proc_infifo_out_packed[16];
	assign proc_infifo_in_data = proc_infifo_out_packed[15:0];
	assign proc_infifo_in_valid = ~proc_infifo_empty;
	assign cmrg_coord_in_1_ready = ~proc_infifo_full;
	assign base_data_seen = base_infifo_in_valid & ~base_infifo_in_eos;
	assign proc_data_seen = proc_infifo_in_valid & ~proc_infifo_in_eos;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			pushed_data_sticky_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				pushed_data_sticky_was_high <= 1'h0;
			else if (clr_pushed_data_lower)
				pushed_data_sticky_was_high <= 1'h0;
			else if (set_pushed_data_lower)
				pushed_data_sticky_was_high <= 1'h1;
		end
	assign pushed_data_sticky_sticky = pushed_data_sticky_was_high;
	assign base_eos_seen = (base_infifo_in_valid & base_infifo_in_eos) & (base_infifo_in_data[9:8] == 2'h0);
	assign base_done_seen = (base_infifo_in_valid & base_infifo_in_eos) & (base_infifo_in_data[9:8] == 2'h1);
	assign base_done = (base_infifo_in_valid & base_infifo_in_eos) & (base_infifo_in_data[9:8] == 2'h1);
	assign proc_done = (proc_infifo_in_valid & proc_infifo_in_eos) & (proc_infifo_in_data[9:8] == 2'h1);
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			pushed_proc_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				pushed_proc_was_high <= 1'h0;
			else if (clr_pushed_proc)
				pushed_proc_was_high <= 1'h0;
			else if (cmrg_fifo_push[1])
				pushed_proc_was_high <= 1'h1;
		end
	assign pushed_proc_sticky = pushed_proc_was_high;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			pushed_stop_lvl_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				pushed_stop_lvl_was_high <= 1'h0;
			else if (clr_pushed_stop_lvl)
				pushed_stop_lvl_was_high <= 1'h0;
			else if ((cmrg_fifo_push[0] & base_infifo_in_valid) & base_infifo_in_eos)
				pushed_stop_lvl_was_high <= 1'h1;
		end
	assign pushed_stop_lvl_sticky = pushed_stop_lvl_was_high;
	assign both_done = ((((base_infifo_in_valid & base_infifo_in_eos) & proc_infifo_in_valid) & proc_infifo_in_eos) & (base_infifo_in_data[9:8] == 2'h1)) & (proc_infifo_in_data[9:8] == 2'h1);
	assign pushing_done = ((((((base_infifo_in_valid & base_infifo_in_eos) & proc_infifo_in_valid) & proc_infifo_in_eos) & (base_infifo_in_data[9:8] == 2'h1)) & (proc_infifo_in_data[9:8] == 2'h1)) & ~base_outfifo_full) & ~proc_outfifo_full;
	assign base_outfifo_in_packed[16] = base_infifo_in_eos;
	assign base_outfifo_in_packed[15:0] = base_infifo_in_data;
	assign cmrg_coord_out_0[16] = base_outfifo_out_packed[16];
	assign cmrg_coord_out_0[15:0] = base_outfifo_out_packed[15:0];
	assign cmrg_coord_out_0_valid = ~base_outfifo_empty;
	assign proc_outfifo_in_packed[16] = proc_infifo_in_eos;
	assign proc_outfifo_in_packed[15:0] = proc_infifo_in_data;
	assign cmrg_coord_out_1[16] = proc_outfifo_out_packed[16];
	assign cmrg_coord_out_1[15:0] = proc_outfifo_out_packed[15:0];
	assign cmrg_coord_out_1_valid = ~proc_outfifo_empty;
	always @(posedge clk or negedge rst_n)
		if (!rst_n)
			proc_seq_current_state <= 1'h1;
		else if (clk_en) begin
			if (flush)
				proc_seq_current_state <= 1'h1;
			else
				proc_seq_current_state <= proc_seq_next_state;
		end
	always @(*) begin
		proc_seq_next_state = proc_seq_current_state;
		case (proc_seq_current_state)
			1'h0: proc_seq_next_state = 1'h0;
			1'h1:
				if (tile_en)
					proc_seq_next_state = 1'h0;
				else
					proc_seq_next_state = 1'h1;
			default:
				;
		endcase
	end
	always @(*)
		case (proc_seq_current_state)
			1'h0: begin : proc_seq_PROCESS_Output
				cmrg_fifo_pop[0] = (base_done ? (proc_done & ~base_outfifo_full) & ~proc_outfifo_full : (base_infifo_in_valid & ~base_infifo_in_eos ? ~base_outfifo_full : (base_infifo_in_valid & base_infifo_in_eos ? ((proc_done | (proc_infifo_in_valid & ~proc_infifo_in_eos)) & ~base_outfifo_full) & ~proc_outfifo_full : 1'h0)));
				cmrg_fifo_pop[1] = (proc_done ? (base_done & ~base_outfifo_full) & ~proc_outfifo_full : (((base_infifo_in_valid & base_infifo_in_eos) & proc_infifo_in_valid) & ~proc_infifo_in_eos ? ~base_outfifo_full & (~proc_outfifo_full | ~pushed_data_sticky_sticky) : (proc_infifo_in_valid & proc_infifo_in_eos ? ~proc_outfifo_full : 1'h0)));
				cmrg_fifo_push[0] = (base_done ? proc_done : (base_infifo_in_valid & ~base_infifo_in_eos ? ~base_outfifo_full : (base_infifo_in_valid & base_infifo_in_eos ? ((proc_done | ((proc_infifo_in_valid & ~proc_infifo_in_eos) & pushed_data_sticky_sticky)) & ~base_outfifo_full) & ~proc_outfifo_full : 1'h0)));
				cmrg_fifo_push[1] = (proc_done ? base_done : (((base_infifo_in_valid & base_infifo_in_eos) & proc_infifo_in_valid) & ~proc_infifo_in_eos ? (~base_outfifo_full & ~proc_outfifo_full) & pushed_data_sticky_sticky : (proc_infifo_in_valid & proc_infifo_in_eos ? ~proc_outfifo_full : 1'h0)));
				clr_pushed_proc = 1'h0;
				clr_pushed_stop_lvl = 1'h0;
				set_pushed_data_lower = (base_infifo_in_valid & ~base_infifo_in_eos) & ~base_outfifo_full;
				clr_pushed_data_lower = base_done | (((((base_infifo_in_valid & base_infifo_in_eos) & proc_infifo_in_valid) & ~proc_infifo_in_eos) & ~base_outfifo_full) & ~proc_outfifo_full);
			end
			1'h1: begin : proc_seq_START_Output
				cmrg_fifo_pop[0] = 1'h0;
				cmrg_fifo_pop[1] = 1'h0;
				cmrg_fifo_push[0] = 1'h0;
				cmrg_fifo_push[1] = 1'h0;
				clr_pushed_proc = 1'h1;
				clr_pushed_stop_lvl = 1'h1;
				set_pushed_data_lower = 1'h0;
				clr_pushed_data_lower = 1'h1;
			end
			default:
				;
		endcase
	reg_fifo_depth_0_w_17_afd_2 base_infifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(base_infifo_in_packed),
		.flush(flush),
		.pop(cmrg_fifo_pop[0]),
		.push(cmrg_coord_in_0_valid),
		.rst_n(rst_n),
		.data_out(base_infifo_out_packed),
		.empty(base_infifo_empty),
		.full(base_infifo_full)
	);
	reg_fifo_depth_0_w_17_afd_2 proc_infifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(proc_infifo_in_packed),
		.flush(flush),
		.pop(cmrg_fifo_pop[1]),
		.push(cmrg_coord_in_1_valid),
		.rst_n(rst_n),
		.data_out(proc_infifo_out_packed),
		.empty(proc_infifo_empty),
		.full(proc_infifo_full)
	);
	reg_fifo_depth_0_w_17_afd_2 base_outfifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(base_outfifo_in_packed),
		.flush(flush),
		.pop(cmrg_coord_out_0_ready),
		.push(cmrg_fifo_push[0]),
		.rst_n(rst_n),
		.data_out(base_outfifo_out_packed),
		.empty(base_outfifo_empty),
		.full(base_outfifo_full)
	);
	reg_fifo_depth_0_w_17_afd_2 proc_outfifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(proc_outfifo_in_packed),
		.flush(flush),
		.pop(cmrg_coord_out_1_ready),
		.push(cmrg_fifo_push[1]),
		.rst_n(rst_n),
		.data_out(proc_outfifo_out_packed),
		.empty(proc_outfifo_empty),
		.full(proc_outfifo_full)
	);
endmodule
module crddrop_flat (
	clk,
	clk_en,
	cmrg_coord_in_0_f_,
	cmrg_coord_in_0_valid_f_,
	cmrg_coord_in_1_f_,
	cmrg_coord_in_1_valid_f_,
	cmrg_coord_out_0_ready_f_,
	cmrg_coord_out_1_ready_f_,
	crddrop_inst_cmrg_enable,
	crddrop_inst_cmrg_stop_lvl,
	crddrop_inst_tile_en,
	flush,
	rst_n,
	cmrg_coord_in_0_ready_f_,
	cmrg_coord_in_1_ready_f_,
	cmrg_coord_out_0_f_,
	cmrg_coord_out_0_valid_f_,
	cmrg_coord_out_1_f_,
	cmrg_coord_out_1_valid_f_
);
	input wire clk;
	input wire clk_en;
	input wire [16:0] cmrg_coord_in_0_f_;
	input wire cmrg_coord_in_0_valid_f_;
	input wire [16:0] cmrg_coord_in_1_f_;
	input wire cmrg_coord_in_1_valid_f_;
	input wire cmrg_coord_out_0_ready_f_;
	input wire cmrg_coord_out_1_ready_f_;
	input wire crddrop_inst_cmrg_enable;
	input wire [15:0] crddrop_inst_cmrg_stop_lvl;
	input wire crddrop_inst_tile_en;
	input wire flush;
	input wire rst_n;
	output wire cmrg_coord_in_0_ready_f_;
	output wire cmrg_coord_in_1_ready_f_;
	output wire [16:0] cmrg_coord_out_0_f_;
	output wire cmrg_coord_out_0_valid_f_;
	output wire [16:0] cmrg_coord_out_1_f_;
	output wire cmrg_coord_out_1_valid_f_;
	crddrop crddrop_inst(
		.clk(clk),
		.clk_en(clk_en),
		.cmrg_coord_in_0(cmrg_coord_in_0_f_),
		.cmrg_coord_in_0_valid(cmrg_coord_in_0_valid_f_),
		.cmrg_coord_in_1(cmrg_coord_in_1_f_),
		.cmrg_coord_in_1_valid(cmrg_coord_in_1_valid_f_),
		.cmrg_coord_out_0_ready(cmrg_coord_out_0_ready_f_),
		.cmrg_coord_out_1_ready(cmrg_coord_out_1_ready_f_),
		.cmrg_enable(crddrop_inst_cmrg_enable),
		.cmrg_stop_lvl(crddrop_inst_cmrg_stop_lvl),
		.flush(flush),
		.rst_n(rst_n),
		.tile_en(crddrop_inst_tile_en),
		.cmrg_coord_in_0_ready(cmrg_coord_in_0_ready_f_),
		.cmrg_coord_in_1_ready(cmrg_coord_in_1_ready_f_),
		.cmrg_coord_out_0(cmrg_coord_out_0_f_),
		.cmrg_coord_out_0_valid(cmrg_coord_out_0_valid_f_),
		.cmrg_coord_out_1(cmrg_coord_out_1_f_),
		.cmrg_coord_out_1_valid(cmrg_coord_out_1_valid_f_)
	);
endmodule
module crdhold (
	clk,
	clk_en,
	cmrg_coord_in_0,
	cmrg_coord_in_0_valid,
	cmrg_coord_in_1,
	cmrg_coord_in_1_valid,
	cmrg_coord_out_0_ready,
	cmrg_coord_out_1_ready,
	cmrg_enable,
	cmrg_stop_lvl,
	flush,
	rst_n,
	tile_en,
	cmrg_coord_in_0_ready,
	cmrg_coord_in_1_ready,
	cmrg_coord_out_0,
	cmrg_coord_out_0_valid,
	cmrg_coord_out_1,
	cmrg_coord_out_1_valid
);
	input wire clk;
	input wire clk_en;
	input wire [16:0] cmrg_coord_in_0;
	input wire cmrg_coord_in_0_valid;
	input wire [16:0] cmrg_coord_in_1;
	input wire cmrg_coord_in_1_valid;
	input wire cmrg_coord_out_0_ready;
	input wire cmrg_coord_out_1_ready;
	input wire cmrg_enable;
	input wire [15:0] cmrg_stop_lvl;
	input wire flush;
	input wire rst_n;
	input wire tile_en;
	output wire cmrg_coord_in_0_ready;
	output wire cmrg_coord_in_1_ready;
	output wire [16:0] cmrg_coord_out_0;
	output wire cmrg_coord_out_0_valid;
	output wire [16:0] cmrg_coord_out_1;
	output wire cmrg_coord_out_1_valid;
	wire base_data_seen;
	wire base_done_seen;
	wire base_eos_seen;
	wire base_infifo_empty;
	wire base_infifo_full;
	wire [15:0] base_infifo_in_data;
	wire base_infifo_in_eos;
	wire [16:0] base_infifo_in_packed;
	wire base_infifo_in_valid;
	wire [16:0] base_infifo_out_packed;
	wire base_outfifo_empty;
	wire base_outfifo_full;
	wire [16:0] base_outfifo_in_packed;
	wire [16:0] base_outfifo_out_packed;
	wire both_done;
	reg clr_pushed_base;
	reg clr_pushed_proc;
	wire cmrg_coord_in_0_eos;
	wire cmrg_coord_in_1_eos;
	reg [1:0] cmrg_fifo_pop;
	reg [1:0] cmrg_fifo_push;
	reg [15:0] data_to_fifo;
	reg eos_to_fifo;
	wire gclk;
	reg [15:0] hold_reg;
	wire proc_data_seen;
	wire proc_done_seen;
	wire proc_eos_seen;
	wire proc_infifo_empty;
	wire proc_infifo_full;
	wire [15:0] proc_infifo_in_data;
	wire proc_infifo_in_eos;
	wire [16:0] proc_infifo_in_packed;
	wire proc_infifo_in_valid;
	wire [16:0] proc_infifo_out_packed;
	wire proc_outfifo_empty;
	wire proc_outfifo_full;
	wire [16:0] proc_outfifo_in_packed;
	wire [16:0] proc_outfifo_out_packed;
	reg [1:0] proc_seq_current_state;
	reg [1:0] proc_seq_next_state;
	wire pushed_base_sticky;
	reg pushed_base_was_high;
	wire pushed_proc_sticky;
	reg pushed_proc_was_high;
	wire pushing_done;
	reg reg_clr;
	reg reg_hold;
	assign gclk = clk & tile_en;
	assign cmrg_coord_in_0_eos = cmrg_coord_in_0[16];
	assign cmrg_coord_in_1_eos = cmrg_coord_in_1[16];
	assign base_infifo_in_packed[16] = cmrg_coord_in_0_eos;
	assign base_infifo_in_packed[15:0] = cmrg_coord_in_0[15:0];
	assign base_infifo_in_eos = base_infifo_out_packed[16];
	assign base_infifo_in_data = base_infifo_out_packed[15:0];
	assign base_infifo_in_valid = ~base_infifo_empty;
	assign cmrg_coord_in_0_ready = ~base_infifo_full;
	assign proc_infifo_in_packed[16] = cmrg_coord_in_1_eos;
	assign proc_infifo_in_packed[15:0] = cmrg_coord_in_1[15:0];
	assign proc_infifo_in_eos = proc_infifo_out_packed[16];
	assign proc_infifo_in_data = proc_infifo_out_packed[15:0];
	assign proc_infifo_in_valid = ~proc_infifo_empty;
	assign cmrg_coord_in_1_ready = ~proc_infifo_full;
	assign base_data_seen = base_infifo_in_valid & ~base_infifo_in_eos;
	assign proc_data_seen = proc_infifo_in_valid & ~proc_infifo_in_eos;
	assign base_eos_seen = (base_infifo_in_valid & base_infifo_in_eos) & (base_infifo_in_data[9:8] == 2'h0);
	assign proc_eos_seen = (proc_infifo_in_valid & proc_infifo_in_eos) & (proc_infifo_in_data[9:8] == 2'h0);
	assign base_done_seen = (base_infifo_in_valid & base_infifo_in_eos) & (base_infifo_in_data[9:8] == 2'h1);
	assign proc_done_seen = (proc_infifo_in_valid & proc_infifo_in_eos) & (proc_infifo_in_data[9:8] == 2'h1);
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			pushed_proc_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				pushed_proc_was_high <= 1'h0;
			else if (clr_pushed_proc)
				pushed_proc_was_high <= 1'h0;
			else if (cmrg_fifo_push[1])
				pushed_proc_was_high <= 1'h1;
		end
	assign pushed_proc_sticky = pushed_proc_was_high;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			pushed_base_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				pushed_base_was_high <= 1'h0;
			else if (clr_pushed_base)
				pushed_base_was_high <= 1'h0;
			else if (cmrg_fifo_push[0])
				pushed_base_was_high <= 1'h1;
		end
	assign pushed_base_sticky = pushed_base_was_high;
	assign both_done = ((((base_infifo_in_valid & base_infifo_in_eos) & proc_infifo_in_valid) & proc_infifo_in_eos) & (base_infifo_in_data[9:8] == 2'h1)) & (proc_infifo_in_data[9:8] == 2'h1);
	assign pushing_done = ((((((base_infifo_in_valid & base_infifo_in_eos) & proc_infifo_in_valid) & proc_infifo_in_eos) & (base_infifo_in_data[9:8] == 2'h1)) & (proc_infifo_in_data[9:8] == 2'h1)) & ~base_outfifo_full) & ~proc_outfifo_full;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			hold_reg <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				hold_reg <= 16'h0000;
			else if (reg_clr)
				hold_reg <= 16'h0000;
			else if (reg_hold)
				hold_reg <= proc_infifo_in_data;
		end
	assign base_outfifo_in_packed[16] = base_infifo_in_eos;
	assign base_outfifo_in_packed[15:0] = base_infifo_in_data;
	assign cmrg_coord_out_0[16] = base_outfifo_out_packed[16];
	assign cmrg_coord_out_0[15:0] = base_outfifo_out_packed[15:0];
	assign cmrg_coord_out_0_valid = ~base_outfifo_empty;
	assign proc_outfifo_in_packed[16] = eos_to_fifo;
	assign proc_outfifo_in_packed[15:0] = data_to_fifo;
	assign cmrg_coord_out_1[16] = proc_outfifo_out_packed[16];
	assign cmrg_coord_out_1[15:0] = proc_outfifo_out_packed[15:0];
	assign cmrg_coord_out_1_valid = ~proc_outfifo_empty;
	always @(posedge clk or negedge rst_n)
		if (!rst_n)
			proc_seq_current_state <= 2'h2;
		else if (clk_en) begin
			if (flush)
				proc_seq_current_state <= 2'h2;
			else
				proc_seq_current_state <= proc_seq_next_state;
		end
	always @(*) begin
		proc_seq_next_state = proc_seq_current_state;
		case (proc_seq_current_state)
			2'h0:
				if (both_done)
					proc_seq_next_state = 2'h1;
				else
					proc_seq_next_state = 2'h0;
			2'h1:
				if (~base_outfifo_full & ~proc_outfifo_full)
					proc_seq_next_state = 2'h2;
			2'h2:
				if (tile_en)
					proc_seq_next_state = 2'h0;
				else
					proc_seq_next_state = 2'h2;
			default: proc_seq_next_state = proc_seq_current_state;
		endcase
	end
	always @(*)
		case (proc_seq_current_state)
			2'h0: begin : proc_seq_DATA_SEEN_Output
				cmrg_fifo_pop[0] = (((base_eos_seen ? 1'h1 : ((base_infifo_in_valid & ~base_infifo_in_eos) & proc_infifo_in_valid) & ~proc_infifo_in_eos) & ~base_outfifo_full) & ~proc_outfifo_full) & ~base_done_seen;
				cmrg_fifo_pop[1] = (proc_eos_seen ? 1'h1 : (base_eos_seen & ~base_outfifo_full) & ~proc_outfifo_full) & ~proc_done_seen;
				cmrg_fifo_push[0] = (((base_eos_seen ? 1'h1 : ((base_infifo_in_valid & ~base_infifo_in_eos) & proc_infifo_in_valid) & ~proc_infifo_in_eos) & ~base_outfifo_full) & ~proc_outfifo_full) & ~base_done_seen;
				cmrg_fifo_push[1] = (((base_eos_seen ? 1'h1 : ((base_infifo_in_valid & ~base_infifo_in_eos) & proc_infifo_in_valid) & ~proc_infifo_in_eos) & ~base_outfifo_full) & ~proc_outfifo_full) & ~base_done_seen;
				data_to_fifo = (base_infifo_in_eos ? base_infifo_in_data : proc_infifo_in_data);
				eos_to_fifo = base_infifo_in_eos;
				clr_pushed_proc = 1'h1;
				clr_pushed_base = 1'h1;
				reg_clr = 1'h1;
				reg_hold = 1'h0;
			end
			2'h1: begin : proc_seq_DONE_Output
				cmrg_fifo_pop[0] = ~proc_outfifo_full & ~base_outfifo_full;
				cmrg_fifo_pop[1] = ~proc_outfifo_full & ~base_outfifo_full;
				cmrg_fifo_push[0] = ~proc_outfifo_full & ~base_outfifo_full;
				cmrg_fifo_push[1] = ~proc_outfifo_full & ~base_outfifo_full;
				data_to_fifo = base_infifo_in_data;
				eos_to_fifo = 1'h1;
				clr_pushed_proc = 1'h1;
				clr_pushed_base = 1'h1;
				reg_clr = 1'h1;
				reg_hold = 1'h0;
			end
			2'h2: begin : proc_seq_START_Output
				cmrg_fifo_pop[0] = 1'h0;
				cmrg_fifo_pop[1] = 1'h0;
				cmrg_fifo_push[0] = 1'h0;
				cmrg_fifo_push[1] = 1'h0;
				data_to_fifo = 16'h0000;
				eos_to_fifo = 1'h0;
				clr_pushed_proc = 1'h1;
				clr_pushed_base = 1'h1;
				reg_clr = 1'h0;
				reg_hold = 1'h0;
			end
			default: begin : proc_seq_default_Output
				cmrg_fifo_pop[0] = 1'h0;
				cmrg_fifo_pop[1] = 1'h0;
				cmrg_fifo_push[0] = 1'h0;
				cmrg_fifo_push[1] = 1'h0;
				data_to_fifo = 16'h0000;
				eos_to_fifo = 1'h0;
				clr_pushed_proc = 1'h1;
				clr_pushed_base = 1'h1;
				reg_clr = 1'h0;
				reg_hold = 1'h0;
			end
		endcase
	reg_fifo_depth_0_w_17_afd_2 base_infifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(base_infifo_in_packed),
		.flush(flush),
		.pop(cmrg_fifo_pop[0]),
		.push(cmrg_coord_in_0_valid),
		.rst_n(rst_n),
		.data_out(base_infifo_out_packed),
		.empty(base_infifo_empty),
		.full(base_infifo_full)
	);
	reg_fifo_depth_0_w_17_afd_2 proc_infifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(proc_infifo_in_packed),
		.flush(flush),
		.pop(cmrg_fifo_pop[1]),
		.push(cmrg_coord_in_1_valid),
		.rst_n(rst_n),
		.data_out(proc_infifo_out_packed),
		.empty(proc_infifo_empty),
		.full(proc_infifo_full)
	);
	reg_fifo_depth_0_w_17_afd_2 base_outfifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(base_outfifo_in_packed),
		.flush(flush),
		.pop(cmrg_coord_out_0_ready),
		.push(cmrg_fifo_push[0]),
		.rst_n(rst_n),
		.data_out(base_outfifo_out_packed),
		.empty(base_outfifo_empty),
		.full(base_outfifo_full)
	);
	reg_fifo_depth_0_w_17_afd_2 proc_outfifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(proc_outfifo_in_packed),
		.flush(flush),
		.pop(cmrg_coord_out_1_ready),
		.push(cmrg_fifo_push[1]),
		.rst_n(rst_n),
		.data_out(proc_outfifo_out_packed),
		.empty(proc_outfifo_empty),
		.full(proc_outfifo_full)
	);
endmodule
module crdhold_flat (
	clk,
	clk_en,
	cmrg_coord_in_0_f_,
	cmrg_coord_in_0_valid_f_,
	cmrg_coord_in_1_f_,
	cmrg_coord_in_1_valid_f_,
	cmrg_coord_out_0_ready_f_,
	cmrg_coord_out_1_ready_f_,
	crdhold_inst_cmrg_enable,
	crdhold_inst_cmrg_stop_lvl,
	crdhold_inst_tile_en,
	flush,
	rst_n,
	cmrg_coord_in_0_ready_f_,
	cmrg_coord_in_1_ready_f_,
	cmrg_coord_out_0_f_,
	cmrg_coord_out_0_valid_f_,
	cmrg_coord_out_1_f_,
	cmrg_coord_out_1_valid_f_
);
	input wire clk;
	input wire clk_en;
	input wire [16:0] cmrg_coord_in_0_f_;
	input wire cmrg_coord_in_0_valid_f_;
	input wire [16:0] cmrg_coord_in_1_f_;
	input wire cmrg_coord_in_1_valid_f_;
	input wire cmrg_coord_out_0_ready_f_;
	input wire cmrg_coord_out_1_ready_f_;
	input wire crdhold_inst_cmrg_enable;
	input wire [15:0] crdhold_inst_cmrg_stop_lvl;
	input wire crdhold_inst_tile_en;
	input wire flush;
	input wire rst_n;
	output wire cmrg_coord_in_0_ready_f_;
	output wire cmrg_coord_in_1_ready_f_;
	output wire [16:0] cmrg_coord_out_0_f_;
	output wire cmrg_coord_out_0_valid_f_;
	output wire [16:0] cmrg_coord_out_1_f_;
	output wire cmrg_coord_out_1_valid_f_;
	crdhold crdhold_inst(
		.clk(clk),
		.clk_en(clk_en),
		.cmrg_coord_in_0(cmrg_coord_in_0_f_),
		.cmrg_coord_in_0_valid(cmrg_coord_in_0_valid_f_),
		.cmrg_coord_in_1(cmrg_coord_in_1_f_),
		.cmrg_coord_in_1_valid(cmrg_coord_in_1_valid_f_),
		.cmrg_coord_out_0_ready(cmrg_coord_out_0_ready_f_),
		.cmrg_coord_out_1_ready(cmrg_coord_out_1_ready_f_),
		.cmrg_enable(crdhold_inst_cmrg_enable),
		.cmrg_stop_lvl(crdhold_inst_cmrg_stop_lvl),
		.flush(flush),
		.rst_n(rst_n),
		.tile_en(crdhold_inst_tile_en),
		.cmrg_coord_in_0_ready(cmrg_coord_in_0_ready_f_),
		.cmrg_coord_in_1_ready(cmrg_coord_in_1_ready_f_),
		.cmrg_coord_out_0(cmrg_coord_out_0_f_),
		.cmrg_coord_out_0_valid(cmrg_coord_out_0_valid_f_),
		.cmrg_coord_out_1(cmrg_coord_out_1_f_),
		.cmrg_coord_out_1_valid(cmrg_coord_out_1_valid_f_)
	);
endmodule
module intersect_unit (
	clk,
	clk_en,
	coord_in_0,
	coord_in_0_valid,
	coord_in_1,
	coord_in_1_valid,
	coord_out_ready,
	flush,
	joiner_op,
	pos_in_0,
	pos_in_0_valid,
	pos_in_1,
	pos_in_1_valid,
	pos_out_0_ready,
	pos_out_1_ready,
	rst_n,
	tile_en,
	coord_in_0_ready,
	coord_in_1_ready,
	coord_out,
	coord_out_valid,
	pos_in_0_ready,
	pos_in_1_ready,
	pos_out_0,
	pos_out_0_valid,
	pos_out_1,
	pos_out_1_valid
);
	input wire clk;
	input wire clk_en;
	input wire [16:0] coord_in_0;
	input wire coord_in_0_valid;
	input wire [16:0] coord_in_1;
	input wire coord_in_1_valid;
	input wire coord_out_ready;
	input wire flush;
	input wire joiner_op;
	input wire [16:0] pos_in_0;
	input wire pos_in_0_valid;
	input wire [16:0] pos_in_1;
	input wire pos_in_1_valid;
	input wire pos_out_0_ready;
	input wire pos_out_1_ready;
	input wire rst_n;
	input wire tile_en;
	output wire coord_in_0_ready;
	output wire coord_in_1_ready;
	output wire [16:0] coord_out;
	output wire coord_out_valid;
	output wire pos_in_0_ready;
	output wire pos_in_1_ready;
	output wire [16:0] pos_out_0;
	output wire pos_out_0_valid;
	output wire [16:0] pos_out_1;
	output wire pos_out_1_valid;
	wire all_valid;
	wire all_valid_join;
	wire any_eos;
	reg [1:0] clr_eos_sticky;
	wire [16:0] coord_fifo_in_packed;
	wire [16:0] coord_fifo_out_packed;
	wire coord_in_0_fifo_eos_in;
	wire [16:0] coord_in_0_fifo_in;
	wire coord_in_0_fifo_valid_in;
	wire coord_in_1_fifo_eos_in;
	wire [16:0] coord_in_1_fifo_in;
	wire coord_in_1_fifo_valid_in;
	wire coord_in_fifo_0_empty;
	wire coord_in_fifo_0_full;
	wire coord_in_fifo_1_empty;
	wire coord_in_fifo_1_full;
	reg [15:0] coord_to_fifo;
	reg coord_to_fifo_eos;
	wire coordinate_fifo_empty;
	wire coordinate_fifo_full;
	wire [1:0] eos_in_sticky;
	wire eos_sticky_0_sticky;
	reg eos_sticky_0_was_high;
	wire eos_sticky_1_sticky;
	reg eos_sticky_1_was_high;
	wire [2:0] fifo_full;
	reg fifo_push;
	wire gclk;
	reg [1:0] inc_pos_cnt;
	reg [2:0] intersect_seq_current_state;
	reg [2:0] intersect_seq_next_state;
	wire [15:0] maybe;
	wire pos0_fifo_empty;
	wire pos0_fifo_full;
	wire [16:0] pos0_fifo_in_packed;
	wire [16:0] pos0_fifo_out_packed;
	wire pos1_fifo_empty;
	wire pos1_fifo_full;
	wire [16:0] pos1_fifo_in_packed;
	wire [16:0] pos1_fifo_out_packed;
	reg [31:0] pos_cnt;
	wire pos_in_0_fifo_eos_in;
	wire [16:0] pos_in_0_fifo_in;
	wire pos_in_0_fifo_valid_in;
	wire pos_in_1_fifo_eos_in;
	wire [16:0] pos_in_1_fifo_in;
	wire pos_in_1_fifo_valid_in;
	wire pos_in_fifo_0_empty;
	wire pos_in_fifo_0_full;
	wire pos_in_fifo_1_empty;
	wire pos_in_fifo_1_full;
	reg [31:0] pos_to_fifo;
	reg [1:0] pos_to_fifo_eos;
	reg [1:0] rst_pos_cnt;
	assign gclk = clk & tile_en;
	assign coord_in_0_fifo_eos_in = coord_in_0_fifo_in[16];
	assign coord_in_0_ready = ~coord_in_fifo_0_full;
	assign coord_in_0_fifo_valid_in = ~coord_in_fifo_0_empty;
	assign pos_in_0_fifo_eos_in = pos_in_0_fifo_in[16];
	assign pos_in_0_ready = ~pos_in_fifo_0_full;
	assign pos_in_0_fifo_valid_in = ~pos_in_fifo_0_empty;
	assign coord_in_1_fifo_eos_in = coord_in_1_fifo_in[16];
	assign coord_in_1_ready = ~coord_in_fifo_1_full;
	assign coord_in_1_fifo_valid_in = ~coord_in_fifo_1_empty;
	assign pos_in_1_fifo_eos_in = pos_in_1_fifo_in[16];
	assign pos_in_1_ready = ~pos_in_fifo_1_full;
	assign pos_in_1_fifo_valid_in = ~pos_in_fifo_1_empty;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			eos_sticky_0_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				eos_sticky_0_was_high <= 1'h0;
			else if (clr_eos_sticky[0])
				eos_sticky_0_was_high <= 1'h0;
			else if (((coord_in_0_fifo_eos_in & coord_in_0_fifo_valid_in) & pos_in_0_fifo_eos_in) & pos_in_0_fifo_valid_in)
				eos_sticky_0_was_high <= 1'h1;
		end
	assign eos_sticky_0_sticky = (((coord_in_0_fifo_eos_in & coord_in_0_fifo_valid_in) & pos_in_0_fifo_eos_in) & pos_in_0_fifo_valid_in) | eos_sticky_0_was_high;
	assign eos_in_sticky[0] = eos_sticky_0_sticky;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			eos_sticky_1_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				eos_sticky_1_was_high <= 1'h0;
			else if (clr_eos_sticky[1])
				eos_sticky_1_was_high <= 1'h0;
			else if (((coord_in_1_fifo_eos_in & coord_in_1_fifo_valid_in) & pos_in_1_fifo_eos_in) & pos_in_1_fifo_valid_in)
				eos_sticky_1_was_high <= 1'h1;
		end
	assign eos_sticky_1_sticky = (((coord_in_1_fifo_eos_in & coord_in_1_fifo_valid_in) & pos_in_1_fifo_eos_in) & pos_in_1_fifo_valid_in) | eos_sticky_1_was_high;
	assign eos_in_sticky[1] = eos_sticky_1_sticky;
	assign all_valid = &{coord_in_0_fifo_valid_in, coord_in_1_fifo_valid_in, pos_in_0_fifo_valid_in, pos_in_1_fifo_valid_in} & ~any_eos;
	assign all_valid_join = &{coord_in_0_fifo_valid_in, coord_in_1_fifo_valid_in, pos_in_0_fifo_valid_in, pos_in_1_fifo_valid_in};
	assign any_eos = |({coord_in_0_fifo_eos_in, coord_in_1_fifo_eos_in, pos_in_0_fifo_eos_in, pos_in_1_fifo_eos_in} & {coord_in_0_fifo_valid_in, coord_in_1_fifo_valid_in, pos_in_0_fifo_valid_in, pos_in_1_fifo_valid_in});
	assign maybe = 16'h0200;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			pos_cnt[0+:16] <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				pos_cnt[0+:16] <= 16'h0000;
			else if (rst_pos_cnt[0])
				pos_cnt[0+:16] <= 16'h0000;
			else if (inc_pos_cnt[0])
				pos_cnt[0+:16] <= pos_cnt[0+:16] + 16'h0001;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			pos_cnt[16+:16] <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				pos_cnt[16+:16] <= 16'h0000;
			else if (rst_pos_cnt[1])
				pos_cnt[16+:16] <= 16'h0000;
			else if (inc_pos_cnt[1])
				pos_cnt[16+:16] <= pos_cnt[16+:16] + 16'h0001;
		end
	assign coord_fifo_in_packed[16] = coord_to_fifo_eos;
	assign coord_fifo_in_packed[15:0] = coord_to_fifo;
	assign coord_out[16] = coord_fifo_out_packed[16];
	assign coord_out[15:0] = coord_fifo_out_packed[15:0];
	assign pos0_fifo_in_packed[16] = pos_to_fifo_eos[0];
	assign pos0_fifo_in_packed[15:0] = pos_to_fifo[0+:16];
	assign pos_out_0[16] = pos0_fifo_out_packed[16];
	assign pos_out_0[15:0] = pos0_fifo_out_packed[15:0];
	assign pos1_fifo_in_packed[16] = pos_to_fifo_eos[1];
	assign pos1_fifo_in_packed[15:0] = pos_to_fifo[16+:16];
	assign pos_out_1[16] = pos1_fifo_out_packed[16];
	assign pos_out_1[15:0] = pos1_fifo_out_packed[15:0];
	assign fifo_full[0] = coordinate_fifo_full;
	assign fifo_full[1] = pos0_fifo_full;
	assign fifo_full[2] = pos1_fifo_full;
	assign coord_out_valid = ~coordinate_fifo_empty;
	assign pos_out_0_valid = ~pos0_fifo_empty;
	assign pos_out_1_valid = ~pos1_fifo_empty;
	always @(posedge clk or negedge rst_n)
		if (!rst_n)
			intersect_seq_current_state <= 3'h3;
		else if (clk_en) begin
			if (flush)
				intersect_seq_current_state <= 3'h3;
			else
				intersect_seq_current_state <= intersect_seq_next_state;
		end
	always @(*) begin
		intersect_seq_next_state = intersect_seq_current_state;
		case (intersect_seq_current_state)
			3'h0:
				if (&eos_in_sticky)
					intersect_seq_next_state = 3'h2;
				else
					intersect_seq_next_state = 3'h0;
			3'h1: intersect_seq_next_state = 3'h3;
			3'h2:
				if (~(&({coord_in_0_fifo_eos_in, coord_in_1_fifo_eos_in, pos_in_0_fifo_eos_in, pos_in_1_fifo_eos_in} & {coord_in_0_fifo_valid_in, coord_in_1_fifo_valid_in, pos_in_0_fifo_valid_in, pos_in_1_fifo_valid_in})) & &{coord_in_0_fifo_valid_in, coord_in_1_fifo_valid_in, pos_in_0_fifo_valid_in, pos_in_1_fifo_valid_in})
					intersect_seq_next_state = 3'h1;
				else
					intersect_seq_next_state = 3'h2;
			3'h3:
				if ((all_valid_join & (joiner_op == 1'h1)) & tile_en)
					intersect_seq_next_state = 3'h5;
				else if ((any_eos & (joiner_op == 1'h0)) & tile_en)
					intersect_seq_next_state = 3'h0;
				else if ((all_valid & (joiner_op == 1'h0)) & tile_en)
					intersect_seq_next_state = 3'h4;
				else
					intersect_seq_next_state = 3'h3;
			3'h4:
				if (any_eos)
					intersect_seq_next_state = 3'h0;
				else
					intersect_seq_next_state = 3'h4;
			3'h5:
				if (&eos_in_sticky)
					intersect_seq_next_state = 3'h2;
				else
					intersect_seq_next_state = 3'h5;
			default: intersect_seq_next_state = intersect_seq_current_state;
		endcase
	end
	always @(*)
		case (intersect_seq_current_state)
			3'h0: begin : intersect_seq_ALIGN_Output
				inc_pos_cnt[0] = (~eos_in_sticky[0] & coord_in_0_fifo_valid_in) & pos_in_0_fifo_valid_in;
				inc_pos_cnt[1] = (~eos_in_sticky[1] & coord_in_1_fifo_valid_in) & pos_in_1_fifo_valid_in;
				rst_pos_cnt[0] = 1'h0;
				rst_pos_cnt[1] = 1'h0;
				fifo_push = 1'h0;
				clr_eos_sticky[0] = 1'h0;
				clr_eos_sticky[1] = 1'h0;
				coord_to_fifo = 16'h0000;
				pos_to_fifo[0+:16] = 16'h0000;
				pos_to_fifo[16+:16] = 16'h0000;
				coord_to_fifo_eos = 1'h0;
				pos_to_fifo_eos[0] = 1'h0;
				pos_to_fifo_eos[1] = 1'h0;
			end
			3'h1: begin : intersect_seq_DONE_Output
				inc_pos_cnt[0] = 1'h0;
				inc_pos_cnt[1] = 1'h0;
				rst_pos_cnt[0] = 1'h1;
				rst_pos_cnt[1] = 1'h1;
				fifo_push = 1'h0;
				clr_eos_sticky[0] = 1'h1;
				clr_eos_sticky[1] = 1'h1;
				coord_to_fifo = 16'h0000;
				pos_to_fifo[0+:16] = 16'h0000;
				pos_to_fifo[16+:16] = 16'h0000;
				coord_to_fifo_eos = 1'h0;
				pos_to_fifo_eos[0] = 1'h0;
				pos_to_fifo_eos[1] = 1'h0;
			end
			3'h2: begin : intersect_seq_DRAIN_Output
				inc_pos_cnt[0] = (~(|fifo_full) & &({coord_in_0_fifo_eos_in, coord_in_1_fifo_eos_in, pos_in_0_fifo_eos_in, pos_in_1_fifo_eos_in} & {coord_in_0_fifo_valid_in, coord_in_1_fifo_valid_in, pos_in_0_fifo_valid_in, pos_in_1_fifo_valid_in})) & &{coord_in_0_fifo_valid_in, coord_in_1_fifo_valid_in, pos_in_0_fifo_valid_in, pos_in_1_fifo_valid_in};
				inc_pos_cnt[1] = (~(|fifo_full) & &({coord_in_0_fifo_eos_in, coord_in_1_fifo_eos_in, pos_in_0_fifo_eos_in, pos_in_1_fifo_eos_in} & {coord_in_0_fifo_valid_in, coord_in_1_fifo_valid_in, pos_in_0_fifo_valid_in, pos_in_1_fifo_valid_in})) & &{coord_in_0_fifo_valid_in, coord_in_1_fifo_valid_in, pos_in_0_fifo_valid_in, pos_in_1_fifo_valid_in};
				rst_pos_cnt[0] = 1'h0;
				rst_pos_cnt[1] = 1'h0;
				fifo_push = (~(|fifo_full) & &({coord_in_0_fifo_eos_in, coord_in_1_fifo_eos_in, pos_in_0_fifo_eos_in, pos_in_1_fifo_eos_in} & {coord_in_0_fifo_valid_in, coord_in_1_fifo_valid_in, pos_in_0_fifo_valid_in, pos_in_1_fifo_valid_in})) & &{coord_in_0_fifo_valid_in, coord_in_1_fifo_valid_in, pos_in_0_fifo_valid_in, pos_in_1_fifo_valid_in};
				clr_eos_sticky[0] = 1'h0;
				clr_eos_sticky[1] = 1'h0;
				coord_to_fifo = coord_in_0_fifo_in[15:0];
				pos_to_fifo[0+:16] = coord_in_0_fifo_in[15:0];
				pos_to_fifo[16+:16] = coord_in_0_fifo_in[15:0];
				coord_to_fifo_eos = any_eos;
				pos_to_fifo_eos[0] = any_eos;
				pos_to_fifo_eos[1] = any_eos;
			end
			3'h3: begin : intersect_seq_IDLE_Output
				inc_pos_cnt[0] = 1'h0;
				inc_pos_cnt[1] = 1'h0;
				rst_pos_cnt[0] = 1'h0;
				rst_pos_cnt[1] = 1'h0;
				fifo_push = 1'h0;
				clr_eos_sticky[0] = 1'h0;
				clr_eos_sticky[1] = 1'h0;
				coord_to_fifo = 16'h0000;
				pos_to_fifo[0+:16] = 16'h0000;
				pos_to_fifo[16+:16] = 16'h0000;
				coord_to_fifo_eos = 1'h0;
				pos_to_fifo_eos[0] = 1'h0;
				pos_to_fifo_eos[1] = 1'h0;
			end
			3'h4: begin : intersect_seq_ITER_Output
				inc_pos_cnt[0] = (all_valid & (coord_in_0_fifo_in <= coord_in_1_fifo_in)) & ~(|fifo_full);
				inc_pos_cnt[1] = (all_valid & (coord_in_0_fifo_in >= coord_in_1_fifo_in)) & ~(|fifo_full);
				rst_pos_cnt[0] = any_eos & ~(|fifo_full);
				rst_pos_cnt[1] = any_eos & ~(|fifo_full);
				fifo_push = ((all_valid & (coord_in_0_fifo_in == coord_in_1_fifo_in)) & ~(|fifo_full)) & ~any_eos;
				clr_eos_sticky[0] = 1'h0;
				clr_eos_sticky[1] = 1'h0;
				coord_to_fifo = coord_in_0_fifo_in[15:0];
				pos_to_fifo[0+:16] = pos_in_0_fifo_in[15:0];
				pos_to_fifo[16+:16] = pos_in_1_fifo_in[15:0];
				coord_to_fifo_eos = 1'h0;
				pos_to_fifo_eos[0] = 1'h0;
				pos_to_fifo_eos[1] = 1'h0;
			end
			3'h5: begin : intersect_seq_UNION_Output
				inc_pos_cnt[0] = ((all_valid_join & ((coord_in_0_fifo_in <= coord_in_1_fifo_in) | coord_in_1_fifo_eos_in)) & ~(|fifo_full)) & ~coord_in_0_fifo_eos_in;
				inc_pos_cnt[1] = ((all_valid_join & ((coord_in_0_fifo_in >= coord_in_1_fifo_in) | coord_in_0_fifo_eos_in)) & ~(|fifo_full)) & ~coord_in_1_fifo_eos_in;
				rst_pos_cnt[0] = any_eos & ~(|fifo_full);
				rst_pos_cnt[1] = any_eos & ~(|fifo_full);
				fifo_push = (all_valid_join & ~(|fifo_full)) & ~(&({coord_in_0_fifo_eos_in, coord_in_1_fifo_eos_in, pos_in_0_fifo_eos_in, pos_in_1_fifo_eos_in} & {coord_in_0_fifo_valid_in, coord_in_1_fifo_valid_in, pos_in_0_fifo_valid_in, pos_in_1_fifo_valid_in}));
				clr_eos_sticky[0] = 1'h0;
				clr_eos_sticky[1] = 1'h0;
				coord_to_fifo = (coord_in_0_fifo_eos_in ? coord_in_1_fifo_in[15:0] : (coord_in_1_fifo_eos_in ? coord_in_0_fifo_in[15:0] : (coord_in_0_fifo_in <= coord_in_1_fifo_in ? coord_in_0_fifo_in[15:0] : coord_in_1_fifo_in[15:0])));
				pos_to_fifo[0+:16] = (coord_in_0_fifo_eos_in ? maybe : (coord_in_1_fifo_eos_in ? pos_in_0_fifo_in[15:0] : (coord_in_0_fifo_in <= coord_in_1_fifo_in ? pos_in_0_fifo_in[15:0] : maybe)));
				pos_to_fifo[16+:16] = (coord_in_1_fifo_eos_in ? maybe : (coord_in_0_fifo_eos_in ? pos_in_1_fifo_in[15:0] : (coord_in_1_fifo_in <= coord_in_0_fifo_in ? pos_in_1_fifo_in[15:0] : maybe)));
				coord_to_fifo_eos = 1'h0;
				pos_to_fifo_eos[0] = (pos_in_0_fifo_eos_in & ~coord_in_0_fifo_eos_in) | (coord_in_0_fifo_eos_in ? 1'h1 : (coord_in_1_fifo_eos_in ? 1'h0 : (coord_in_0_fifo_in <= coord_in_1_fifo_in ? 1'h0 : 1'h1)));
				pos_to_fifo_eos[1] = (pos_in_1_fifo_eos_in & ~coord_in_1_fifo_eos_in) | (coord_in_1_fifo_eos_in ? 1'h1 : (coord_in_0_fifo_eos_in ? 1'h0 : (coord_in_1_fifo_in <= coord_in_0_fifo_in ? 1'h0 : 1'h1)));
			end
			default: begin : intersect_seq_default_Output
				inc_pos_cnt[0] = 1'h0;
				inc_pos_cnt[1] = 1'h0;
				rst_pos_cnt[0] = 1'h0;
				rst_pos_cnt[1] = 1'h0;
				fifo_push = 1'h0;
				clr_eos_sticky[0] = 1'h0;
				clr_eos_sticky[1] = 1'h0;
				coord_to_fifo = 16'h0000;
				pos_to_fifo[0+:16] = 16'h0000;
				pos_to_fifo[16+:16] = 16'h0000;
				coord_to_fifo_eos = 1'h0;
				pos_to_fifo_eos[0] = 1'h0;
				pos_to_fifo_eos[1] = 1'h0;
			end
		endcase
	reg_fifo_depth_0_w_17_afd_2 coord_in_fifo_0(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(coord_in_0),
		.flush(flush),
		.pop(inc_pos_cnt[0]),
		.push(coord_in_0_valid),
		.rst_n(rst_n),
		.data_out(coord_in_0_fifo_in),
		.empty(coord_in_fifo_0_empty),
		.full(coord_in_fifo_0_full)
	);
	reg_fifo_depth_0_w_17_afd_2 pos_in_fifo_0(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(pos_in_0),
		.flush(flush),
		.pop(inc_pos_cnt[0]),
		.push(pos_in_0_valid),
		.rst_n(rst_n),
		.data_out(pos_in_0_fifo_in),
		.empty(pos_in_fifo_0_empty),
		.full(pos_in_fifo_0_full)
	);
	reg_fifo_depth_0_w_17_afd_2 coord_in_fifo_1(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(coord_in_1),
		.flush(flush),
		.pop(inc_pos_cnt[1]),
		.push(coord_in_1_valid),
		.rst_n(rst_n),
		.data_out(coord_in_1_fifo_in),
		.empty(coord_in_fifo_1_empty),
		.full(coord_in_fifo_1_full)
	);
	reg_fifo_depth_0_w_17_afd_2 pos_in_fifo_1(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(pos_in_1),
		.flush(flush),
		.pop(inc_pos_cnt[1]),
		.push(pos_in_1_valid),
		.rst_n(rst_n),
		.data_out(pos_in_1_fifo_in),
		.empty(pos_in_fifo_1_empty),
		.full(pos_in_fifo_1_full)
	);
	reg_fifo_depth_0_w_17_afd_2 coordinate_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(coord_fifo_in_packed),
		.flush(flush),
		.pop(coord_out_ready),
		.push(fifo_push),
		.rst_n(rst_n),
		.data_out(coord_fifo_out_packed),
		.empty(coordinate_fifo_empty),
		.full(coordinate_fifo_full)
	);
	reg_fifo_depth_0_w_17_afd_2 pos0_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(pos0_fifo_in_packed),
		.flush(flush),
		.pop(pos_out_0_ready),
		.push(fifo_push),
		.rst_n(rst_n),
		.data_out(pos0_fifo_out_packed),
		.empty(pos0_fifo_empty),
		.full(pos0_fifo_full)
	);
	reg_fifo_depth_0_w_17_afd_2 pos1_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(pos1_fifo_in_packed),
		.flush(flush),
		.pop(pos_out_1_ready),
		.push(fifo_push),
		.rst_n(rst_n),
		.data_out(pos1_fifo_out_packed),
		.empty(pos1_fifo_empty),
		.full(pos1_fifo_full)
	);
endmodule
module intersect_unit_flat (
	clk,
	clk_en,
	coord_in_0_f_,
	coord_in_0_valid_f_,
	coord_in_1_f_,
	coord_in_1_valid_f_,
	coord_out_ready_f_,
	flush,
	intersect_unit_inst_joiner_op,
	intersect_unit_inst_tile_en,
	pos_in_0_f_,
	pos_in_0_valid_f_,
	pos_in_1_f_,
	pos_in_1_valid_f_,
	pos_out_0_ready_f_,
	pos_out_1_ready_f_,
	rst_n,
	coord_in_0_ready_f_,
	coord_in_1_ready_f_,
	coord_out_f_,
	coord_out_valid_f_,
	pos_in_0_ready_f_,
	pos_in_1_ready_f_,
	pos_out_0_f_,
	pos_out_0_valid_f_,
	pos_out_1_f_,
	pos_out_1_valid_f_
);
	input wire clk;
	input wire clk_en;
	input wire [16:0] coord_in_0_f_;
	input wire coord_in_0_valid_f_;
	input wire [16:0] coord_in_1_f_;
	input wire coord_in_1_valid_f_;
	input wire coord_out_ready_f_;
	input wire flush;
	input wire intersect_unit_inst_joiner_op;
	input wire intersect_unit_inst_tile_en;
	input wire [16:0] pos_in_0_f_;
	input wire pos_in_0_valid_f_;
	input wire [16:0] pos_in_1_f_;
	input wire pos_in_1_valid_f_;
	input wire pos_out_0_ready_f_;
	input wire pos_out_1_ready_f_;
	input wire rst_n;
	output wire coord_in_0_ready_f_;
	output wire coord_in_1_ready_f_;
	output wire [16:0] coord_out_f_;
	output wire coord_out_valid_f_;
	output wire pos_in_0_ready_f_;
	output wire pos_in_1_ready_f_;
	output wire [16:0] pos_out_0_f_;
	output wire pos_out_0_valid_f_;
	output wire [16:0] pos_out_1_f_;
	output wire pos_out_1_valid_f_;
	intersect_unit intersect_unit_inst(
		.clk(clk),
		.clk_en(clk_en),
		.coord_in_0(coord_in_0_f_),
		.coord_in_0_valid(coord_in_0_valid_f_),
		.coord_in_1(coord_in_1_f_),
		.coord_in_1_valid(coord_in_1_valid_f_),
		.coord_out_ready(coord_out_ready_f_),
		.flush(flush),
		.joiner_op(intersect_unit_inst_joiner_op),
		.pos_in_0(pos_in_0_f_),
		.pos_in_0_valid(pos_in_0_valid_f_),
		.pos_in_1(pos_in_1_f_),
		.pos_in_1_valid(pos_in_1_valid_f_),
		.pos_out_0_ready(pos_out_0_ready_f_),
		.pos_out_1_ready(pos_out_1_ready_f_),
		.rst_n(rst_n),
		.tile_en(intersect_unit_inst_tile_en),
		.coord_in_0_ready(coord_in_0_ready_f_),
		.coord_in_1_ready(coord_in_1_ready_f_),
		.coord_out(coord_out_f_),
		.coord_out_valid(coord_out_valid_f_),
		.pos_in_0_ready(pos_in_0_ready_f_),
		.pos_in_1_ready(pos_in_1_ready_f_),
		.pos_out_0(pos_out_0_f_),
		.pos_out_0_valid(pos_out_0_valid_f_),
		.pos_out_1(pos_out_1_f_),
		.pos_out_1_valid(pos_out_1_valid_f_)
	);
endmodule
module reg_cr (
	clk,
	clk_en,
	data_in,
	data_in_valid,
	data_out_ready,
	default_value,
	flush,
	rst_n,
	stop_lvl,
	tile_en,
	data_in_ready,
	data_out,
	data_out_valid
);
	input wire clk;
	input wire clk_en;
	input wire [16:0] data_in;
	input wire data_in_valid;
	input wire data_out_ready;
	input wire [15:0] default_value;
	input wire flush;
	input wire rst_n;
	input wire [15:0] stop_lvl;
	input wire tile_en;
	output wire data_in_ready;
	output wire [16:0] data_out;
	output wire data_out_valid;
	reg [15:0] accum_reg;
	reg [2:0] accum_seq_current_state;
	reg [2:0] accum_seq_next_state;
	reg clr_once_popped;
	reg [15:0] data_to_fifo;
	wire gclk;
	wire [16:0] infifo_in_packed;
	wire [15:0] infifo_out_data;
	wire infifo_out_eos;
	wire [16:0] infifo_out_packed;
	wire infifo_out_valid;
	reg infifo_pop;
	wire infifo_push;
	wire input_fifo_empty;
	wire input_fifo_full;
	wire outfifo_full;
	reg outfifo_in_eos;
	wire [16:0] outfifo_in_packed;
	wire [16:0] outfifo_out_packed;
	wire outfifo_pop;
	reg outfifo_push;
	wire output_fifo_empty;
	reg reg_accum;
	reg reg_clr;
	reg set_once_popped;
	wire set_once_popped_sticky;
	reg set_once_popped_was_high;
	assign gclk = clk & tile_en;
	assign data_in_ready = ~input_fifo_full;
	assign infifo_in_packed[16:0] = data_in;
	assign infifo_out_eos = infifo_out_packed[16];
	assign infifo_out_data = infifo_out_packed[15:0];
	assign infifo_push = data_in_valid;
	assign infifo_out_valid = ~input_fifo_empty;
	assign outfifo_in_packed[16] = outfifo_in_eos;
	assign outfifo_in_packed[15:0] = data_to_fifo;
	assign data_out = outfifo_out_packed[16:0];
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			set_once_popped_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				set_once_popped_was_high <= 1'h0;
			else if (clr_once_popped)
				set_once_popped_was_high <= 1'h0;
			else if (set_once_popped)
				set_once_popped_was_high <= 1'h1;
		end
	assign set_once_popped_sticky = set_once_popped_was_high;
	assign data_out_valid = ~output_fifo_empty;
	assign outfifo_pop = data_out_ready;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			accum_reg <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				accum_reg <= 16'h0000;
			else if (reg_clr)
				accum_reg <= default_value;
			else if (reg_accum)
				accum_reg <= accum_reg + infifo_out_data;
		end
	always @(posedge clk or negedge rst_n)
		if (!rst_n)
			accum_seq_current_state <= 3'h3;
		else if (clk_en) begin
			if (flush)
				accum_seq_current_state <= 3'h3;
			else
				accum_seq_current_state <= accum_seq_next_state;
		end
	always @(*) begin
		accum_seq_next_state = accum_seq_current_state;
		case (accum_seq_current_state)
			3'h0:
				if (infifo_out_valid & infifo_out_eos)
					accum_seq_next_state = 3'h2;
				else
					accum_seq_next_state = 3'h0;
			3'h1:
				if (~outfifo_full)
					accum_seq_next_state = 3'h3;
				else
					accum_seq_next_state = 3'h1;
			3'h2:
				if (~outfifo_full)
					accum_seq_next_state = 3'h4;
				else
					accum_seq_next_state = 3'h2;
			3'h3:
				if (infifo_out_valid & ~infifo_out_eos)
					accum_seq_next_state = 3'h0;
				else if ((infifo_out_valid & infifo_out_eos) & (infifo_out_data[9:8] == 2'h1))
					accum_seq_next_state = 3'h1;
				else if ((infifo_out_valid & infifo_out_eos) & (infifo_out_data[9:8] == 2'h0))
					accum_seq_next_state = 3'h2;
				else
					accum_seq_next_state = 3'h3;
			3'h4:
				if (~outfifo_full)
					accum_seq_next_state = 3'h3;
				else
					accum_seq_next_state = 3'h4;
			default: accum_seq_next_state = accum_seq_current_state;
		endcase
	end
	always @(*)
		case (accum_seq_current_state)
			3'h0: begin : accum_seq_ACCUM_Output
				infifo_pop = infifo_out_valid & ~infifo_out_eos;
				outfifo_push = 1'h0;
				reg_clr = 1'h0;
				reg_accum = infifo_out_valid & ~infifo_out_eos;
				data_to_fifo = 16'h0000;
				outfifo_in_eos = 1'h0;
				set_once_popped = 1'h0;
				clr_once_popped = 1'h0;
			end
			3'h1: begin : accum_seq_DONE_Output
				infifo_pop = ~outfifo_full;
				outfifo_push = ~outfifo_full;
				reg_clr = 1'h1;
				reg_accum = 1'h0;
				data_to_fifo = infifo_out_data;
				outfifo_in_eos = infifo_out_eos;
				set_once_popped = 1'h0;
				clr_once_popped = 1'h1;
			end
			3'h2: begin : accum_seq_OUTPUT_Output
				infifo_pop = 1'h0;
				outfifo_push = ~outfifo_full;
				reg_clr = 1'h0;
				reg_accum = 1'h0;
				data_to_fifo = accum_reg;
				outfifo_in_eos = 1'h0;
				set_once_popped = 1'h0;
				clr_once_popped = 1'h0;
			end
			3'h3: begin : accum_seq_START_Output
				infifo_pop = 1'h0;
				outfifo_push = 1'h0;
				reg_clr = 1'h0;
				reg_accum = 1'h0;
				data_to_fifo = 16'h0000;
				outfifo_in_eos = 1'h0;
				set_once_popped = 1'h0;
				clr_once_popped = 1'h0;
			end
			3'h4: begin : accum_seq_STOP_PASS_Output
				infifo_pop = ((~outfifo_full & infifo_out_valid) & infifo_out_eos) & (infifo_out_data[9:8] == 2'h0);
				outfifo_push = (((~outfifo_full & infifo_out_valid) & infifo_out_eos) & (infifo_out_data[9:8] == 2'h0)) & (infifo_out_data[7:0] > 8'h00);
				reg_clr = 1'h1;
				reg_accum = 1'h0;
				data_to_fifo = infifo_out_data - 16'h0001;
				outfifo_in_eos = 1'h1;
				set_once_popped = 1'h0;
				clr_once_popped = 1'h1;
			end
			default: begin : accum_seq_default_Output
				infifo_pop = 1'h0;
				outfifo_push = 1'h0;
				reg_clr = 1'h0;
				reg_accum = 1'h0;
				data_to_fifo = 16'h0000;
				outfifo_in_eos = 1'h0;
				set_once_popped = 1'h0;
				clr_once_popped = 1'h0;
			end
		endcase
	reg_fifo_depth_0_w_17_afd_2 input_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(infifo_in_packed),
		.flush(flush),
		.pop(infifo_pop),
		.push(infifo_push),
		.rst_n(rst_n),
		.data_out(infifo_out_packed),
		.empty(input_fifo_empty),
		.full(input_fifo_full)
	);
	reg_fifo_depth_0_w_17_afd_2 output_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(outfifo_in_packed),
		.flush(flush),
		.pop(outfifo_pop),
		.push(outfifo_push),
		.rst_n(rst_n),
		.data_out(outfifo_out_packed),
		.empty(output_fifo_empty),
		.full(outfifo_full)
	);
endmodule
module reg_cr_flat (
	clk,
	clk_en,
	data_in_f_,
	data_in_valid_f_,
	data_out_ready_f_,
	flush,
	reg_cr_inst_default_value,
	reg_cr_inst_stop_lvl,
	reg_cr_inst_tile_en,
	rst_n,
	data_in_ready_f_,
	data_out_f_,
	data_out_valid_f_
);
	input wire clk;
	input wire clk_en;
	input wire [16:0] data_in_f_;
	input wire data_in_valid_f_;
	input wire data_out_ready_f_;
	input wire flush;
	input wire [15:0] reg_cr_inst_default_value;
	input wire [15:0] reg_cr_inst_stop_lvl;
	input wire reg_cr_inst_tile_en;
	input wire rst_n;
	output wire data_in_ready_f_;
	output wire [16:0] data_out_f_;
	output wire data_out_valid_f_;
	reg_cr reg_cr_inst(
		.clk(clk),
		.clk_en(clk_en),
		.data_in(data_in_f_),
		.data_in_valid(data_in_valid_f_),
		.data_out_ready(data_out_ready_f_),
		.default_value(reg_cr_inst_default_value),
		.flush(flush),
		.rst_n(rst_n),
		.stop_lvl(reg_cr_inst_stop_lvl),
		.tile_en(reg_cr_inst_tile_en),
		.data_in_ready(data_in_ready_f_),
		.data_out(data_out_f_),
		.data_out_valid(data_out_valid_f_)
	);
endmodule
module reg_fifo_depth_0_w_17_afd_2 (
	clk,
	clk_en,
	data_in,
	flush,
	pop,
	push,
	rst_n,
	almost_full,
	data_out,
	empty,
	full,
	valid
);
	input wire clk;
	input wire clk_en;
	input wire [16:0] data_in;
	input wire flush;
	input wire pop;
	input wire push;
	input wire rst_n;
	output wire almost_full;
	output wire [16:0] data_out;
	output wire empty;
	output wire full;
	output wire valid;
	assign data_out = data_in;
	assign valid = push;
	assign empty = ~push;
	assign full = ~pop;
	assign almost_full = ~pop;
endmodule
module reg_fifo_depth_2_w_17_afd_2 (
	clk,
	clk_en,
	data_in,
	flush,
	pop,
	push,
	rst_n,
	almost_full,
	data_out,
	empty,
	full,
	valid
);
	input wire clk;
	input wire clk_en;
	input wire [16:0] data_in;
	input wire flush;
	input wire pop;
	input wire push;
	input wire rst_n;
	output wire almost_full;
	output reg [16:0] data_out;
	output wire empty;
	output wire full;
	output reg valid;
	reg [1:0] num_items;
	wire passthru;
	reg rd_ptr;
	wire read;
	reg [33:0] reg_array;
	reg wr_ptr;
	wire write;
	assign full = num_items == 2'h2;
	assign almost_full = num_items >= 2'h0;
	assign empty = num_items == 2'h0;
	assign read = (pop & ~passthru) & ~empty;
	assign passthru = 1'h0;
	assign write = (push & ~passthru) & ~full;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			num_items <= 2'h0;
		else if (flush)
			num_items <= 2'h0;
		else if (clk_en) begin
			if (write & ~read)
				num_items <= num_items + 2'h1;
			else if (~write & read)
				num_items <= num_items - 2'h1;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			reg_array <= 34'h000000000;
		else if (flush)
			reg_array <= 34'h000000000;
		else if (clk_en) begin
			if (write)
				reg_array[17 * wr_ptr+:17] <= data_in;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			wr_ptr <= 1'h0;
		else if (flush)
			wr_ptr <= 1'h0;
		else if (clk_en) begin
			if (write) begin
				if (wr_ptr == 1'h1)
					wr_ptr <= 1'h0;
				else
					wr_ptr <= wr_ptr + 1'h1;
			end
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			rd_ptr <= 1'h0;
		else if (flush)
			rd_ptr <= 1'h0;
		else if (clk_en) begin
			if (read)
				rd_ptr <= rd_ptr + 1'h1;
		end
	always @(*)
		if (passthru)
			data_out = data_in;
		else
			data_out = reg_array[17 * rd_ptr+:17];
	always @(*) valid = ~empty | passthru;
endmodule
module Or4x32 (
	I0,
	I1,
	I2,
	I3,
	O
);
	input [31:0] I0;
	input [31:0] I1;
	input [31:0] I2;
	input [31:0] I3;
	output wire [31:0] O;
	wire orr_inst0_out;
	wire orr_inst1_out;
	wire orr_inst10_out;
	wire orr_inst11_out;
	wire orr_inst12_out;
	wire orr_inst13_out;
	wire orr_inst14_out;
	wire orr_inst15_out;
	wire orr_inst16_out;
	wire orr_inst17_out;
	wire orr_inst18_out;
	wire orr_inst19_out;
	wire orr_inst2_out;
	wire orr_inst20_out;
	wire orr_inst21_out;
	wire orr_inst22_out;
	wire orr_inst23_out;
	wire orr_inst24_out;
	wire orr_inst25_out;
	wire orr_inst26_out;
	wire orr_inst27_out;
	wire orr_inst28_out;
	wire orr_inst29_out;
	wire orr_inst3_out;
	wire orr_inst30_out;
	wire orr_inst31_out;
	wire orr_inst4_out;
	wire orr_inst5_out;
	wire orr_inst6_out;
	wire orr_inst7_out;
	wire orr_inst8_out;
	wire orr_inst9_out;
	wire [3:0] orr_inst0_in;
	assign orr_inst0_in = {I3[0], I2[0], I1[0], I0[0]};
	coreir_orr #(.width(4)) orr_inst0(
		.in(orr_inst0_in),
		.out(orr_inst0_out)
	);
	wire [3:0] orr_inst1_in;
	assign orr_inst1_in = {I3[1], I2[1], I1[1], I0[1]};
	coreir_orr #(.width(4)) orr_inst1(
		.in(orr_inst1_in),
		.out(orr_inst1_out)
	);
	wire [3:0] orr_inst10_in;
	assign orr_inst10_in = {I3[10], I2[10], I1[10], I0[10]};
	coreir_orr #(.width(4)) orr_inst10(
		.in(orr_inst10_in),
		.out(orr_inst10_out)
	);
	wire [3:0] orr_inst11_in;
	assign orr_inst11_in = {I3[11], I2[11], I1[11], I0[11]};
	coreir_orr #(.width(4)) orr_inst11(
		.in(orr_inst11_in),
		.out(orr_inst11_out)
	);
	wire [3:0] orr_inst12_in;
	assign orr_inst12_in = {I3[12], I2[12], I1[12], I0[12]};
	coreir_orr #(.width(4)) orr_inst12(
		.in(orr_inst12_in),
		.out(orr_inst12_out)
	);
	wire [3:0] orr_inst13_in;
	assign orr_inst13_in = {I3[13], I2[13], I1[13], I0[13]};
	coreir_orr #(.width(4)) orr_inst13(
		.in(orr_inst13_in),
		.out(orr_inst13_out)
	);
	wire [3:0] orr_inst14_in;
	assign orr_inst14_in = {I3[14], I2[14], I1[14], I0[14]};
	coreir_orr #(.width(4)) orr_inst14(
		.in(orr_inst14_in),
		.out(orr_inst14_out)
	);
	wire [3:0] orr_inst15_in;
	assign orr_inst15_in = {I3[15], I2[15], I1[15], I0[15]};
	coreir_orr #(.width(4)) orr_inst15(
		.in(orr_inst15_in),
		.out(orr_inst15_out)
	);
	wire [3:0] orr_inst16_in;
	assign orr_inst16_in = {I3[16], I2[16], I1[16], I0[16]};
	coreir_orr #(.width(4)) orr_inst16(
		.in(orr_inst16_in),
		.out(orr_inst16_out)
	);
	wire [3:0] orr_inst17_in;
	assign orr_inst17_in = {I3[17], I2[17], I1[17], I0[17]};
	coreir_orr #(.width(4)) orr_inst17(
		.in(orr_inst17_in),
		.out(orr_inst17_out)
	);
	wire [3:0] orr_inst18_in;
	assign orr_inst18_in = {I3[18], I2[18], I1[18], I0[18]};
	coreir_orr #(.width(4)) orr_inst18(
		.in(orr_inst18_in),
		.out(orr_inst18_out)
	);
	wire [3:0] orr_inst19_in;
	assign orr_inst19_in = {I3[19], I2[19], I1[19], I0[19]};
	coreir_orr #(.width(4)) orr_inst19(
		.in(orr_inst19_in),
		.out(orr_inst19_out)
	);
	wire [3:0] orr_inst2_in;
	assign orr_inst2_in = {I3[2], I2[2], I1[2], I0[2]};
	coreir_orr #(.width(4)) orr_inst2(
		.in(orr_inst2_in),
		.out(orr_inst2_out)
	);
	wire [3:0] orr_inst20_in;
	assign orr_inst20_in = {I3[20], I2[20], I1[20], I0[20]};
	coreir_orr #(.width(4)) orr_inst20(
		.in(orr_inst20_in),
		.out(orr_inst20_out)
	);
	wire [3:0] orr_inst21_in;
	assign orr_inst21_in = {I3[21], I2[21], I1[21], I0[21]};
	coreir_orr #(.width(4)) orr_inst21(
		.in(orr_inst21_in),
		.out(orr_inst21_out)
	);
	wire [3:0] orr_inst22_in;
	assign orr_inst22_in = {I3[22], I2[22], I1[22], I0[22]};
	coreir_orr #(.width(4)) orr_inst22(
		.in(orr_inst22_in),
		.out(orr_inst22_out)
	);
	wire [3:0] orr_inst23_in;
	assign orr_inst23_in = {I3[23], I2[23], I1[23], I0[23]};
	coreir_orr #(.width(4)) orr_inst23(
		.in(orr_inst23_in),
		.out(orr_inst23_out)
	);
	wire [3:0] orr_inst24_in;
	assign orr_inst24_in = {I3[24], I2[24], I1[24], I0[24]};
	coreir_orr #(.width(4)) orr_inst24(
		.in(orr_inst24_in),
		.out(orr_inst24_out)
	);
	wire [3:0] orr_inst25_in;
	assign orr_inst25_in = {I3[25], I2[25], I1[25], I0[25]};
	coreir_orr #(.width(4)) orr_inst25(
		.in(orr_inst25_in),
		.out(orr_inst25_out)
	);
	wire [3:0] orr_inst26_in;
	assign orr_inst26_in = {I3[26], I2[26], I1[26], I0[26]};
	coreir_orr #(.width(4)) orr_inst26(
		.in(orr_inst26_in),
		.out(orr_inst26_out)
	);
	wire [3:0] orr_inst27_in;
	assign orr_inst27_in = {I3[27], I2[27], I1[27], I0[27]};
	coreir_orr #(.width(4)) orr_inst27(
		.in(orr_inst27_in),
		.out(orr_inst27_out)
	);
	wire [3:0] orr_inst28_in;
	assign orr_inst28_in = {I3[28], I2[28], I1[28], I0[28]};
	coreir_orr #(.width(4)) orr_inst28(
		.in(orr_inst28_in),
		.out(orr_inst28_out)
	);
	wire [3:0] orr_inst29_in;
	assign orr_inst29_in = {I3[29], I2[29], I1[29], I0[29]};
	coreir_orr #(.width(4)) orr_inst29(
		.in(orr_inst29_in),
		.out(orr_inst29_out)
	);
	wire [3:0] orr_inst3_in;
	assign orr_inst3_in = {I3[3], I2[3], I1[3], I0[3]};
	coreir_orr #(.width(4)) orr_inst3(
		.in(orr_inst3_in),
		.out(orr_inst3_out)
	);
	wire [3:0] orr_inst30_in;
	assign orr_inst30_in = {I3[30], I2[30], I1[30], I0[30]};
	coreir_orr #(.width(4)) orr_inst30(
		.in(orr_inst30_in),
		.out(orr_inst30_out)
	);
	wire [3:0] orr_inst31_in;
	assign orr_inst31_in = {I3[31], I2[31], I1[31], I0[31]};
	coreir_orr #(.width(4)) orr_inst31(
		.in(orr_inst31_in),
		.out(orr_inst31_out)
	);
	wire [3:0] orr_inst4_in;
	assign orr_inst4_in = {I3[4], I2[4], I1[4], I0[4]};
	coreir_orr #(.width(4)) orr_inst4(
		.in(orr_inst4_in),
		.out(orr_inst4_out)
	);
	wire [3:0] orr_inst5_in;
	assign orr_inst5_in = {I3[5], I2[5], I1[5], I0[5]};
	coreir_orr #(.width(4)) orr_inst5(
		.in(orr_inst5_in),
		.out(orr_inst5_out)
	);
	wire [3:0] orr_inst6_in;
	assign orr_inst6_in = {I3[6], I2[6], I1[6], I0[6]};
	coreir_orr #(.width(4)) orr_inst6(
		.in(orr_inst6_in),
		.out(orr_inst6_out)
	);
	wire [3:0] orr_inst7_in;
	assign orr_inst7_in = {I3[7], I2[7], I1[7], I0[7]};
	coreir_orr #(.width(4)) orr_inst7(
		.in(orr_inst7_in),
		.out(orr_inst7_out)
	);
	wire [3:0] orr_inst8_in;
	assign orr_inst8_in = {I3[8], I2[8], I1[8], I0[8]};
	coreir_orr #(.width(4)) orr_inst8(
		.in(orr_inst8_in),
		.out(orr_inst8_out)
	);
	wire [3:0] orr_inst9_in;
	assign orr_inst9_in = {I3[9], I2[9], I1[9], I0[9]};
	coreir_orr #(.width(4)) orr_inst9(
		.in(orr_inst9_in),
		.out(orr_inst9_out)
	);
	assign O = {orr_inst31_out, orr_inst30_out, orr_inst29_out, orr_inst28_out, orr_inst27_out, orr_inst26_out, orr_inst25_out, orr_inst24_out, orr_inst23_out, orr_inst22_out, orr_inst21_out, orr_inst20_out, orr_inst19_out, orr_inst18_out, orr_inst17_out, orr_inst16_out, orr_inst15_out, orr_inst14_out, orr_inst13_out, orr_inst12_out, orr_inst11_out, orr_inst10_out, orr_inst9_out, orr_inst8_out, orr_inst7_out, orr_inst6_out, orr_inst5_out, orr_inst4_out, orr_inst3_out, orr_inst2_out, orr_inst1_out, orr_inst0_out};
endmodule
module Or3x8 (
	I0,
	I1,
	I2,
	O
);
	input [7:0] I0;
	input [7:0] I1;
	input [7:0] I2;
	output wire [7:0] O;
	wire orr_inst0_out;
	wire orr_inst1_out;
	wire orr_inst2_out;
	wire orr_inst3_out;
	wire orr_inst4_out;
	wire orr_inst5_out;
	wire orr_inst6_out;
	wire orr_inst7_out;
	wire [2:0] orr_inst0_in;
	assign orr_inst0_in = {I2[0], I1[0], I0[0]};
	coreir_orr #(.width(3)) orr_inst0(
		.in(orr_inst0_in),
		.out(orr_inst0_out)
	);
	wire [2:0] orr_inst1_in;
	assign orr_inst1_in = {I2[1], I1[1], I0[1]};
	coreir_orr #(.width(3)) orr_inst1(
		.in(orr_inst1_in),
		.out(orr_inst1_out)
	);
	wire [2:0] orr_inst2_in;
	assign orr_inst2_in = {I2[2], I1[2], I0[2]};
	coreir_orr #(.width(3)) orr_inst2(
		.in(orr_inst2_in),
		.out(orr_inst2_out)
	);
	wire [2:0] orr_inst3_in;
	assign orr_inst3_in = {I2[3], I1[3], I0[3]};
	coreir_orr #(.width(3)) orr_inst3(
		.in(orr_inst3_in),
		.out(orr_inst3_out)
	);
	wire [2:0] orr_inst4_in;
	assign orr_inst4_in = {I2[4], I1[4], I0[4]};
	coreir_orr #(.width(3)) orr_inst4(
		.in(orr_inst4_in),
		.out(orr_inst4_out)
	);
	wire [2:0] orr_inst5_in;
	assign orr_inst5_in = {I2[5], I1[5], I0[5]};
	coreir_orr #(.width(3)) orr_inst5(
		.in(orr_inst5_in),
		.out(orr_inst5_out)
	);
	wire [2:0] orr_inst6_in;
	assign orr_inst6_in = {I2[6], I1[6], I0[6]};
	coreir_orr #(.width(3)) orr_inst6(
		.in(orr_inst6_in),
		.out(orr_inst6_out)
	);
	wire [2:0] orr_inst7_in;
	assign orr_inst7_in = {I2[7], I1[7], I0[7]};
	coreir_orr #(.width(3)) orr_inst7(
		.in(orr_inst7_in),
		.out(orr_inst7_out)
	);
	assign O = {orr_inst7_out, orr_inst6_out, orr_inst5_out, orr_inst4_out, orr_inst3_out, orr_inst2_out, orr_inst1_out, orr_inst0_out};
endmodule
module Or3x32 (
	I0,
	I1,
	I2,
	O
);
	input [31:0] I0;
	input [31:0] I1;
	input [31:0] I2;
	output wire [31:0] O;
	wire orr_inst0_out;
	wire orr_inst1_out;
	wire orr_inst10_out;
	wire orr_inst11_out;
	wire orr_inst12_out;
	wire orr_inst13_out;
	wire orr_inst14_out;
	wire orr_inst15_out;
	wire orr_inst16_out;
	wire orr_inst17_out;
	wire orr_inst18_out;
	wire orr_inst19_out;
	wire orr_inst2_out;
	wire orr_inst20_out;
	wire orr_inst21_out;
	wire orr_inst22_out;
	wire orr_inst23_out;
	wire orr_inst24_out;
	wire orr_inst25_out;
	wire orr_inst26_out;
	wire orr_inst27_out;
	wire orr_inst28_out;
	wire orr_inst29_out;
	wire orr_inst3_out;
	wire orr_inst30_out;
	wire orr_inst31_out;
	wire orr_inst4_out;
	wire orr_inst5_out;
	wire orr_inst6_out;
	wire orr_inst7_out;
	wire orr_inst8_out;
	wire orr_inst9_out;
	wire [2:0] orr_inst0_in;
	assign orr_inst0_in = {I2[0], I1[0], I0[0]};
	coreir_orr #(.width(3)) orr_inst0(
		.in(orr_inst0_in),
		.out(orr_inst0_out)
	);
	wire [2:0] orr_inst1_in;
	assign orr_inst1_in = {I2[1], I1[1], I0[1]};
	coreir_orr #(.width(3)) orr_inst1(
		.in(orr_inst1_in),
		.out(orr_inst1_out)
	);
	wire [2:0] orr_inst10_in;
	assign orr_inst10_in = {I2[10], I1[10], I0[10]};
	coreir_orr #(.width(3)) orr_inst10(
		.in(orr_inst10_in),
		.out(orr_inst10_out)
	);
	wire [2:0] orr_inst11_in;
	assign orr_inst11_in = {I2[11], I1[11], I0[11]};
	coreir_orr #(.width(3)) orr_inst11(
		.in(orr_inst11_in),
		.out(orr_inst11_out)
	);
	wire [2:0] orr_inst12_in;
	assign orr_inst12_in = {I2[12], I1[12], I0[12]};
	coreir_orr #(.width(3)) orr_inst12(
		.in(orr_inst12_in),
		.out(orr_inst12_out)
	);
	wire [2:0] orr_inst13_in;
	assign orr_inst13_in = {I2[13], I1[13], I0[13]};
	coreir_orr #(.width(3)) orr_inst13(
		.in(orr_inst13_in),
		.out(orr_inst13_out)
	);
	wire [2:0] orr_inst14_in;
	assign orr_inst14_in = {I2[14], I1[14], I0[14]};
	coreir_orr #(.width(3)) orr_inst14(
		.in(orr_inst14_in),
		.out(orr_inst14_out)
	);
	wire [2:0] orr_inst15_in;
	assign orr_inst15_in = {I2[15], I1[15], I0[15]};
	coreir_orr #(.width(3)) orr_inst15(
		.in(orr_inst15_in),
		.out(orr_inst15_out)
	);
	wire [2:0] orr_inst16_in;
	assign orr_inst16_in = {I2[16], I1[16], I0[16]};
	coreir_orr #(.width(3)) orr_inst16(
		.in(orr_inst16_in),
		.out(orr_inst16_out)
	);
	wire [2:0] orr_inst17_in;
	assign orr_inst17_in = {I2[17], I1[17], I0[17]};
	coreir_orr #(.width(3)) orr_inst17(
		.in(orr_inst17_in),
		.out(orr_inst17_out)
	);
	wire [2:0] orr_inst18_in;
	assign orr_inst18_in = {I2[18], I1[18], I0[18]};
	coreir_orr #(.width(3)) orr_inst18(
		.in(orr_inst18_in),
		.out(orr_inst18_out)
	);
	wire [2:0] orr_inst19_in;
	assign orr_inst19_in = {I2[19], I1[19], I0[19]};
	coreir_orr #(.width(3)) orr_inst19(
		.in(orr_inst19_in),
		.out(orr_inst19_out)
	);
	wire [2:0] orr_inst2_in;
	assign orr_inst2_in = {I2[2], I1[2], I0[2]};
	coreir_orr #(.width(3)) orr_inst2(
		.in(orr_inst2_in),
		.out(orr_inst2_out)
	);
	wire [2:0] orr_inst20_in;
	assign orr_inst20_in = {I2[20], I1[20], I0[20]};
	coreir_orr #(.width(3)) orr_inst20(
		.in(orr_inst20_in),
		.out(orr_inst20_out)
	);
	wire [2:0] orr_inst21_in;
	assign orr_inst21_in = {I2[21], I1[21], I0[21]};
	coreir_orr #(.width(3)) orr_inst21(
		.in(orr_inst21_in),
		.out(orr_inst21_out)
	);
	wire [2:0] orr_inst22_in;
	assign orr_inst22_in = {I2[22], I1[22], I0[22]};
	coreir_orr #(.width(3)) orr_inst22(
		.in(orr_inst22_in),
		.out(orr_inst22_out)
	);
	wire [2:0] orr_inst23_in;
	assign orr_inst23_in = {I2[23], I1[23], I0[23]};
	coreir_orr #(.width(3)) orr_inst23(
		.in(orr_inst23_in),
		.out(orr_inst23_out)
	);
	wire [2:0] orr_inst24_in;
	assign orr_inst24_in = {I2[24], I1[24], I0[24]};
	coreir_orr #(.width(3)) orr_inst24(
		.in(orr_inst24_in),
		.out(orr_inst24_out)
	);
	wire [2:0] orr_inst25_in;
	assign orr_inst25_in = {I2[25], I1[25], I0[25]};
	coreir_orr #(.width(3)) orr_inst25(
		.in(orr_inst25_in),
		.out(orr_inst25_out)
	);
	wire [2:0] orr_inst26_in;
	assign orr_inst26_in = {I2[26], I1[26], I0[26]};
	coreir_orr #(.width(3)) orr_inst26(
		.in(orr_inst26_in),
		.out(orr_inst26_out)
	);
	wire [2:0] orr_inst27_in;
	assign orr_inst27_in = {I2[27], I1[27], I0[27]};
	coreir_orr #(.width(3)) orr_inst27(
		.in(orr_inst27_in),
		.out(orr_inst27_out)
	);
	wire [2:0] orr_inst28_in;
	assign orr_inst28_in = {I2[28], I1[28], I0[28]};
	coreir_orr #(.width(3)) orr_inst28(
		.in(orr_inst28_in),
		.out(orr_inst28_out)
	);
	wire [2:0] orr_inst29_in;
	assign orr_inst29_in = {I2[29], I1[29], I0[29]};
	coreir_orr #(.width(3)) orr_inst29(
		.in(orr_inst29_in),
		.out(orr_inst29_out)
	);
	wire [2:0] orr_inst3_in;
	assign orr_inst3_in = {I2[3], I1[3], I0[3]};
	coreir_orr #(.width(3)) orr_inst3(
		.in(orr_inst3_in),
		.out(orr_inst3_out)
	);
	wire [2:0] orr_inst30_in;
	assign orr_inst30_in = {I2[30], I1[30], I0[30]};
	coreir_orr #(.width(3)) orr_inst30(
		.in(orr_inst30_in),
		.out(orr_inst30_out)
	);
	wire [2:0] orr_inst31_in;
	assign orr_inst31_in = {I2[31], I1[31], I0[31]};
	coreir_orr #(.width(3)) orr_inst31(
		.in(orr_inst31_in),
		.out(orr_inst31_out)
	);
	wire [2:0] orr_inst4_in;
	assign orr_inst4_in = {I2[4], I1[4], I0[4]};
	coreir_orr #(.width(3)) orr_inst4(
		.in(orr_inst4_in),
		.out(orr_inst4_out)
	);
	wire [2:0] orr_inst5_in;
	assign orr_inst5_in = {I2[5], I1[5], I0[5]};
	coreir_orr #(.width(3)) orr_inst5(
		.in(orr_inst5_in),
		.out(orr_inst5_out)
	);
	wire [2:0] orr_inst6_in;
	assign orr_inst6_in = {I2[6], I1[6], I0[6]};
	coreir_orr #(.width(3)) orr_inst6(
		.in(orr_inst6_in),
		.out(orr_inst6_out)
	);
	wire [2:0] orr_inst7_in;
	assign orr_inst7_in = {I2[7], I1[7], I0[7]};
	coreir_orr #(.width(3)) orr_inst7(
		.in(orr_inst7_in),
		.out(orr_inst7_out)
	);
	wire [2:0] orr_inst8_in;
	assign orr_inst8_in = {I2[8], I1[8], I0[8]};
	coreir_orr #(.width(3)) orr_inst8(
		.in(orr_inst8_in),
		.out(orr_inst8_out)
	);
	wire [2:0] orr_inst9_in;
	assign orr_inst9_in = {I2[9], I1[9], I0[9]};
	coreir_orr #(.width(3)) orr_inst9(
		.in(orr_inst9_in),
		.out(orr_inst9_out)
	);
	assign O = {orr_inst31_out, orr_inst30_out, orr_inst29_out, orr_inst28_out, orr_inst27_out, orr_inst26_out, orr_inst25_out, orr_inst24_out, orr_inst23_out, orr_inst22_out, orr_inst21_out, orr_inst20_out, orr_inst19_out, orr_inst18_out, orr_inst17_out, orr_inst16_out, orr_inst15_out, orr_inst14_out, orr_inst13_out, orr_inst12_out, orr_inst11_out, orr_inst10_out, orr_inst9_out, orr_inst8_out, orr_inst7_out, orr_inst6_out, orr_inst5_out, orr_inst4_out, orr_inst3_out, orr_inst2_out, orr_inst1_out, orr_inst0_out};
endmodule
module MuxWrapperAOI_1_1_RegularReadyValid (
	I,
	O,
	ready_in,
	ready_out,
	valid_in,
	valid_out
);
	input [0:0] I;
	output wire [0:0] O;
	input ready_in;
	output wire ready_out;
	input valid_in;
	output wire valid_out;
	assign O = I;
	assign ready_out = ready_in;
	assign valid_out = valid_in;
endmodule
module MuxWrapperAOI_1_1_ConstReadyValid (
	I,
	O,
	ready_in,
	ready_out,
	valid_in,
	valid_out
);
	input [0:0] I;
	output wire [0:0] O;
	input ready_in;
	output wire ready_out;
	input valid_in;
	output wire valid_out;
	assign O = I;
	assign ready_out = ready_in;
	assign valid_out = valid_in;
endmodule
module MuxWrapperAOI_1_17_RegularReadyValid (
	I,
	O,
	ready_in,
	ready_out,
	valid_in,
	valid_out
);
	input [16:0] I;
	output wire [16:0] O;
	input ready_in;
	output wire ready_out;
	input valid_in;
	output wire valid_out;
	assign O = I;
	assign ready_out = ready_in;
	assign valid_out = valid_in;
endmodule
module MuxWrapperAOI_1_17_ConstReadyValid (
	I,
	O,
	ready_in,
	ready_out,
	valid_in,
	valid_out
);
	input [16:0] I;
	output wire [16:0] O;
	input ready_in;
	output wire ready_out;
	input valid_in;
	output wire valid_out;
	assign O = I;
	assign ready_out = ready_in;
	assign valid_out = valid_in;
endmodule
module MuxWithDefaultWrapper_6_32_8_0 (
	I,
	S,
	EN,
	O
);
	input [191:0] I;
	input [7:0] S;
	input [0:0] EN;
	output wire [31:0] O;
	wire [31:0] const_0_32_out;
	wire [7:0] const_6_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_ult_inst0_out;
	wire [31:0] mux_aoi_2_32_inst0_O;
	wire [1:0] mux_aoi_2_32_inst0_out_sel;
	wire [31:0] mux_aoi_6_32_inst0_O;
	wire [7:0] mux_aoi_6_32_inst0_out_sel;
	coreir_const #(
		.value(32'h00000000),
		.width(32)
	) const_0_32(.out(const_0_32_out));
	coreir_const #(
		.value(8'h06),
		.width(8)
	) const_6_8(.out(const_6_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_ult_inst0_out),
		.in1(EN[0]),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_ult #(.width(8)) magma_Bits_8_ult_inst0(
		.in0(S),
		.in1(const_6_8_out),
		.out(magma_Bits_8_ult_inst0_out)
	);
	wire [63:0] mux_aoi_2_32_inst0_I;
	assign mux_aoi_2_32_inst0_I[32+:32] = mux_aoi_6_32_inst0_O;
	assign mux_aoi_2_32_inst0_I[0+:32] = const_0_32_out;
	mux_aoi_2_32 mux_aoi_2_32_inst0(
		.I(mux_aoi_2_32_inst0_I),
		.O(mux_aoi_2_32_inst0_O),
		.S(magma_Bit_and_inst0_out),
		.out_sel(mux_aoi_2_32_inst0_out_sel)
	);
	wire [191:0] mux_aoi_6_32_inst0_I;
	assign mux_aoi_6_32_inst0_I[160+:32] = I[160+:32];
	assign mux_aoi_6_32_inst0_I[128+:32] = I[128+:32];
	assign mux_aoi_6_32_inst0_I[96+:32] = I[96+:32];
	assign mux_aoi_6_32_inst0_I[64+:32] = I[64+:32];
	assign mux_aoi_6_32_inst0_I[32+:32] = I[32+:32];
	assign mux_aoi_6_32_inst0_I[0+:32] = I[0+:32];
	mux_aoi_6_32 mux_aoi_6_32_inst0(
		.I(mux_aoi_6_32_inst0_I),
		.O(mux_aoi_6_32_inst0_O),
		.S(S[2:0]),
		.out_sel(mux_aoi_6_32_inst0_out_sel)
	);
	assign O = mux_aoi_2_32_inst0_O;
endmodule
module MuxWithDefaultWrapper_16_32_8_0 (
	I,
	S,
	EN,
	O
);
	input [511:0] I;
	input [7:0] S;
	input [0:0] EN;
	output wire [31:0] O;
	wire [31:0] const_0_32_out;
	wire [7:0] const_16_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_ult_inst0_out;
	wire [31:0] mux_aoi_16_32_inst0_O;
	wire [15:0] mux_aoi_16_32_inst0_out_sel;
	wire [31:0] mux_aoi_2_32_inst0_O;
	wire [1:0] mux_aoi_2_32_inst0_out_sel;
	coreir_const #(
		.value(32'h00000000),
		.width(32)
	) const_0_32(.out(const_0_32_out));
	coreir_const #(
		.value(8'h10),
		.width(8)
	) const_16_8(.out(const_16_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_ult_inst0_out),
		.in1(EN[0]),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_ult #(.width(8)) magma_Bits_8_ult_inst0(
		.in0(S),
		.in1(const_16_8_out),
		.out(magma_Bits_8_ult_inst0_out)
	);
	wire [511:0] mux_aoi_16_32_inst0_I;
	assign mux_aoi_16_32_inst0_I[480+:32] = I[480+:32];
	assign mux_aoi_16_32_inst0_I[448+:32] = I[448+:32];
	assign mux_aoi_16_32_inst0_I[416+:32] = I[416+:32];
	assign mux_aoi_16_32_inst0_I[384+:32] = I[384+:32];
	assign mux_aoi_16_32_inst0_I[352+:32] = I[352+:32];
	assign mux_aoi_16_32_inst0_I[320+:32] = I[320+:32];
	assign mux_aoi_16_32_inst0_I[288+:32] = I[288+:32];
	assign mux_aoi_16_32_inst0_I[256+:32] = I[256+:32];
	assign mux_aoi_16_32_inst0_I[224+:32] = I[224+:32];
	assign mux_aoi_16_32_inst0_I[192+:32] = I[192+:32];
	assign mux_aoi_16_32_inst0_I[160+:32] = I[160+:32];
	assign mux_aoi_16_32_inst0_I[128+:32] = I[128+:32];
	assign mux_aoi_16_32_inst0_I[96+:32] = I[96+:32];
	assign mux_aoi_16_32_inst0_I[64+:32] = I[64+:32];
	assign mux_aoi_16_32_inst0_I[32+:32] = I[32+:32];
	assign mux_aoi_16_32_inst0_I[0+:32] = I[0+:32];
	mux_aoi_16_32 mux_aoi_16_32_inst0(
		.I(mux_aoi_16_32_inst0_I),
		.O(mux_aoi_16_32_inst0_O),
		.S(S[3:0]),
		.out_sel(mux_aoi_16_32_inst0_out_sel)
	);
	wire [63:0] mux_aoi_2_32_inst0_I;
	assign mux_aoi_2_32_inst0_I[32+:32] = mux_aoi_16_32_inst0_O;
	assign mux_aoi_2_32_inst0_I[0+:32] = const_0_32_out;
	mux_aoi_2_32 mux_aoi_2_32_inst0(
		.I(mux_aoi_2_32_inst0_I),
		.O(mux_aoi_2_32_inst0_O),
		.S(magma_Bit_and_inst0_out),
		.out_sel(mux_aoi_2_32_inst0_out_sel)
	);
	assign O = mux_aoi_2_32_inst0_O;
endmodule
module MuxWithDefaultWrapper_13_32_8_0 (
	I,
	S,
	EN,
	O
);
	input [415:0] I;
	input [7:0] S;
	input [0:0] EN;
	output wire [31:0] O;
	wire [31:0] const_0_32_out;
	wire [7:0] const_13_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_ult_inst0_out;
	wire [31:0] mux_aoi_13_32_inst0_O;
	wire [15:0] mux_aoi_13_32_inst0_out_sel;
	wire [31:0] mux_aoi_2_32_inst0_O;
	wire [1:0] mux_aoi_2_32_inst0_out_sel;
	coreir_const #(
		.value(32'h00000000),
		.width(32)
	) const_0_32(.out(const_0_32_out));
	coreir_const #(
		.value(8'h0d),
		.width(8)
	) const_13_8(.out(const_13_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_ult_inst0_out),
		.in1(EN[0]),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_ult #(.width(8)) magma_Bits_8_ult_inst0(
		.in0(S),
		.in1(const_13_8_out),
		.out(magma_Bits_8_ult_inst0_out)
	);
	wire [415:0] mux_aoi_13_32_inst0_I;
	assign mux_aoi_13_32_inst0_I[384+:32] = I[384+:32];
	assign mux_aoi_13_32_inst0_I[352+:32] = I[352+:32];
	assign mux_aoi_13_32_inst0_I[320+:32] = I[320+:32];
	assign mux_aoi_13_32_inst0_I[288+:32] = I[288+:32];
	assign mux_aoi_13_32_inst0_I[256+:32] = I[256+:32];
	assign mux_aoi_13_32_inst0_I[224+:32] = I[224+:32];
	assign mux_aoi_13_32_inst0_I[192+:32] = I[192+:32];
	assign mux_aoi_13_32_inst0_I[160+:32] = I[160+:32];
	assign mux_aoi_13_32_inst0_I[128+:32] = I[128+:32];
	assign mux_aoi_13_32_inst0_I[96+:32] = I[96+:32];
	assign mux_aoi_13_32_inst0_I[64+:32] = I[64+:32];
	assign mux_aoi_13_32_inst0_I[32+:32] = I[32+:32];
	assign mux_aoi_13_32_inst0_I[0+:32] = I[0+:32];
	mux_aoi_13_32 mux_aoi_13_32_inst0(
		.I(mux_aoi_13_32_inst0_I),
		.O(mux_aoi_13_32_inst0_O),
		.S(S[3:0]),
		.out_sel(mux_aoi_13_32_inst0_out_sel)
	);
	wire [63:0] mux_aoi_2_32_inst0_I;
	assign mux_aoi_2_32_inst0_I[32+:32] = mux_aoi_13_32_inst0_O;
	assign mux_aoi_2_32_inst0_I[0+:32] = const_0_32_out;
	mux_aoi_2_32 mux_aoi_2_32_inst0(
		.I(mux_aoi_2_32_inst0_I),
		.O(mux_aoi_2_32_inst0_O),
		.S(magma_Bit_and_inst0_out),
		.out_sel(mux_aoi_2_32_inst0_out_sel)
	);
	assign O = mux_aoi_2_32_inst0_O;
endmodule
module Chain_2_16 (
	accessor_output,
	chain_data_in,
	chain_en,
	clk_en,
	curr_tile_data_out,
	flush,
	data_out_tile
);
	input wire [1:0] accessor_output;
	input wire [31:0] chain_data_in;
	input wire chain_en;
	input wire clk_en;
	input wire [31:0] curr_tile_data_out;
	input wire flush;
	output reg [31:0] data_out_tile;
	always @(*) begin
		if (accessor_output[0])
			data_out_tile[0+:16] = curr_tile_data_out[0+:16];
		else if (chain_en)
			data_out_tile[0+:16] = chain_data_in[0+:16];
		else
			data_out_tile[0+:16] = 16'h0000;
		if (accessor_output[1])
			data_out_tile[16+:16] = curr_tile_data_out[16+:16];
		else if (chain_en)
			data_out_tile[16+:16] = chain_data_in[16+:16];
		else
			data_out_tile[16+:16] = 16'h0000;
	end
endmodule
module MemCore_inner (
	CONFIG_SPACE_0,
	CONFIG_SPACE_1,
	CONFIG_SPACE_10,
	CONFIG_SPACE_11,
	CONFIG_SPACE_12,
	CONFIG_SPACE_13,
	CONFIG_SPACE_14,
	CONFIG_SPACE_15,
	CONFIG_SPACE_16,
	CONFIG_SPACE_17,
	CONFIG_SPACE_18,
	CONFIG_SPACE_19,
	CONFIG_SPACE_2,
	CONFIG_SPACE_20,
	CONFIG_SPACE_21,
	CONFIG_SPACE_22,
	CONFIG_SPACE_23,
	CONFIG_SPACE_24,
	CONFIG_SPACE_25,
	CONFIG_SPACE_26,
	CONFIG_SPACE_27,
	CONFIG_SPACE_28,
	CONFIG_SPACE_29,
	CONFIG_SPACE_3,
	CONFIG_SPACE_30,
	CONFIG_SPACE_31,
	CONFIG_SPACE_32,
	CONFIG_SPACE_33,
	CONFIG_SPACE_34,
	CONFIG_SPACE_35,
	CONFIG_SPACE_36,
	CONFIG_SPACE_37,
	CONFIG_SPACE_38,
	CONFIG_SPACE_39,
	CONFIG_SPACE_4,
	CONFIG_SPACE_40,
	CONFIG_SPACE_41,
	CONFIG_SPACE_42,
	CONFIG_SPACE_43,
	CONFIG_SPACE_44,
	CONFIG_SPACE_45,
	CONFIG_SPACE_5,
	CONFIG_SPACE_6,
	CONFIG_SPACE_7,
	CONFIG_SPACE_8,
	CONFIG_SPACE_9,
	MEM_input_width_17_num_0,
	MEM_input_width_17_num_0_valid,
	MEM_input_width_17_num_1,
	MEM_input_width_17_num_1_valid,
	MEM_input_width_17_num_2,
	MEM_input_width_17_num_2_valid,
	MEM_input_width_17_num_3,
	MEM_input_width_17_num_3_valid,
	MEM_input_width_1_num_0,
	MEM_input_width_1_num_1,
	MEM_output_width_17_num_0_ready,
	MEM_output_width_17_num_1_ready,
	MEM_output_width_17_num_2_ready,
	clk,
	clk_en,
	config_addr_in,
	config_data_in,
	config_en,
	config_read,
	config_write,
	flush,
	mode,
	mode_excl,
	rst_n,
	tile_en,
	MEM_input_width_17_num_0_ready,
	MEM_input_width_17_num_1_ready,
	MEM_input_width_17_num_2_ready,
	MEM_input_width_17_num_3_ready,
	MEM_output_width_17_num_0,
	MEM_output_width_17_num_0_valid,
	MEM_output_width_17_num_1,
	MEM_output_width_17_num_1_valid,
	MEM_output_width_17_num_2,
	MEM_output_width_17_num_2_valid,
	MEM_output_width_1_num_0,
	MEM_output_width_1_num_1,
	MEM_output_width_1_num_2,
	config_data_out
);
	input wire [31:0] CONFIG_SPACE_0;
	input wire [31:0] CONFIG_SPACE_1;
	input wire [31:0] CONFIG_SPACE_10;
	input wire [31:0] CONFIG_SPACE_11;
	input wire [31:0] CONFIG_SPACE_12;
	input wire [31:0] CONFIG_SPACE_13;
	input wire [31:0] CONFIG_SPACE_14;
	input wire [31:0] CONFIG_SPACE_15;
	input wire [31:0] CONFIG_SPACE_16;
	input wire [31:0] CONFIG_SPACE_17;
	input wire [31:0] CONFIG_SPACE_18;
	input wire [31:0] CONFIG_SPACE_19;
	input wire [31:0] CONFIG_SPACE_2;
	input wire [31:0] CONFIG_SPACE_20;
	input wire [31:0] CONFIG_SPACE_21;
	input wire [31:0] CONFIG_SPACE_22;
	input wire [31:0] CONFIG_SPACE_23;
	input wire [31:0] CONFIG_SPACE_24;
	input wire [31:0] CONFIG_SPACE_25;
	input wire [31:0] CONFIG_SPACE_26;
	input wire [31:0] CONFIG_SPACE_27;
	input wire [31:0] CONFIG_SPACE_28;
	input wire [31:0] CONFIG_SPACE_29;
	input wire [31:0] CONFIG_SPACE_3;
	input wire [31:0] CONFIG_SPACE_30;
	input wire [31:0] CONFIG_SPACE_31;
	input wire [31:0] CONFIG_SPACE_32;
	input wire [31:0] CONFIG_SPACE_33;
	input wire [31:0] CONFIG_SPACE_34;
	input wire [31:0] CONFIG_SPACE_35;
	input wire [31:0] CONFIG_SPACE_36;
	input wire [31:0] CONFIG_SPACE_37;
	input wire [31:0] CONFIG_SPACE_38;
	input wire [31:0] CONFIG_SPACE_39;
	input wire [31:0] CONFIG_SPACE_4;
	input wire [31:0] CONFIG_SPACE_40;
	input wire [31:0] CONFIG_SPACE_41;
	input wire [31:0] CONFIG_SPACE_42;
	input wire [31:0] CONFIG_SPACE_43;
	input wire [31:0] CONFIG_SPACE_44;
	input wire [18:0] CONFIG_SPACE_45;
	input wire [31:0] CONFIG_SPACE_5;
	input wire [31:0] CONFIG_SPACE_6;
	input wire [31:0] CONFIG_SPACE_7;
	input wire [31:0] CONFIG_SPACE_8;
	input wire [31:0] CONFIG_SPACE_9;
	input wire [16:0] MEM_input_width_17_num_0;
	input wire MEM_input_width_17_num_0_valid;
	input wire [16:0] MEM_input_width_17_num_1;
	input wire MEM_input_width_17_num_1_valid;
	input wire [16:0] MEM_input_width_17_num_2;
	input wire MEM_input_width_17_num_2_valid;
	input wire [16:0] MEM_input_width_17_num_3;
	input wire MEM_input_width_17_num_3_valid;
	input wire MEM_input_width_1_num_0;
	input wire MEM_input_width_1_num_1;
	input wire MEM_output_width_17_num_0_ready;
	input wire MEM_output_width_17_num_1_ready;
	input wire MEM_output_width_17_num_2_ready;
	input wire clk;
	input wire clk_en;
	input wire [7:0] config_addr_in;
	input wire [31:0] config_data_in;
	input wire [1:0] config_en;
	input wire config_read;
	input wire config_write;
	input wire flush;
	input wire [1:0] mode;
	input wire mode_excl;
	input wire rst_n;
	input wire tile_en;
	output reg MEM_input_width_17_num_0_ready;
	output reg MEM_input_width_17_num_1_ready;
	output reg MEM_input_width_17_num_2_ready;
	output reg MEM_input_width_17_num_3_ready;
	output reg [16:0] MEM_output_width_17_num_0;
	output reg MEM_output_width_17_num_0_valid;
	output reg [16:0] MEM_output_width_17_num_1;
	output reg MEM_output_width_17_num_1_valid;
	output reg [16:0] MEM_output_width_17_num_2;
	output reg MEM_output_width_17_num_2_valid;
	output reg MEM_output_width_1_num_0;
	output reg MEM_output_width_1_num_1;
	output reg MEM_output_width_1_num_2;
	output wire [63:0] config_data_out;
	wire [1458:0] CONFIG_SPACE;
	wire [15:0] config_data_in_shrt;
	wire [31:0] config_data_out_shrt;
	wire [8:0] config_seq_addr_out;
	wire config_seq_clk_en;
	reg [63:0] config_seq_rd_data_stg;
	wire config_seq_ren_out;
	wire config_seq_wen_out;
	wire [63:0] config_seq_wr_data;
	wire gclk;
	wire [16:0] input_width_17_num_0_fifo_out;
	reg input_width_17_num_0_fifo_out_ready;
	wire input_width_17_num_0_fifo_out_valid;
	wire input_width_17_num_0_input_fifo_empty;
	wire input_width_17_num_0_input_fifo_full;
	wire [16:0] input_width_17_num_1_fifo_out;
	reg input_width_17_num_1_fifo_out_ready;
	wire input_width_17_num_1_fifo_out_valid;
	wire input_width_17_num_1_input_fifo_empty;
	wire input_width_17_num_1_input_fifo_full;
	wire [16:0] input_width_17_num_2_fifo_out;
	reg input_width_17_num_2_fifo_out_ready;
	wire input_width_17_num_2_fifo_out_valid;
	wire input_width_17_num_2_input_fifo_empty;
	wire input_width_17_num_2_input_fifo_full;
	wire [16:0] input_width_17_num_3_fifo_out;
	reg input_width_17_num_3_fifo_out_ready;
	wire input_width_17_num_3_fifo_out_valid;
	wire input_width_17_num_3_input_fifo_empty;
	wire input_width_17_num_3_input_fifo_full;
	wire mem_ctrl_fiber_access_16_flat_clk;
	wire [8:0] mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_addr_to_mem_lifted_lifted;
	wire [3:0] mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_buffet_capacity_log_0;
	wire [3:0] mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_buffet_capacity_log_1;
	reg [63:0] mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_data_from_mem_lifted_lifted;
	wire [63:0] mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_data_to_mem_lifted_lifted;
	wire mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_ren_to_mem_lifted_lifted;
	wire mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_tile_en;
	wire mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_wen_to_mem_lifted_lifted;
	wire mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_block_mode;
	wire mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_dense;
	wire [15:0] mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_dim_size;
	wire mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_do_repeat;
	wire [15:0] mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_inner_dim_offset;
	wire mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_lookup;
	wire [15:0] mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_repeat_factor;
	wire mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_repeat_outer_inner_n;
	wire mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_root;
	wire mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_spacc_mode;
	wire [15:0] mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_stop_lvl;
	wire mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_tile_en;
	wire mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_tile_en;
	wire mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_block_mode;
	wire mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_compressed;
	wire mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_init_blank;
	wire mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_lowest_level;
	wire mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_spacc_mode;
	wire [15:0] mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_stop_lvl;
	wire mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_tile_en;
	wire [16:0] mem_ctrl_fiber_access_16_flat_read_scanner_block_rd_out_f_;
	wire mem_ctrl_fiber_access_16_flat_read_scanner_block_rd_out_valid_f_;
	wire [16:0] mem_ctrl_fiber_access_16_flat_read_scanner_coord_out_f_;
	wire mem_ctrl_fiber_access_16_flat_read_scanner_coord_out_valid_f_;
	wire [16:0] mem_ctrl_fiber_access_16_flat_read_scanner_pos_out_f_;
	wire mem_ctrl_fiber_access_16_flat_read_scanner_pos_out_valid_f_;
	wire mem_ctrl_fiber_access_16_flat_read_scanner_us_pos_in_ready_f_;
	wire mem_ctrl_fiber_access_16_flat_write_scanner_addr_in_ready_f_;
	wire mem_ctrl_fiber_access_16_flat_write_scanner_block_wr_in_ready_f_;
	wire mem_ctrl_fiber_access_16_flat_write_scanner_data_in_ready_f_;
	wire mem_ctrl_stencil_valid_flat_clk;
	wire mem_ctrl_stencil_valid_flat_stencil_valid_f_;
	wire [3:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality;
	wire [10:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_0;
	wire [10:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_1;
	wire [10:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_2;
	wire [10:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_3;
	wire [10:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_4;
	wire [10:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_5;
	wire mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable;
	wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr;
	wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0;
	wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1;
	wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2;
	wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3;
	wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4;
	wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5;
	wire mem_ctrl_strg_ram_64_512_delay1_flat_clk;
	wire [16:0] mem_ctrl_strg_ram_64_512_delay1_flat_data_out_f_;
	wire mem_ctrl_strg_ram_64_512_delay1_flat_ready_f_;
	wire [8:0] mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_addr_out_lifted;
	reg [63:0] mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_data_from_strg_lifted;
	wire [63:0] mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_data_to_strg_lifted;
	wire mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_ren_to_strg_lifted;
	wire mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_wen_to_strg_lifted;
	wire mem_ctrl_strg_ram_64_512_delay1_flat_valid_out_f_;
	wire mem_ctrl_strg_ub_vec_flat_accessor_output_f_b_0;
	wire mem_ctrl_strg_ub_vec_flat_accessor_output_f_b_1;
	wire mem_ctrl_strg_ub_vec_flat_clk;
	wire [16:0] mem_ctrl_strg_ub_vec_flat_data_out_f_0;
	wire [16:0] mem_ctrl_strg_ub_vec_flat_data_out_f_1;
	wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_addr_out_lifted;
	wire [2:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr;
	wire [2:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0;
	wire [2:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1;
	wire [2:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2;
	wire [2:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr;
	wire [2:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0;
	wire [2:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1;
	wire [2:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2;
	wire mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2;
	wire mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2;
	wire [2:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2;
	wire [2:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_agg_read_padding;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_agg_read_padding;
	wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_sram_shared_addr_gen_0_starting_addr;
	wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_sram_shared_addr_gen_1_starting_addr;
	wire [1:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_mode_0;
	wire [1:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_mode_1;
	wire mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en;
	reg [63:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_data_from_strg_lifted;
	wire [63:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_data_to_strg_lifted;
	wire mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_ren_to_strg_lifted;
	wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr;
	wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0;
	wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1;
	wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2;
	wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3;
	wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4;
	wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5;
	wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr;
	wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0;
	wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1;
	wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2;
	wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3;
	wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4;
	wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5;
	wire mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable;
	wire [9:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_delay;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5;
	wire mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable;
	wire [9:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_delay;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4;
	wire [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5;
	wire mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_shared_tb_0;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5;
	wire mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable;
	wire [9:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_delay;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5;
	wire mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable;
	wire [9:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_delay;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5;
	wire mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_wen_to_strg_lifted;
	wire memory_0_clk_en;
	reg [63:0] memory_0_data_in_p0;
	wire [63:0] memory_0_data_out_p0;
	reg [8:0] memory_0_read_addr_p0;
	reg memory_0_read_enable_p0;
	reg [8:0] memory_0_write_addr_p0;
	reg memory_0_write_enable_p0;
	reg [16:0] output_width_17_num_0_fifo_in;
	wire output_width_17_num_0_fifo_in_ready;
	reg output_width_17_num_0_fifo_in_valid;
	wire [16:0] output_width_17_num_0_output_fifo_data_out;
	wire output_width_17_num_0_output_fifo_empty;
	wire output_width_17_num_0_output_fifo_full;
	reg [16:0] output_width_17_num_1_fifo_in;
	wire output_width_17_num_1_fifo_in_ready;
	reg output_width_17_num_1_fifo_in_valid;
	wire [16:0] output_width_17_num_1_output_fifo_data_out;
	wire output_width_17_num_1_output_fifo_empty;
	wire output_width_17_num_1_output_fifo_full;
	reg [16:0] output_width_17_num_2_fifo_in;
	wire output_width_17_num_2_fifo_in_ready;
	reg output_width_17_num_2_fifo_in_valid;
	wire [16:0] output_width_17_num_2_output_fifo_data_out;
	wire output_width_17_num_2_output_fifo_empty;
	wire output_width_17_num_2_output_fifo_full;
	assign gclk = clk & tile_en;
	assign mem_ctrl_fiber_access_16_flat_clk = gclk & (mode == 2'h0);
	assign mem_ctrl_strg_ub_vec_flat_clk = gclk & (mode == 2'h1);
	assign mem_ctrl_strg_ram_64_512_delay1_flat_clk = gclk & (mode == 2'h2);
	assign mem_ctrl_stencil_valid_flat_clk = gclk;
	assign input_width_17_num_0_fifo_out_valid = ~input_width_17_num_0_input_fifo_empty;
	always @(*) begin
		input_width_17_num_0_fifo_out_ready = 1'h1;
		if (mode == 2'h0)
			input_width_17_num_0_fifo_out_ready = mem_ctrl_fiber_access_16_flat_read_scanner_us_pos_in_ready_f_;
		else
			input_width_17_num_0_fifo_out_ready = 1'h1;
	end
	always @(*) begin
		MEM_input_width_17_num_0_ready = 1'h1;
		if (mode == 2'h0)
			MEM_input_width_17_num_0_ready = ~input_width_17_num_0_input_fifo_full;
		else if (mode == 2'h1)
			MEM_input_width_17_num_0_ready = 1'h1;
		else if (mode == 2'h2)
			MEM_input_width_17_num_0_ready = 1'h1;
	end
	assign input_width_17_num_1_fifo_out_valid = ~input_width_17_num_1_input_fifo_empty;
	always @(*) begin
		input_width_17_num_1_fifo_out_ready = 1'h1;
		if (mode == 2'h0)
			input_width_17_num_1_fifo_out_ready = mem_ctrl_fiber_access_16_flat_write_scanner_addr_in_ready_f_;
		else
			input_width_17_num_1_fifo_out_ready = 1'h1;
	end
	always @(*) begin
		MEM_input_width_17_num_1_ready = 1'h1;
		if (mode == 2'h0)
			MEM_input_width_17_num_1_ready = ~input_width_17_num_1_input_fifo_full;
		else if (mode == 2'h1)
			MEM_input_width_17_num_1_ready = 1'h1;
		else if (mode == 2'h2)
			MEM_input_width_17_num_1_ready = 1'h1;
	end
	assign input_width_17_num_2_fifo_out_valid = ~input_width_17_num_2_input_fifo_empty;
	always @(*) begin
		input_width_17_num_2_fifo_out_ready = 1'h1;
		if (mode == 2'h0)
			input_width_17_num_2_fifo_out_ready = mem_ctrl_fiber_access_16_flat_write_scanner_block_wr_in_ready_f_;
		else
			input_width_17_num_2_fifo_out_ready = 1'h1;
	end
	always @(*) begin
		MEM_input_width_17_num_2_ready = 1'h1;
		if (mode == 2'h0)
			MEM_input_width_17_num_2_ready = ~input_width_17_num_2_input_fifo_full;
		else if (mode == 2'h1)
			MEM_input_width_17_num_2_ready = 1'h1;
		else if (mode == 2'h2)
			MEM_input_width_17_num_2_ready = 1'h1;
	end
	assign input_width_17_num_3_fifo_out_valid = ~input_width_17_num_3_input_fifo_empty;
	always @(*) begin
		input_width_17_num_3_fifo_out_ready = 1'h1;
		if (mode == 2'h0)
			input_width_17_num_3_fifo_out_ready = mem_ctrl_fiber_access_16_flat_write_scanner_data_in_ready_f_;
		else
			input_width_17_num_3_fifo_out_ready = 1'h1;
	end
	always @(*) begin
		MEM_input_width_17_num_3_ready = 1'h1;
		if (mode == 2'h0)
			MEM_input_width_17_num_3_ready = ~input_width_17_num_3_input_fifo_full;
		else if (mode == 2'h1)
			MEM_input_width_17_num_3_ready = 1'h1;
	end
	assign output_width_17_num_0_fifo_in_ready = ~output_width_17_num_0_output_fifo_full;
	always @(*) begin
		output_width_17_num_0_fifo_in = 17'h00000;
		output_width_17_num_0_fifo_in_valid = 1'h0;
		output_width_17_num_0_fifo_in = mem_ctrl_fiber_access_16_flat_read_scanner_block_rd_out_f_;
		output_width_17_num_0_fifo_in_valid = mem_ctrl_fiber_access_16_flat_read_scanner_block_rd_out_valid_f_;
	end
	always @(*) begin
		MEM_output_width_17_num_0 = 17'h00000;
		if (mode == 2'h0)
			MEM_output_width_17_num_0 = output_width_17_num_0_output_fifo_data_out;
		else if (mode == 2'h1)
			MEM_output_width_17_num_0 = mem_ctrl_strg_ub_vec_flat_data_out_f_0;
		else if (mode == 2'h2)
			MEM_output_width_17_num_0 = mem_ctrl_strg_ram_64_512_delay1_flat_data_out_f_;
	end
	always @(*) begin
		MEM_output_width_17_num_0_valid = 1'h0;
		if (mode == 2'h0)
			MEM_output_width_17_num_0_valid = ~output_width_17_num_0_output_fifo_empty;
		else if (mode == 2'h1)
			MEM_output_width_17_num_0_valid = 1'h1;
		else if (mode == 2'h2)
			MEM_output_width_17_num_0_valid = 1'h1;
	end
	assign output_width_17_num_1_fifo_in_ready = ~output_width_17_num_1_output_fifo_full;
	always @(*) begin
		output_width_17_num_1_fifo_in = 17'h00000;
		output_width_17_num_1_fifo_in_valid = 1'h0;
		output_width_17_num_1_fifo_in = mem_ctrl_fiber_access_16_flat_read_scanner_coord_out_f_;
		output_width_17_num_1_fifo_in_valid = mem_ctrl_fiber_access_16_flat_read_scanner_coord_out_valid_f_;
	end
	always @(*) begin
		MEM_output_width_17_num_1 = 17'h00000;
		if (mode == 2'h0)
			MEM_output_width_17_num_1 = output_width_17_num_1_output_fifo_data_out;
		else if (mode == 2'h1)
			MEM_output_width_17_num_1 = mem_ctrl_strg_ub_vec_flat_data_out_f_1;
	end
	always @(*) begin
		MEM_output_width_17_num_1_valid = 1'h0;
		if (mode == 2'h0)
			MEM_output_width_17_num_1_valid = ~output_width_17_num_1_output_fifo_empty;
		else if (mode == 2'h1)
			MEM_output_width_17_num_1_valid = 1'h1;
	end
	assign output_width_17_num_2_fifo_in_ready = ~output_width_17_num_2_output_fifo_full;
	always @(*) begin
		output_width_17_num_2_fifo_in = 17'h00000;
		output_width_17_num_2_fifo_in_valid = 1'h0;
		output_width_17_num_2_fifo_in = mem_ctrl_fiber_access_16_flat_read_scanner_pos_out_f_;
		output_width_17_num_2_fifo_in_valid = mem_ctrl_fiber_access_16_flat_read_scanner_pos_out_valid_f_;
	end
	always @(*) begin
		MEM_output_width_17_num_2 = 17'h00000;
		if (mode == 2'h0)
			MEM_output_width_17_num_2 = output_width_17_num_2_output_fifo_data_out;
		else
			MEM_output_width_17_num_2 = 17'h00000;
	end
	always @(*) begin
		MEM_output_width_17_num_2_valid = 1'h0;
		if (mode == 2'h0)
			MEM_output_width_17_num_2_valid = ~output_width_17_num_2_output_fifo_empty;
		else
			MEM_output_width_17_num_2_valid = 1'h0;
	end
	always @(*) begin
		MEM_output_width_1_num_0 = 1'h0;
		if (mode == 2'h1)
			MEM_output_width_1_num_0 = mem_ctrl_strg_ub_vec_flat_accessor_output_f_b_0;
		else if (mode == 2'h2)
			MEM_output_width_1_num_0 = mem_ctrl_strg_ram_64_512_delay1_flat_ready_f_;
	end
	always @(*) begin
		MEM_output_width_1_num_1 = 1'h0;
		if (mode == 2'h1)
			MEM_output_width_1_num_1 = mem_ctrl_strg_ub_vec_flat_accessor_output_f_b_1;
		else if (mode == 2'h2)
			MEM_output_width_1_num_1 = mem_ctrl_strg_ram_64_512_delay1_flat_valid_out_f_;
	end
	always @(*) begin
		MEM_output_width_1_num_2 = 1'h0;
		if (mode_excl == 1'h1)
			MEM_output_width_1_num_2 = mem_ctrl_stencil_valid_flat_stencil_valid_f_;
		else
			MEM_output_width_1_num_2 = 1'h0;
	end
	always @(*) begin
		memory_0_data_in_p0 = 64'h0000000000000000;
		memory_0_write_addr_p0 = 9'h000;
		memory_0_write_enable_p0 = 1'h0;
		memory_0_read_addr_p0 = 9'h000;
		memory_0_read_enable_p0 = 1'h0;
		if (|config_en) begin
			memory_0_data_in_p0 = config_seq_wr_data;
			memory_0_write_addr_p0 = config_seq_addr_out;
			memory_0_write_enable_p0 = config_seq_wen_out;
			memory_0_read_addr_p0 = config_seq_addr_out;
			memory_0_read_enable_p0 = config_seq_ren_out;
		end
		else if (mode == 2'h0) begin
			memory_0_data_in_p0 = mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_data_to_mem_lifted_lifted;
			memory_0_write_addr_p0 = mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_addr_to_mem_lifted_lifted;
			memory_0_write_enable_p0 = mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_wen_to_mem_lifted_lifted;
			memory_0_read_addr_p0 = mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_addr_to_mem_lifted_lifted;
			memory_0_read_enable_p0 = mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_ren_to_mem_lifted_lifted;
		end
		else if (mode == 2'h1) begin
			memory_0_data_in_p0 = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_data_to_strg_lifted;
			memory_0_write_addr_p0 = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_addr_out_lifted;
			memory_0_write_enable_p0 = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_wen_to_strg_lifted;
			memory_0_read_addr_p0 = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_addr_out_lifted;
			memory_0_read_enable_p0 = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_ren_to_strg_lifted;
		end
		else if (mode == 2'h2) begin
			memory_0_data_in_p0 = mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_data_to_strg_lifted;
			memory_0_write_addr_p0 = mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_addr_out_lifted;
			memory_0_write_enable_p0 = mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_wen_to_strg_lifted;
			memory_0_read_addr_p0 = mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_addr_out_lifted;
			memory_0_read_enable_p0 = mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_ren_to_strg_lifted;
		end
	end
	always @(*) begin
		mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_data_from_mem_lifted_lifted = memory_0_data_out_p0;
		mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_data_from_strg_lifted = memory_0_data_out_p0;
		mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_data_from_strg_lifted = memory_0_data_out_p0;
		config_seq_rd_data_stg = memory_0_data_out_p0;
	end
	assign config_data_in_shrt = config_data_in[15:0];
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	assign config_data_out[0+:32] = sv2v_cast_32(config_data_out_shrt[0+:16]);
	assign config_data_out[32+:32] = sv2v_cast_32(config_data_out_shrt[16+:16]);
	assign config_seq_clk_en = clk_en | |config_en;
	assign memory_0_clk_en = clk_en | |config_en;
	assign {mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_buffet_capacity_log_0, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_buffet_capacity_log_1, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_tile_en, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_block_mode, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_dense, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_dim_size, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_do_repeat, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_inner_dim_offset, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_lookup, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_repeat_factor, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_repeat_outer_inner_n, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_root, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_spacc_mode, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_stop_lvl, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_tile_en, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_tile_en, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_block_mode, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_compressed, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_init_blank, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_lowest_level, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_spacc_mode, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_stop_lvl, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_tile_en} = CONFIG_SPACE[103:0];
	assign {mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_agg_read_padding, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_agg_read_padding, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_sram_shared_addr_gen_0_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_sram_shared_addr_gen_1_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_mode_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_mode_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_delay, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_delay, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_shared_tb_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_delay, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_delay, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5} = CONFIG_SPACE[1275:0];
	assign {mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality, mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_0, mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_1, mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_2, mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_3, mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_4, mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_5, mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable, mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr, mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0, mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1, mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2, mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3, mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4, mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5} = CONFIG_SPACE[1458:1276];
	assign CONFIG_SPACE[31:0] = CONFIG_SPACE_0;
	assign CONFIG_SPACE[63:32] = CONFIG_SPACE_1;
	assign CONFIG_SPACE[95:64] = CONFIG_SPACE_2;
	assign CONFIG_SPACE[127:96] = CONFIG_SPACE_3;
	assign CONFIG_SPACE[159:128] = CONFIG_SPACE_4;
	assign CONFIG_SPACE[191:160] = CONFIG_SPACE_5;
	assign CONFIG_SPACE[223:192] = CONFIG_SPACE_6;
	assign CONFIG_SPACE[255:224] = CONFIG_SPACE_7;
	assign CONFIG_SPACE[287:256] = CONFIG_SPACE_8;
	assign CONFIG_SPACE[319:288] = CONFIG_SPACE_9;
	assign CONFIG_SPACE[351:320] = CONFIG_SPACE_10;
	assign CONFIG_SPACE[383:352] = CONFIG_SPACE_11;
	assign CONFIG_SPACE[415:384] = CONFIG_SPACE_12;
	assign CONFIG_SPACE[447:416] = CONFIG_SPACE_13;
	assign CONFIG_SPACE[479:448] = CONFIG_SPACE_14;
	assign CONFIG_SPACE[511:480] = CONFIG_SPACE_15;
	assign CONFIG_SPACE[543:512] = CONFIG_SPACE_16;
	assign CONFIG_SPACE[575:544] = CONFIG_SPACE_17;
	assign CONFIG_SPACE[607:576] = CONFIG_SPACE_18;
	assign CONFIG_SPACE[639:608] = CONFIG_SPACE_19;
	assign CONFIG_SPACE[671:640] = CONFIG_SPACE_20;
	assign CONFIG_SPACE[703:672] = CONFIG_SPACE_21;
	assign CONFIG_SPACE[735:704] = CONFIG_SPACE_22;
	assign CONFIG_SPACE[767:736] = CONFIG_SPACE_23;
	assign CONFIG_SPACE[799:768] = CONFIG_SPACE_24;
	assign CONFIG_SPACE[831:800] = CONFIG_SPACE_25;
	assign CONFIG_SPACE[863:832] = CONFIG_SPACE_26;
	assign CONFIG_SPACE[895:864] = CONFIG_SPACE_27;
	assign CONFIG_SPACE[927:896] = CONFIG_SPACE_28;
	assign CONFIG_SPACE[959:928] = CONFIG_SPACE_29;
	assign CONFIG_SPACE[991:960] = CONFIG_SPACE_30;
	assign CONFIG_SPACE[1023:992] = CONFIG_SPACE_31;
	assign CONFIG_SPACE[1055:1024] = CONFIG_SPACE_32;
	assign CONFIG_SPACE[1087:1056] = CONFIG_SPACE_33;
	assign CONFIG_SPACE[1119:1088] = CONFIG_SPACE_34;
	assign CONFIG_SPACE[1151:1120] = CONFIG_SPACE_35;
	assign CONFIG_SPACE[1183:1152] = CONFIG_SPACE_36;
	assign CONFIG_SPACE[1215:1184] = CONFIG_SPACE_37;
	assign CONFIG_SPACE[1247:1216] = CONFIG_SPACE_38;
	assign CONFIG_SPACE[1279:1248] = CONFIG_SPACE_39;
	assign CONFIG_SPACE[1311:1280] = CONFIG_SPACE_40;
	assign CONFIG_SPACE[1343:1312] = CONFIG_SPACE_41;
	assign CONFIG_SPACE[1375:1344] = CONFIG_SPACE_42;
	assign CONFIG_SPACE[1407:1376] = CONFIG_SPACE_43;
	assign CONFIG_SPACE[1439:1408] = CONFIG_SPACE_44;
	assign CONFIG_SPACE[1458:1440] = CONFIG_SPACE_45;
	fiber_access_16_flat mem_ctrl_fiber_access_16_flat(
		.clk(mem_ctrl_fiber_access_16_flat_clk),
		.clk_en(clk_en),
		.fiber_access_16_inst_buffet_buffet_capacity_log_0(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_buffet_capacity_log_0),
		.fiber_access_16_inst_buffet_buffet_capacity_log_1(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_buffet_capacity_log_1),
		.fiber_access_16_inst_buffet_data_from_mem_lifted_lifted(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_data_from_mem_lifted_lifted),
		.fiber_access_16_inst_buffet_tile_en(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_tile_en),
		.fiber_access_16_inst_read_scanner_block_mode(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_block_mode),
		.fiber_access_16_inst_read_scanner_dense(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_dense),
		.fiber_access_16_inst_read_scanner_dim_size(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_dim_size),
		.fiber_access_16_inst_read_scanner_do_repeat(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_do_repeat),
		.fiber_access_16_inst_read_scanner_inner_dim_offset(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_inner_dim_offset),
		.fiber_access_16_inst_read_scanner_lookup(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_lookup),
		.fiber_access_16_inst_read_scanner_repeat_factor(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_repeat_factor),
		.fiber_access_16_inst_read_scanner_repeat_outer_inner_n(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_repeat_outer_inner_n),
		.fiber_access_16_inst_read_scanner_root(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_root),
		.fiber_access_16_inst_read_scanner_spacc_mode(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_spacc_mode),
		.fiber_access_16_inst_read_scanner_stop_lvl(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_stop_lvl),
		.fiber_access_16_inst_read_scanner_tile_en(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_tile_en),
		.fiber_access_16_inst_tile_en(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_tile_en),
		.fiber_access_16_inst_write_scanner_block_mode(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_block_mode),
		.fiber_access_16_inst_write_scanner_compressed(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_compressed),
		.fiber_access_16_inst_write_scanner_init_blank(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_init_blank),
		.fiber_access_16_inst_write_scanner_lowest_level(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_lowest_level),
		.fiber_access_16_inst_write_scanner_spacc_mode(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_spacc_mode),
		.fiber_access_16_inst_write_scanner_stop_lvl(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_stop_lvl),
		.fiber_access_16_inst_write_scanner_tile_en(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_tile_en),
		.flush(flush),
		.read_scanner_block_rd_out_ready_f_(output_width_17_num_0_fifo_in_ready),
		.read_scanner_coord_out_ready_f_(output_width_17_num_1_fifo_in_ready),
		.read_scanner_pos_out_ready_f_(output_width_17_num_2_fifo_in_ready),
		.read_scanner_us_pos_in_f_(input_width_17_num_0_fifo_out),
		.read_scanner_us_pos_in_valid_f_(input_width_17_num_0_fifo_out_valid),
		.rst_n(rst_n),
		.write_scanner_addr_in_f_(input_width_17_num_1_fifo_out),
		.write_scanner_addr_in_valid_f_(input_width_17_num_1_fifo_out_valid),
		.write_scanner_block_wr_in_f_(input_width_17_num_2_fifo_out),
		.write_scanner_block_wr_in_valid_f_(input_width_17_num_2_fifo_out_valid),
		.write_scanner_data_in_f_(input_width_17_num_3_fifo_out),
		.write_scanner_data_in_valid_f_(input_width_17_num_3_fifo_out_valid),
		.fiber_access_16_inst_buffet_addr_to_mem_lifted_lifted(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_addr_to_mem_lifted_lifted),
		.fiber_access_16_inst_buffet_data_to_mem_lifted_lifted(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_data_to_mem_lifted_lifted),
		.fiber_access_16_inst_buffet_ren_to_mem_lifted_lifted(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_ren_to_mem_lifted_lifted),
		.fiber_access_16_inst_buffet_wen_to_mem_lifted_lifted(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_wen_to_mem_lifted_lifted),
		.read_scanner_block_rd_out_f_(mem_ctrl_fiber_access_16_flat_read_scanner_block_rd_out_f_),
		.read_scanner_block_rd_out_valid_f_(mem_ctrl_fiber_access_16_flat_read_scanner_block_rd_out_valid_f_),
		.read_scanner_coord_out_f_(mem_ctrl_fiber_access_16_flat_read_scanner_coord_out_f_),
		.read_scanner_coord_out_valid_f_(mem_ctrl_fiber_access_16_flat_read_scanner_coord_out_valid_f_),
		.read_scanner_pos_out_f_(mem_ctrl_fiber_access_16_flat_read_scanner_pos_out_f_),
		.read_scanner_pos_out_valid_f_(mem_ctrl_fiber_access_16_flat_read_scanner_pos_out_valid_f_),
		.read_scanner_us_pos_in_ready_f_(mem_ctrl_fiber_access_16_flat_read_scanner_us_pos_in_ready_f_),
		.write_scanner_addr_in_ready_f_(mem_ctrl_fiber_access_16_flat_write_scanner_addr_in_ready_f_),
		.write_scanner_block_wr_in_ready_f_(mem_ctrl_fiber_access_16_flat_write_scanner_block_wr_in_ready_f_),
		.write_scanner_data_in_ready_f_(mem_ctrl_fiber_access_16_flat_write_scanner_data_in_ready_f_)
	);
	strg_ub_vec_flat mem_ctrl_strg_ub_vec_flat(
		.chain_data_in_f_0(MEM_input_width_17_num_0),
		.chain_data_in_f_1(MEM_input_width_17_num_1),
		.clk(mem_ctrl_strg_ub_vec_flat_clk),
		.clk_en(clk_en),
		.data_in_f_0(MEM_input_width_17_num_2),
		.data_in_f_1(MEM_input_width_17_num_3),
		.flush(flush),
		.rst_n(rst_n),
		.strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr),
		.strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0),
		.strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1),
		.strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2),
		.strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr),
		.strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0),
		.strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1),
		.strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2),
		.strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable),
		.strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr),
		.strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0),
		.strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1),
		.strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2),
		.strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable),
		.strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr),
		.strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0),
		.strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1),
		.strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2),
		.strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality),
		.strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0),
		.strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1),
		.strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2),
		.strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality),
		.strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0),
		.strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1),
		.strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2),
		.strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_agg_read_padding(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_agg_read_padding),
		.strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_agg_read_padding(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_agg_read_padding),
		.strg_ub_vec_inst_agg_sram_shared_agg_sram_shared_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_sram_shared_addr_gen_0_starting_addr),
		.strg_ub_vec_inst_agg_sram_shared_agg_sram_shared_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_sram_shared_addr_gen_1_starting_addr),
		.strg_ub_vec_inst_agg_sram_shared_mode_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_mode_0),
		.strg_ub_vec_inst_agg_sram_shared_mode_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_mode_1),
		.strg_ub_vec_inst_chain_chain_en(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en),
		.strg_ub_vec_inst_data_from_strg_lifted(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_data_from_strg_lifted),
		.strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr),
		.strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0),
		.strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1),
		.strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2),
		.strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3),
		.strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4),
		.strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5),
		.strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr),
		.strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0),
		.strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1),
		.strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2),
		.strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3),
		.strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4),
		.strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5),
		.strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality),
		.strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0),
		.strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1),
		.strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2),
		.strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3),
		.strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4),
		.strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5),
		.strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality),
		.strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0),
		.strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1),
		.strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2),
		.strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3),
		.strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4),
		.strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5),
		.strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable),
		.strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_delay(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_delay),
		.strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr),
		.strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0),
		.strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1),
		.strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2),
		.strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3),
		.strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4),
		.strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5),
		.strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable),
		.strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_delay(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_delay),
		.strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr),
		.strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0),
		.strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1),
		.strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2),
		.strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3),
		.strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4),
		.strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5),
		.strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality),
		.strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0),
		.strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1),
		.strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2),
		.strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3),
		.strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4),
		.strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5),
		.strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality),
		.strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0),
		.strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1),
		.strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2),
		.strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3),
		.strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4),
		.strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5),
		.strg_ub_vec_inst_tb_only_shared_tb_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_shared_tb_0),
		.strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr),
		.strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0),
		.strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1),
		.strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2),
		.strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3),
		.strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4),
		.strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5),
		.strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr),
		.strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0),
		.strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1),
		.strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2),
		.strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3),
		.strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4),
		.strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5),
		.strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable),
		.strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_delay(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_delay),
		.strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr),
		.strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0),
		.strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1),
		.strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2),
		.strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3),
		.strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4),
		.strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5),
		.strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable),
		.strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_delay(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_delay),
		.strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr),
		.strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0),
		.strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1),
		.strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2),
		.strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3),
		.strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4),
		.strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5),
		.strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr),
		.strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0),
		.strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1),
		.strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2),
		.strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3),
		.strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4),
		.strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5),
		.strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr),
		.strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0),
		.strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1),
		.strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2),
		.strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3),
		.strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4),
		.strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5),
		.accessor_output_f_b_0(mem_ctrl_strg_ub_vec_flat_accessor_output_f_b_0),
		.accessor_output_f_b_1(mem_ctrl_strg_ub_vec_flat_accessor_output_f_b_1),
		.data_out_f_0(mem_ctrl_strg_ub_vec_flat_data_out_f_0),
		.data_out_f_1(mem_ctrl_strg_ub_vec_flat_data_out_f_1),
		.strg_ub_vec_inst_addr_out_lifted(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_addr_out_lifted),
		.strg_ub_vec_inst_data_to_strg_lifted(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_data_to_strg_lifted),
		.strg_ub_vec_inst_ren_to_strg_lifted(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_ren_to_strg_lifted),
		.strg_ub_vec_inst_wen_to_strg_lifted(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_wen_to_strg_lifted)
	);
	strg_ram_64_512_delay1_flat mem_ctrl_strg_ram_64_512_delay1_flat(
		.clk(mem_ctrl_strg_ram_64_512_delay1_flat_clk),
		.clk_en(clk_en),
		.data_in_f_(MEM_input_width_17_num_0),
		.flush(flush),
		.rd_addr_in_f_(MEM_input_width_17_num_1),
		.ren_f_(MEM_input_width_1_num_0),
		.rst_n(rst_n),
		.strg_ram_64_512_delay1_inst_data_from_strg_lifted(mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_data_from_strg_lifted),
		.wen_f_(MEM_input_width_1_num_1),
		.wr_addr_in_f_(MEM_input_width_17_num_2),
		.data_out_f_(mem_ctrl_strg_ram_64_512_delay1_flat_data_out_f_),
		.ready_f_(mem_ctrl_strg_ram_64_512_delay1_flat_ready_f_),
		.strg_ram_64_512_delay1_inst_addr_out_lifted(mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_addr_out_lifted),
		.strg_ram_64_512_delay1_inst_data_to_strg_lifted(mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_data_to_strg_lifted),
		.strg_ram_64_512_delay1_inst_ren_to_strg_lifted(mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_ren_to_strg_lifted),
		.strg_ram_64_512_delay1_inst_wen_to_strg_lifted(mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_wen_to_strg_lifted),
		.valid_out_f_(mem_ctrl_strg_ram_64_512_delay1_flat_valid_out_f_)
	);
	stencil_valid_flat mem_ctrl_stencil_valid_flat(
		.clk(mem_ctrl_stencil_valid_flat_clk),
		.clk_en(clk_en),
		.flush(flush),
		.rst_n(rst_n),
		.stencil_valid_inst_loops_stencil_valid_dimensionality(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality),
		.stencil_valid_inst_loops_stencil_valid_ranges_0(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_0),
		.stencil_valid_inst_loops_stencil_valid_ranges_1(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_1),
		.stencil_valid_inst_loops_stencil_valid_ranges_2(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_2),
		.stencil_valid_inst_loops_stencil_valid_ranges_3(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_3),
		.stencil_valid_inst_loops_stencil_valid_ranges_4(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_4),
		.stencil_valid_inst_loops_stencil_valid_ranges_5(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_5),
		.stencil_valid_inst_stencil_valid_sched_gen_enable(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable),
		.stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr),
		.stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0),
		.stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1),
		.stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2),
		.stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3),
		.stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4),
		.stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5),
		.stencil_valid_f_(mem_ctrl_stencil_valid_flat_stencil_valid_f_)
	);
	reg_fifo_depth_2_w_17_afd_2 input_width_17_num_0_input_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(MEM_input_width_17_num_0),
		.flush(flush),
		.pop(input_width_17_num_0_fifo_out_ready),
		.push(MEM_input_width_17_num_0_valid),
		.rst_n(rst_n),
		.data_out(input_width_17_num_0_fifo_out),
		.empty(input_width_17_num_0_input_fifo_empty),
		.full(input_width_17_num_0_input_fifo_full)
	);
	reg_fifo_depth_2_w_17_afd_2 input_width_17_num_1_input_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(MEM_input_width_17_num_1),
		.flush(flush),
		.pop(input_width_17_num_1_fifo_out_ready),
		.push(MEM_input_width_17_num_1_valid),
		.rst_n(rst_n),
		.data_out(input_width_17_num_1_fifo_out),
		.empty(input_width_17_num_1_input_fifo_empty),
		.full(input_width_17_num_1_input_fifo_full)
	);
	reg_fifo_depth_2_w_17_afd_2 input_width_17_num_2_input_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(MEM_input_width_17_num_2),
		.flush(flush),
		.pop(input_width_17_num_2_fifo_out_ready),
		.push(MEM_input_width_17_num_2_valid),
		.rst_n(rst_n),
		.data_out(input_width_17_num_2_fifo_out),
		.empty(input_width_17_num_2_input_fifo_empty),
		.full(input_width_17_num_2_input_fifo_full)
	);
	reg_fifo_depth_2_w_17_afd_2 input_width_17_num_3_input_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(MEM_input_width_17_num_3),
		.flush(flush),
		.pop(input_width_17_num_3_fifo_out_ready),
		.push(MEM_input_width_17_num_3_valid),
		.rst_n(rst_n),
		.data_out(input_width_17_num_3_fifo_out),
		.empty(input_width_17_num_3_input_fifo_empty),
		.full(input_width_17_num_3_input_fifo_full)
	);
	reg_fifo_depth_2_w_17_afd_2 output_width_17_num_0_output_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(output_width_17_num_0_fifo_in),
		.flush(flush),
		.pop(MEM_output_width_17_num_0_ready),
		.push(output_width_17_num_0_fifo_in_valid),
		.rst_n(rst_n),
		.data_out(output_width_17_num_0_output_fifo_data_out),
		.empty(output_width_17_num_0_output_fifo_empty),
		.full(output_width_17_num_0_output_fifo_full)
	);
	reg_fifo_depth_2_w_17_afd_2 output_width_17_num_1_output_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(output_width_17_num_1_fifo_in),
		.flush(flush),
		.pop(MEM_output_width_17_num_1_ready),
		.push(output_width_17_num_1_fifo_in_valid),
		.rst_n(rst_n),
		.data_out(output_width_17_num_1_output_fifo_data_out),
		.empty(output_width_17_num_1_output_fifo_empty),
		.full(output_width_17_num_1_output_fifo_full)
	);
	reg_fifo_depth_2_w_17_afd_2 output_width_17_num_2_output_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(output_width_17_num_2_fifo_in),
		.flush(flush),
		.pop(MEM_output_width_17_num_2_ready),
		.push(output_width_17_num_2_fifo_in_valid),
		.rst_n(rst_n),
		.data_out(output_width_17_num_2_output_fifo_data_out),
		.empty(output_width_17_num_2_output_fifo_empty),
		.full(output_width_17_num_2_output_fifo_full)
	);
	sram_sp__0 memory_0(
		.clk(gclk),
		.clk_en(memory_0_clk_en),
		.data_in_p0(memory_0_data_in_p0),
		.flush(flush),
		.read_addr_p0(memory_0_read_addr_p0),
		.read_enable_p0(memory_0_read_enable_p0),
		.write_addr_p0(memory_0_write_addr_p0),
		.write_enable_p0(memory_0_write_enable_p0),
		.data_out_p0(memory_0_data_out_p0)
	);
	storage_config_seq_2_64_16 config_seq(
		.clk(gclk),
		.clk_en(config_seq_clk_en),
		.config_addr_in(config_addr_in),
		.config_data_in(config_data_in_shrt),
		.config_en(config_en),
		.config_rd(config_read),
		.config_wr(config_write),
		.flush(flush),
		.rd_data_stg(config_seq_rd_data_stg),
		.rst_n(rst_n),
		.addr_out(config_seq_addr_out),
		.rd_data_out(config_data_out_shrt),
		.ren_out(config_seq_ren_out),
		.wen_out(config_seq_wen_out),
		.wr_data(config_seq_wr_data)
	);
endmodule
module MemCore_inner_W (
	CONFIG_SPACE_0,
	CONFIG_SPACE_1,
	CONFIG_SPACE_10,
	CONFIG_SPACE_11,
	CONFIG_SPACE_12,
	CONFIG_SPACE_13,
	CONFIG_SPACE_14,
	CONFIG_SPACE_15,
	CONFIG_SPACE_16,
	CONFIG_SPACE_17,
	CONFIG_SPACE_18,
	CONFIG_SPACE_19,
	CONFIG_SPACE_2,
	CONFIG_SPACE_20,
	CONFIG_SPACE_21,
	CONFIG_SPACE_22,
	CONFIG_SPACE_23,
	CONFIG_SPACE_24,
	CONFIG_SPACE_25,
	CONFIG_SPACE_26,
	CONFIG_SPACE_27,
	CONFIG_SPACE_28,
	CONFIG_SPACE_29,
	CONFIG_SPACE_3,
	CONFIG_SPACE_30,
	CONFIG_SPACE_31,
	CONFIG_SPACE_32,
	CONFIG_SPACE_33,
	CONFIG_SPACE_34,
	CONFIG_SPACE_35,
	CONFIG_SPACE_36,
	CONFIG_SPACE_37,
	CONFIG_SPACE_38,
	CONFIG_SPACE_39,
	CONFIG_SPACE_4,
	CONFIG_SPACE_40,
	CONFIG_SPACE_41,
	CONFIG_SPACE_42,
	CONFIG_SPACE_43,
	CONFIG_SPACE_44,
	CONFIG_SPACE_45,
	CONFIG_SPACE_5,
	CONFIG_SPACE_6,
	CONFIG_SPACE_7,
	CONFIG_SPACE_8,
	CONFIG_SPACE_9,
	MEM_input_width_17_num_0,
	MEM_input_width_17_num_0_valid,
	MEM_input_width_17_num_1,
	MEM_input_width_17_num_1_valid,
	MEM_input_width_17_num_2,
	MEM_input_width_17_num_2_valid,
	MEM_input_width_17_num_3,
	MEM_input_width_17_num_3_valid,
	MEM_input_width_1_num_0,
	MEM_input_width_1_num_1,
	MEM_output_width_17_num_0_ready,
	MEM_output_width_17_num_1_ready,
	MEM_output_width_17_num_2_ready,
	clk,
	clk_en,
	config_addr_in,
	config_data_in,
	config_en,
	config_read,
	config_write,
	flush,
	mode,
	mode_excl,
	rst_n,
	tile_en,
	MEM_input_width_17_num_0_ready,
	MEM_input_width_17_num_1_ready,
	MEM_input_width_17_num_2_ready,
	MEM_input_width_17_num_3_ready,
	MEM_output_width_17_num_0,
	MEM_output_width_17_num_0_valid,
	MEM_output_width_17_num_1,
	MEM_output_width_17_num_1_valid,
	MEM_output_width_17_num_2,
	MEM_output_width_17_num_2_valid,
	MEM_output_width_1_num_0,
	MEM_output_width_1_num_1,
	MEM_output_width_1_num_2,
	config_data_out_0,
	config_data_out_1
);
	input wire [31:0] CONFIG_SPACE_0;
	input wire [31:0] CONFIG_SPACE_1;
	input wire [31:0] CONFIG_SPACE_10;
	input wire [31:0] CONFIG_SPACE_11;
	input wire [31:0] CONFIG_SPACE_12;
	input wire [31:0] CONFIG_SPACE_13;
	input wire [31:0] CONFIG_SPACE_14;
	input wire [31:0] CONFIG_SPACE_15;
	input wire [31:0] CONFIG_SPACE_16;
	input wire [31:0] CONFIG_SPACE_17;
	input wire [31:0] CONFIG_SPACE_18;
	input wire [31:0] CONFIG_SPACE_19;
	input wire [31:0] CONFIG_SPACE_2;
	input wire [31:0] CONFIG_SPACE_20;
	input wire [31:0] CONFIG_SPACE_21;
	input wire [31:0] CONFIG_SPACE_22;
	input wire [31:0] CONFIG_SPACE_23;
	input wire [31:0] CONFIG_SPACE_24;
	input wire [31:0] CONFIG_SPACE_25;
	input wire [31:0] CONFIG_SPACE_26;
	input wire [31:0] CONFIG_SPACE_27;
	input wire [31:0] CONFIG_SPACE_28;
	input wire [31:0] CONFIG_SPACE_29;
	input wire [31:0] CONFIG_SPACE_3;
	input wire [31:0] CONFIG_SPACE_30;
	input wire [31:0] CONFIG_SPACE_31;
	input wire [31:0] CONFIG_SPACE_32;
	input wire [31:0] CONFIG_SPACE_33;
	input wire [31:0] CONFIG_SPACE_34;
	input wire [31:0] CONFIG_SPACE_35;
	input wire [31:0] CONFIG_SPACE_36;
	input wire [31:0] CONFIG_SPACE_37;
	input wire [31:0] CONFIG_SPACE_38;
	input wire [31:0] CONFIG_SPACE_39;
	input wire [31:0] CONFIG_SPACE_4;
	input wire [31:0] CONFIG_SPACE_40;
	input wire [31:0] CONFIG_SPACE_41;
	input wire [31:0] CONFIG_SPACE_42;
	input wire [31:0] CONFIG_SPACE_43;
	input wire [31:0] CONFIG_SPACE_44;
	input wire [18:0] CONFIG_SPACE_45;
	input wire [31:0] CONFIG_SPACE_5;
	input wire [31:0] CONFIG_SPACE_6;
	input wire [31:0] CONFIG_SPACE_7;
	input wire [31:0] CONFIG_SPACE_8;
	input wire [31:0] CONFIG_SPACE_9;
	input wire [16:0] MEM_input_width_17_num_0;
	input wire MEM_input_width_17_num_0_valid;
	input wire [16:0] MEM_input_width_17_num_1;
	input wire MEM_input_width_17_num_1_valid;
	input wire [16:0] MEM_input_width_17_num_2;
	input wire MEM_input_width_17_num_2_valid;
	input wire [16:0] MEM_input_width_17_num_3;
	input wire MEM_input_width_17_num_3_valid;
	input wire MEM_input_width_1_num_0;
	input wire MEM_input_width_1_num_1;
	input wire MEM_output_width_17_num_0_ready;
	input wire MEM_output_width_17_num_1_ready;
	input wire MEM_output_width_17_num_2_ready;
	input wire clk;
	input wire clk_en;
	input wire [7:0] config_addr_in;
	input wire [31:0] config_data_in;
	input wire [1:0] config_en;
	input wire config_read;
	input wire config_write;
	input wire flush;
	input wire [1:0] mode;
	input wire mode_excl;
	input wire rst_n;
	input wire tile_en;
	output wire MEM_input_width_17_num_0_ready;
	output wire MEM_input_width_17_num_1_ready;
	output wire MEM_input_width_17_num_2_ready;
	output wire MEM_input_width_17_num_3_ready;
	output wire [16:0] MEM_output_width_17_num_0;
	output wire MEM_output_width_17_num_0_valid;
	output wire [16:0] MEM_output_width_17_num_1;
	output wire MEM_output_width_17_num_1_valid;
	output wire [16:0] MEM_output_width_17_num_2;
	output wire MEM_output_width_17_num_2_valid;
	output wire MEM_output_width_1_num_0;
	output wire MEM_output_width_1_num_1;
	output wire MEM_output_width_1_num_2;
	output wire [31:0] config_data_out_0;
	output wire [31:0] config_data_out_1;
	wire [63:0] MemCore_inner_config_data_out;
	assign config_data_out_0 = MemCore_inner_config_data_out[0+:32];
	assign config_data_out_1 = MemCore_inner_config_data_out[32+:32];
	MemCore_inner MemCore_inner(
		.CONFIG_SPACE_0(CONFIG_SPACE_0),
		.CONFIG_SPACE_1(CONFIG_SPACE_1),
		.CONFIG_SPACE_10(CONFIG_SPACE_10),
		.CONFIG_SPACE_11(CONFIG_SPACE_11),
		.CONFIG_SPACE_12(CONFIG_SPACE_12),
		.CONFIG_SPACE_13(CONFIG_SPACE_13),
		.CONFIG_SPACE_14(CONFIG_SPACE_14),
		.CONFIG_SPACE_15(CONFIG_SPACE_15),
		.CONFIG_SPACE_16(CONFIG_SPACE_16),
		.CONFIG_SPACE_17(CONFIG_SPACE_17),
		.CONFIG_SPACE_18(CONFIG_SPACE_18),
		.CONFIG_SPACE_19(CONFIG_SPACE_19),
		.CONFIG_SPACE_2(CONFIG_SPACE_2),
		.CONFIG_SPACE_20(CONFIG_SPACE_20),
		.CONFIG_SPACE_21(CONFIG_SPACE_21),
		.CONFIG_SPACE_22(CONFIG_SPACE_22),
		.CONFIG_SPACE_23(CONFIG_SPACE_23),
		.CONFIG_SPACE_24(CONFIG_SPACE_24),
		.CONFIG_SPACE_25(CONFIG_SPACE_25),
		.CONFIG_SPACE_26(CONFIG_SPACE_26),
		.CONFIG_SPACE_27(CONFIG_SPACE_27),
		.CONFIG_SPACE_28(CONFIG_SPACE_28),
		.CONFIG_SPACE_29(CONFIG_SPACE_29),
		.CONFIG_SPACE_3(CONFIG_SPACE_3),
		.CONFIG_SPACE_30(CONFIG_SPACE_30),
		.CONFIG_SPACE_31(CONFIG_SPACE_31),
		.CONFIG_SPACE_32(CONFIG_SPACE_32),
		.CONFIG_SPACE_33(CONFIG_SPACE_33),
		.CONFIG_SPACE_34(CONFIG_SPACE_34),
		.CONFIG_SPACE_35(CONFIG_SPACE_35),
		.CONFIG_SPACE_36(CONFIG_SPACE_36),
		.CONFIG_SPACE_37(CONFIG_SPACE_37),
		.CONFIG_SPACE_38(CONFIG_SPACE_38),
		.CONFIG_SPACE_39(CONFIG_SPACE_39),
		.CONFIG_SPACE_4(CONFIG_SPACE_4),
		.CONFIG_SPACE_40(CONFIG_SPACE_40),
		.CONFIG_SPACE_41(CONFIG_SPACE_41),
		.CONFIG_SPACE_42(CONFIG_SPACE_42),
		.CONFIG_SPACE_43(CONFIG_SPACE_43),
		.CONFIG_SPACE_44(CONFIG_SPACE_44),
		.CONFIG_SPACE_45(CONFIG_SPACE_45),
		.CONFIG_SPACE_5(CONFIG_SPACE_5),
		.CONFIG_SPACE_6(CONFIG_SPACE_6),
		.CONFIG_SPACE_7(CONFIG_SPACE_7),
		.CONFIG_SPACE_8(CONFIG_SPACE_8),
		.CONFIG_SPACE_9(CONFIG_SPACE_9),
		.MEM_input_width_17_num_0(MEM_input_width_17_num_0),
		.MEM_input_width_17_num_0_valid(MEM_input_width_17_num_0_valid),
		.MEM_input_width_17_num_1(MEM_input_width_17_num_1),
		.MEM_input_width_17_num_1_valid(MEM_input_width_17_num_1_valid),
		.MEM_input_width_17_num_2(MEM_input_width_17_num_2),
		.MEM_input_width_17_num_2_valid(MEM_input_width_17_num_2_valid),
		.MEM_input_width_17_num_3(MEM_input_width_17_num_3),
		.MEM_input_width_17_num_3_valid(MEM_input_width_17_num_3_valid),
		.MEM_input_width_1_num_0(MEM_input_width_1_num_0),
		.MEM_input_width_1_num_1(MEM_input_width_1_num_1),
		.MEM_output_width_17_num_0_ready(MEM_output_width_17_num_0_ready),
		.MEM_output_width_17_num_1_ready(MEM_output_width_17_num_1_ready),
		.MEM_output_width_17_num_2_ready(MEM_output_width_17_num_2_ready),
		.clk(clk),
		.clk_en(clk_en),
		.config_addr_in(config_addr_in),
		.config_data_in(config_data_in),
		.config_en(config_en),
		.config_read(config_read),
		.config_write(config_write),
		.flush(flush),
		.mode(mode),
		.mode_excl(mode_excl),
		.rst_n(rst_n),
		.tile_en(tile_en),
		.MEM_input_width_17_num_0_ready(MEM_input_width_17_num_0_ready),
		.MEM_input_width_17_num_1_ready(MEM_input_width_17_num_1_ready),
		.MEM_input_width_17_num_2_ready(MEM_input_width_17_num_2_ready),
		.MEM_input_width_17_num_3_ready(MEM_input_width_17_num_3_ready),
		.MEM_output_width_17_num_0(MEM_output_width_17_num_0),
		.MEM_output_width_17_num_0_valid(MEM_output_width_17_num_0_valid),
		.MEM_output_width_17_num_1(MEM_output_width_17_num_1),
		.MEM_output_width_17_num_1_valid(MEM_output_width_17_num_1_valid),
		.MEM_output_width_17_num_2(MEM_output_width_17_num_2),
		.MEM_output_width_17_num_2_valid(MEM_output_width_17_num_2_valid),
		.MEM_output_width_1_num_0(MEM_output_width_1_num_0),
		.MEM_output_width_1_num_1(MEM_output_width_1_num_1),
		.MEM_output_width_1_num_2(MEM_output_width_1_num_2),
		.config_data_out(MemCore_inner_config_data_out)
	);
endmodule
module addr_gen_3_16 (
	clk,
	clk_en,
	flush,
	mux_sel,
	restart,
	rst_n,
	starting_addr,
	step,
	strides,
	addr_out
);
	input wire clk;
	input wire clk_en;
	input wire flush;
	input wire [1:0] mux_sel;
	input wire restart;
	input wire rst_n;
	input wire [15:0] starting_addr;
	input wire step;
	input wire [47:0] strides;
	output wire [15:0] addr_out;
	wire [15:0] calc_addr;
	reg [15:0] current_addr;
	wire [15:0] strt_addr;
	assign strt_addr = starting_addr;
	assign addr_out = calc_addr;
	assign calc_addr = current_addr;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			current_addr <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				current_addr <= strt_addr;
			else if (step) begin
				if (restart)
					current_addr <= strt_addr;
				else
					current_addr <= current_addr + strides[mux_sel * 16+:16];
			end
		end
endmodule
module addr_gen_3_3 (
	clk,
	clk_en,
	flush,
	mux_sel,
	restart,
	rst_n,
	starting_addr,
	step,
	strides,
	addr_out
);
	input wire clk;
	input wire clk_en;
	input wire flush;
	input wire [1:0] mux_sel;
	input wire restart;
	input wire rst_n;
	input wire [2:0] starting_addr;
	input wire step;
	input wire [8:0] strides;
	output wire [2:0] addr_out;
	wire [2:0] calc_addr;
	reg [2:0] current_addr;
	wire [2:0] strt_addr;
	assign strt_addr = starting_addr;
	assign addr_out = calc_addr;
	assign calc_addr = current_addr;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			current_addr <= 3'h0;
		else if (clk_en) begin
			if (flush)
				current_addr <= strt_addr;
			else if (step) begin
				if (restart)
					current_addr <= strt_addr;
				else
					current_addr <= current_addr + strides[mux_sel * 3+:3];
			end
		end
endmodule
module addr_gen_6_16 (
	clk,
	clk_en,
	flush,
	mux_sel,
	restart,
	rst_n,
	starting_addr,
	step,
	strides,
	addr_out
);
	input wire clk;
	input wire clk_en;
	input wire flush;
	input wire [2:0] mux_sel;
	input wire restart;
	input wire rst_n;
	input wire [15:0] starting_addr;
	input wire step;
	input wire [95:0] strides;
	output wire [15:0] addr_out;
	wire [15:0] calc_addr;
	reg [15:0] current_addr;
	wire [15:0] strt_addr;
	assign strt_addr = starting_addr;
	assign addr_out = calc_addr;
	assign calc_addr = current_addr;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			current_addr <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				current_addr <= strt_addr;
			else if (step) begin
				if (restart)
					current_addr <= strt_addr;
				else
					current_addr <= current_addr + strides[mux_sel * 16+:16];
			end
		end
endmodule
module addr_gen_6_16_delay_addr_10 (
	clk,
	clk_en,
	delay,
	flush,
	mux_sel,
	restart,
	rst_n,
	starting_addr,
	step,
	strides,
	addr_out,
	delay_out,
	delayed_addr_out
);
	input wire clk;
	input wire clk_en;
	input wire [9:0] delay;
	input wire flush;
	input wire [2:0] mux_sel;
	input wire restart;
	input wire rst_n;
	input wire [15:0] starting_addr;
	input wire step;
	input wire [95:0] strides;
	output wire [15:0] addr_out;
	output wire [9:0] delay_out;
	output wire [15:0] delayed_addr_out;
	wire [15:0] calc_addr;
	reg [15:0] current_addr;
	wire [15:0] strt_addr;
	assign delay_out = delay;
	assign strt_addr = starting_addr;
	assign addr_out = calc_addr;
	assign calc_addr = current_addr;
	function automatic [15:0] sv2v_cast_16;
		input reg [15:0] inp;
		sv2v_cast_16 = inp;
	endfunction
	assign delayed_addr_out = current_addr + sv2v_cast_16(delay);
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			current_addr <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				current_addr <= strt_addr;
			else if (step) begin
				if (restart)
					current_addr <= strt_addr;
				else
					current_addr <= current_addr + strides[mux_sel * 16+:16];
			end
		end
endmodule
module addr_gen_6_4 (
	clk,
	clk_en,
	flush,
	mux_sel,
	restart,
	rst_n,
	starting_addr,
	step,
	strides,
	addr_out
);
	input wire clk;
	input wire clk_en;
	input wire flush;
	input wire [2:0] mux_sel;
	input wire restart;
	input wire rst_n;
	input wire [3:0] starting_addr;
	input wire step;
	input wire [23:0] strides;
	output wire [3:0] addr_out;
	wire [3:0] calc_addr;
	reg [3:0] current_addr;
	wire [3:0] strt_addr;
	assign strt_addr = starting_addr;
	assign addr_out = calc_addr;
	assign calc_addr = current_addr;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			current_addr <= 4'h0;
		else if (clk_en) begin
			if (flush)
				current_addr <= strt_addr;
			else if (step) begin
				if (restart)
					current_addr <= strt_addr;
				else
					current_addr <= current_addr + strides[mux_sel * 4+:4];
			end
		end
endmodule
module addr_gen_6_9 (
	clk,
	clk_en,
	flush,
	mux_sel,
	restart,
	rst_n,
	starting_addr,
	step,
	strides,
	addr_out
);
	input wire clk;
	input wire clk_en;
	input wire flush;
	input wire [2:0] mux_sel;
	input wire restart;
	input wire rst_n;
	input wire [8:0] starting_addr;
	input wire step;
	input wire [53:0] strides;
	output wire [8:0] addr_out;
	wire [8:0] calc_addr;
	reg [8:0] current_addr;
	wire [8:0] strt_addr;
	assign strt_addr = starting_addr;
	assign addr_out = calc_addr;
	assign calc_addr = current_addr;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			current_addr <= 9'h000;
		else if (clk_en) begin
			if (flush)
				current_addr <= strt_addr;
			else if (step) begin
				if (restart)
					current_addr <= strt_addr;
				else
					current_addr <= current_addr + strides[mux_sel * 9+:9];
			end
		end
endmodule
module agg_sram_shared_addr_gen (
	clk,
	clk_en,
	flush,
	mode,
	rst_n,
	sram_read,
	sram_read_addr,
	starting_addr,
	step,
	addr_out
);
	input wire clk;
	input wire clk_en;
	input wire flush;
	input wire [1:0] mode;
	input wire rst_n;
	input wire [1:0] sram_read;
	input wire [17:0] sram_read_addr;
	input wire [8:0] starting_addr;
	input wire step;
	output wire [8:0] addr_out;
	reg [35:0] addr_fifo;
	wire [8:0] addr_fifo_in;
	reg [8:0] addr_fifo_out;
	wire addr_fifo_wr_en;
	reg [8:0] lin_addr_cnter;
	reg [1:0] rd_ptr;
	reg [1:0] wr_ptr;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			lin_addr_cnter <= 9'h000;
		else if (clk_en) begin
			if (flush)
				lin_addr_cnter <= 9'h000;
			else if (mode[1] == 1'h0) begin
				if (step) begin
					if (lin_addr_cnter == 9'h1ff)
						lin_addr_cnter <= 9'h000;
					else
						lin_addr_cnter <= lin_addr_cnter + 9'h001;
				end
			end
		end
	assign addr_fifo_wr_en = (mode[0] ? sram_read[1] : sram_read[0]);
	assign addr_fifo_in = (mode[0] ? sram_read_addr[9+:9] : sram_read_addr[0+:9]);
	always @(posedge clk or negedge rst_n)
		if (~rst_n) begin
			wr_ptr <= 2'h0;
			rd_ptr <= 2'h0;
			addr_fifo <= 36'h000000000;
			addr_fifo_out <= 9'h000;
		end
		else if (clk_en) begin
			if (flush) begin
				wr_ptr <= 2'h0;
				rd_ptr <= 2'h0;
				addr_fifo <= 36'h000000000;
				addr_fifo_out <= 9'h000;
			end
			else if (mode[1] == 1'h1) begin
				if (addr_fifo_wr_en) begin
					wr_ptr <= wr_ptr + 2'h1;
					addr_fifo[wr_ptr * 9+:9] <= addr_fifo_in;
				end
				if (step)
					rd_ptr <= rd_ptr + 2'h1;
				addr_fifo_out <= addr_fifo[rd_ptr * 9+:9];
			end
		end
	assign addr_out = (mode[1] ? addr_fifo_out : lin_addr_cnter + starting_addr);
endmodule
module agg_sram_shared_sched_gen (
	agg_read_padding,
	agg_write,
	agg_write_addr_l2b,
	agg_write_mux_sel,
	agg_write_restart,
	clk,
	clk_en,
	flush,
	mode,
	rst_n,
	sram_read_d,
	valid_output
);
	input wire [7:0] agg_read_padding;
	input wire agg_write;
	input wire [1:0] agg_write_addr_l2b;
	input wire [2:0] agg_write_mux_sel;
	input wire agg_write_restart;
	input wire clk;
	input wire clk_en;
	input wire flush;
	input wire [1:0] mode;
	input wire rst_n;
	input wire [1:0] sram_read_d;
	output reg valid_output;
	reg agg_write_4_r;
	reg [7:0] pad_cnt;
	reg pad_cnt_en;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			agg_write_4_r <= 1'h0;
		else if (clk_en) begin
			if (flush)
				agg_write_4_r <= 1'h0;
			else if (mode[1] == 1'h0)
				agg_write_4_r <= agg_write & &agg_write_addr_l2b;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n) begin
			pad_cnt_en <= 1'h0;
			pad_cnt <= 8'h00;
		end
		else if (clk_en) begin
			if (flush) begin
				pad_cnt_en <= 1'h0;
				pad_cnt <= 8'h00;
			end
			else if ((mode[1] == 1'h0) & (agg_read_padding != 8'h00)) begin
				if (agg_write & ((agg_write_mux_sel != 3'h0) | agg_write_restart))
					pad_cnt_en <= 1'h1;
				else if (pad_cnt == agg_read_padding)
					pad_cnt_en <= 1'h0;
				if (pad_cnt == agg_read_padding)
					pad_cnt <= 8'h00;
				else if (pad_cnt_en | (agg_write & ((agg_write_mux_sel != 3'h0) | agg_write_restart)))
					pad_cnt <= pad_cnt + 8'h01;
			end
		end
	always @(*)
		if (mode[1] == 1'h0) begin
			if (agg_read_padding != 8'h00)
				valid_output = (agg_read_padding == pad_cnt) | agg_write_4_r;
			else
				valid_output = agg_write_4_r;
		end
		else
			valid_output = (mode[0] ? sram_read_d[1] : sram_read_d[0]);
endmodule
module arbiter_2_in_PRIO_algo (
	clk,
	clk_en,
	flush,
	request_in,
	resource_ready,
	rst_n,
	grant_out
);
	input wire clk;
	input wire clk_en;
	input wire flush;
	input wire [1:0] request_in;
	input wire resource_ready;
	input wire rst_n;
	output wire [1:0] grant_out;
	reg [1:0] grant_line;
	wire [1:0] grant_line_ready;
	wire [1:0] grant_out_consolation;
	wire [1:0] grant_out_priority;
	reg tmp_done;
	reg tmp_out_first;
	always @(*) grant_line = (request_in[1] ? 2'h2 : 2'h1);
	assign grant_line_ready[0] = grant_line[0] & resource_ready;
	assign grant_out_priority[0] = grant_line_ready[0] & request_in[0];
	assign grant_line_ready[1] = grant_line[1] & resource_ready;
	assign grant_out_priority[1] = grant_line_ready[1] & request_in[1];
	always @(*) begin
		tmp_done = 1'h0;
		tmp_out_first = 1'h0;
		if (~tmp_done) begin
			if (request_in[0]) begin
				tmp_out_first = 1'h0;
				tmp_done = 1'h1;
			end
		end
		if (~tmp_done) begin
			if (request_in[1]) begin
				tmp_out_first = 1'h1;
				tmp_done = 1'h1;
			end
		end
	end
	assign grant_out_consolation[0] = (resource_ready & request_in[0]) & (tmp_out_first == 1'h0);
	assign grant_out[0] = (|grant_out_priority ? grant_out_priority[0] : grant_out_consolation[0]);
	assign grant_out_consolation[1] = (resource_ready & request_in[1]) & (tmp_out_first == 1'h1);
	assign grant_out[1] = (|grant_out_priority ? grant_out_priority[1] : grant_out_consolation[1]);
endmodule
module arbiter_4_in_RR_algo (
	clk,
	clk_en,
	flush,
	request_in,
	resource_ready,
	rst_n,
	grant_out
);
	input wire clk;
	input wire clk_en;
	input wire flush;
	input wire [3:0] request_in;
	input wire resource_ready;
	input wire rst_n;
	output wire [3:0] grant_out;
	reg [3:0] grant_line;
	wire [3:0] grant_line_ready;
	wire [3:0] grant_out_consolation;
	wire [3:0] grant_out_priority;
	reg tmp_done;
	reg [1:0] tmp_out_first;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			grant_line <= 4'h1;
		else if (clk_en) begin
			if (flush)
				grant_line <= 4'h1;
			else
				grant_line <= {grant_line[2:0], grant_line[3]};
		end
	assign grant_line_ready[0] = grant_line[0] & resource_ready;
	assign grant_out_priority[0] = grant_line_ready[0] & request_in[0];
	assign grant_line_ready[1] = grant_line[1] & resource_ready;
	assign grant_out_priority[1] = grant_line_ready[1] & request_in[1];
	assign grant_line_ready[2] = grant_line[2] & resource_ready;
	assign grant_out_priority[2] = grant_line_ready[2] & request_in[2];
	assign grant_line_ready[3] = grant_line[3] & resource_ready;
	assign grant_out_priority[3] = grant_line_ready[3] & request_in[3];
	always @(*) begin
		tmp_done = 1'h0;
		tmp_out_first = 2'h0;
		if (~tmp_done) begin
			if (request_in[0]) begin
				tmp_out_first = 2'h0;
				tmp_done = 1'h1;
			end
		end
		if (~tmp_done) begin
			if (request_in[1]) begin
				tmp_out_first = 2'h1;
				tmp_done = 1'h1;
			end
		end
		if (~tmp_done) begin
			if (request_in[2]) begin
				tmp_out_first = 2'h2;
				tmp_done = 1'h1;
			end
		end
		if (~tmp_done) begin
			if (request_in[3]) begin
				tmp_out_first = 2'h3;
				tmp_done = 1'h1;
			end
		end
	end
	assign grant_out_consolation[0] = (resource_ready & request_in[0]) & (tmp_out_first == 2'h0);
	assign grant_out[0] = (|grant_out_priority ? grant_out_priority[0] : grant_out_consolation[0]);
	assign grant_out_consolation[1] = (resource_ready & request_in[1]) & (tmp_out_first == 2'h1);
	assign grant_out[1] = (|grant_out_priority ? grant_out_priority[1] : grant_out_consolation[1]);
	assign grant_out_consolation[2] = (resource_ready & request_in[2]) & (tmp_out_first == 2'h2);
	assign grant_out[2] = (|grant_out_priority ? grant_out_priority[2] : grant_out_consolation[2]);
	assign grant_out_consolation[3] = (resource_ready & request_in[3]) & (tmp_out_first == 2'h3);
	assign grant_out[3] = (|grant_out_priority ? grant_out_priority[3] : grant_out_consolation[3]);
endmodule
module buffet_like_16 (
	buffet_capacity_log,
	clk,
	clk_en,
	data_from_mem,
	flush,
	rd_ID,
	rd_ID_valid,
	rd_addr,
	rd_addr_valid,
	rd_op,
	rd_op_valid,
	rd_rsp_data_ready,
	rst_n,
	tile_en,
	wr_ID,
	wr_ID_valid,
	wr_addr,
	wr_addr_valid,
	wr_data,
	wr_data_valid,
	addr_to_mem,
	data_to_mem,
	rd_ID_ready,
	rd_addr_ready,
	rd_op_ready,
	rd_rsp_data,
	rd_rsp_data_valid,
	ren_to_mem,
	wen_to_mem,
	wr_ID_ready,
	wr_addr_ready,
	wr_data_ready
);
	input wire [7:0] buffet_capacity_log;
	input wire clk;
	input wire clk_en;
	input wire [63:0] data_from_mem;
	input wire flush;
	input wire [16:0] rd_ID;
	input wire rd_ID_valid;
	input wire [16:0] rd_addr;
	input wire rd_addr_valid;
	input wire [16:0] rd_op;
	input wire rd_op_valid;
	input wire rd_rsp_data_ready;
	input wire rst_n;
	input wire tile_en;
	input wire [16:0] wr_ID;
	input wire wr_ID_valid;
	input wire [16:0] wr_addr;
	input wire wr_addr_valid;
	input wire [16:0] wr_data;
	input wire wr_data_valid;
	output wire [8:0] addr_to_mem;
	output wire [63:0] data_to_mem;
	output wire rd_ID_ready;
	output wire rd_addr_ready;
	output wire rd_op_ready;
	output wire [16:0] rd_rsp_data;
	output wire rd_rsp_data_valid;
	output wire ren_to_mem;
	output wire wen_to_mem;
	output wire wr_ID_ready;
	output wire wr_addr_ready;
	output wire wr_data_ready;
	reg PREVIOUS_WR_OP;
	wire [15:0] addr_to_mem_local;
	wire any_sram_lock;
	wire [3:0] base_rr;
	wire [31:0] blk_base;
	wire [31:0] blk_bounds;
	wire [31:0] blk_fifo_0_data_in;
	wire [31:0] blk_fifo_0_data_out;
	wire blk_fifo_0_empty;
	wire blk_fifo_0_full;
	wire [31:0] blk_fifo_1_data_in;
	wire [31:0] blk_fifo_1_data_out;
	wire blk_fifo_1_empty;
	wire blk_fifo_1_full;
	wire [1:0] blk_full;
	wire [1:0] blk_valid;
	wire [31:0] buffet_base;
	wire [31:0] buffet_capacity;
	wire [31:0] buffet_capacity_mask;
	reg [15:0] cached_read_word_addr_0;
	reg [15:0] cached_read_word_addr_1;
	wire [15:0] chosen_read_0;
	wire [15:0] chosen_read_1;
	reg clr_cached_read_0;
	reg clr_cached_read_1;
	reg clr_write_wide_word_0;
	reg clr_write_wide_word_1;
	reg [15:0] curr_base_0;
	reg [15:0] curr_base_1;
	wire [15:0] curr_base_pre_0;
	wire [15:0] curr_base_pre_1;
	reg [15:0] curr_bounds_0;
	reg [15:0] curr_bounds_1;
	reg [31:0] curr_capacity_pre;
	reg [15:0] decode_ret_size_request_full_blk_bounds;
	reg decode_sel_done_size_request_full_blk_bounds;
	reg [1:0] en_curr_base;
	reg [1:0] en_curr_bounds;
	wire first_base_set_0_sticky;
	reg first_base_set_0_was_high;
	wire first_base_set_1_sticky;
	reg first_base_set_1_was_high;
	wire gclk;
	wire joined_in_fifo;
	reg [15:0] last_read_ID;
	reg [1:0] last_read_addr;
	reg [15:0] last_read_addr_wide;
	wire [3:0] mem_acq;
	reg [2:0] num_bits_valid_mask_0_sum;
	reg [2:0] num_bits_valid_mask_1_sum;
	reg [1:0] pop_blk;
	wire pop_in_fifos;
	reg [1:0] pop_in_full;
	reg [1:0] push_blk;
	wire rd_ID_fifo_empty;
	wire rd_ID_fifo_full;
	wire [15:0] rd_ID_fifo_out_data;
	wire rd_ID_fifo_pop;
	wire rd_ID_fifo_valid;
	wire rd_addr_fifo_empty;
	wire rd_addr_fifo_full;
	wire [15:0] rd_addr_fifo_out_addr;
	wire rd_addr_fifo_pop;
	wire rd_addr_fifo_valid;
	wire rd_op_fifo_empty;
	wire rd_op_fifo_full;
	wire [15:0] rd_op_fifo_out_op;
	wire rd_op_fifo_pop;
	wire rd_op_fifo_valid;
	wire rd_rsp_fifo_almost_full;
	wire [16:0] rd_rsp_fifo_data_out;
	wire rd_rsp_fifo_empty;
	wire rd_rsp_fifo_full;
	wire [16:0] rd_rsp_fifo_in_data;
	wire rd_rsp_fifo_push;
	reg [15:0] read_ID_d1;
	reg read_d1;
	reg read_from_sram_write_side_0;
	reg read_from_sram_write_side_1;
	reg read_fsm_0_current_state;
	reg read_fsm_0_next_state;
	reg read_fsm_1_current_state;
	reg read_fsm_1_next_state;
	wire read_joined;
	wire read_pop;
	reg [1:0] read_pop_full;
	reg [63:0] read_wide_word_0;
	reg [63:0] read_wide_word_1;
	wire read_wide_word_valid_sticky_0_sticky;
	reg read_wide_word_valid_sticky_0_was_high;
	wire read_wide_word_valid_sticky_1_sticky;
	reg read_wide_word_valid_sticky_1_was_high;
	reg [1:0] ren_full;
	reg ren_full_delayed_0;
	reg ren_full_delayed_1;
	wire rr_arbiter_resource_ready;
	reg set_cached_read_0;
	reg set_cached_read_1;
	reg set_read_word_addr_0;
	reg set_read_word_addr_1;
	reg set_wide_word_addr_0;
	reg set_wide_word_addr_1;
	reg set_write_wide_word_0;
	reg set_write_wide_word_1;
	reg [1:0] size_request_full;
	reg sram_lock_0;
	reg sram_lock_1;
	wire [15:0] tmp_addr_0;
	wire [15:0] tmp_addr_1;
	wire [15:0] tmp_rd_base;
	wire [15:0] tmp_wr_base;
	wire use_cached_read_0;
	wire use_cached_read_1;
	wire valid_from_mem;
	reg [1:0] wen_full;
	wire wr_ID_fifo_empty;
	wire wr_ID_fifo_full;
	wire [15:0] wr_ID_fifo_out_data;
	wire wr_ID_fifo_pop;
	wire wr_ID_fifo_valid;
	wire wr_addr_fifo_empty;
	wire wr_addr_fifo_full;
	wire [15:0] wr_addr_fifo_out_data;
	wire wr_addr_fifo_pop;
	wire wr_addr_fifo_valid;
	wire [16:0] wr_data_fifo_data_out;
	wire wr_data_fifo_empty;
	wire wr_data_fifo_full;
	wire [15:0] wr_data_fifo_out_data;
	wire wr_data_fifo_out_op;
	wire wr_data_fifo_pop;
	wire wr_data_fifo_valid;
	reg [1:0] write_fsm_0_current_state;
	reg [1:0] write_fsm_0_next_state;
	reg [1:0] write_fsm_1_current_state;
	reg [1:0] write_fsm_1_next_state;
	wire write_full_word_0;
	wire write_full_word_1;
	reg write_to_sram_0;
	reg write_to_sram_1;
	wire [63:0] write_wide_word_comb_in_0;
	wire [63:0] write_wide_word_comb_in_1;
	wire [63:0] write_wide_word_comb_out_0;
	wire [63:0] write_wide_word_comb_out_1;
	wire [3:0] write_wide_word_mask_comb_0;
	wire [3:0] write_wide_word_mask_comb_1;
	wire [3:0] write_wide_word_mask_reg_in_0;
	wire [3:0] write_wide_word_mask_reg_in_1;
	wire [3:0] write_wide_word_mask_reg_out_0;
	wire [3:0] write_wide_word_mask_reg_out_1;
	reg [3:0] write_wide_word_mask_reg_strg_0;
	reg [3:0] write_wide_word_mask_reg_strg_1;
	wire [63:0] write_wide_word_modified_0;
	wire [63:0] write_wide_word_modified_1;
	reg [63:0] write_wide_word_reg_0;
	reg [63:0] write_wide_word_reg_1;
	reg [15:0] write_word_addr_reg_0;
	reg [15:0] write_word_addr_reg_1;
	wire write_word_addr_valid_sticky_0_sticky;
	reg write_word_addr_valid_sticky_0_was_high;
	wire write_word_addr_valid_sticky_1_sticky;
	reg write_word_addr_valid_sticky_1_was_high;
	assign gclk = clk & tile_en;
	assign buffet_capacity_mask[0] = (buffet_capacity_log[0+:4] > 4'h0) & (buffet_capacity_log[0+:4] != 4'h0);
	assign buffet_capacity_mask[1] = (buffet_capacity_log[0+:4] > 4'h1) & (buffet_capacity_log[0+:4] != 4'h0);
	assign buffet_capacity_mask[2] = (buffet_capacity_log[0+:4] > 4'h2) & (buffet_capacity_log[0+:4] != 4'h0);
	assign buffet_capacity_mask[3] = (buffet_capacity_log[0+:4] > 4'h3) & (buffet_capacity_log[0+:4] != 4'h0);
	assign buffet_capacity_mask[4] = (buffet_capacity_log[0+:4] > 4'h4) & (buffet_capacity_log[0+:4] != 4'h0);
	assign buffet_capacity_mask[5] = (buffet_capacity_log[0+:4] > 4'h5) & (buffet_capacity_log[0+:4] != 4'h0);
	assign buffet_capacity_mask[6] = (buffet_capacity_log[0+:4] > 4'h6) & (buffet_capacity_log[0+:4] != 4'h0);
	assign buffet_capacity_mask[7] = (buffet_capacity_log[0+:4] > 4'h7) & (buffet_capacity_log[0+:4] != 4'h0);
	assign buffet_capacity_mask[8] = (buffet_capacity_log[0+:4] > 4'h8) & (buffet_capacity_log[0+:4] != 4'h0);
	assign buffet_capacity_mask[9] = (buffet_capacity_log[0+:4] > 4'h9) & (buffet_capacity_log[0+:4] != 4'h0);
	assign buffet_capacity_mask[10] = (buffet_capacity_log[0+:4] > 4'ha) & (buffet_capacity_log[0+:4] != 4'h0);
	assign buffet_capacity_mask[11] = (buffet_capacity_log[0+:4] > 4'hb) & (buffet_capacity_log[0+:4] != 4'h0);
	assign buffet_capacity_mask[12] = (buffet_capacity_log[0+:4] > 4'hc) & (buffet_capacity_log[0+:4] != 4'h0);
	assign buffet_capacity_mask[13] = (buffet_capacity_log[0+:4] > 4'hd) & (buffet_capacity_log[0+:4] != 4'h0);
	assign buffet_capacity_mask[14] = (buffet_capacity_log[0+:4] > 4'he) & (buffet_capacity_log[0+:4] != 4'h0);
	assign buffet_capacity_mask[15] = (buffet_capacity_log[0+:4] > 4'hf) & (buffet_capacity_log[0+:4] != 4'h0);
	assign buffet_capacity_mask[16] = (buffet_capacity_log[4+:4] > 4'h0) & (buffet_capacity_log[4+:4] != 4'h0);
	assign buffet_capacity_mask[17] = (buffet_capacity_log[4+:4] > 4'h1) & (buffet_capacity_log[4+:4] != 4'h0);
	assign buffet_capacity_mask[18] = (buffet_capacity_log[4+:4] > 4'h2) & (buffet_capacity_log[4+:4] != 4'h0);
	assign buffet_capacity_mask[19] = (buffet_capacity_log[4+:4] > 4'h3) & (buffet_capacity_log[4+:4] != 4'h0);
	assign buffet_capacity_mask[20] = (buffet_capacity_log[4+:4] > 4'h4) & (buffet_capacity_log[4+:4] != 4'h0);
	assign buffet_capacity_mask[21] = (buffet_capacity_log[4+:4] > 4'h5) & (buffet_capacity_log[4+:4] != 4'h0);
	assign buffet_capacity_mask[22] = (buffet_capacity_log[4+:4] > 4'h6) & (buffet_capacity_log[4+:4] != 4'h0);
	assign buffet_capacity_mask[23] = (buffet_capacity_log[4+:4] > 4'h7) & (buffet_capacity_log[4+:4] != 4'h0);
	assign buffet_capacity_mask[24] = (buffet_capacity_log[4+:4] > 4'h8) & (buffet_capacity_log[4+:4] != 4'h0);
	assign buffet_capacity_mask[25] = (buffet_capacity_log[4+:4] > 4'h9) & (buffet_capacity_log[4+:4] != 4'h0);
	assign buffet_capacity_mask[26] = (buffet_capacity_log[4+:4] > 4'ha) & (buffet_capacity_log[4+:4] != 4'h0);
	assign buffet_capacity_mask[27] = (buffet_capacity_log[4+:4] > 4'hb) & (buffet_capacity_log[4+:4] != 4'h0);
	assign buffet_capacity_mask[28] = (buffet_capacity_log[4+:4] > 4'hc) & (buffet_capacity_log[4+:4] != 4'h0);
	assign buffet_capacity_mask[29] = (buffet_capacity_log[4+:4] > 4'hd) & (buffet_capacity_log[4+:4] != 4'h0);
	assign buffet_capacity_mask[30] = (buffet_capacity_log[4+:4] > 4'he) & (buffet_capacity_log[4+:4] != 4'h0);
	assign buffet_capacity_mask[31] = (buffet_capacity_log[4+:4] > 4'hf) & (buffet_capacity_log[4+:4] != 4'h0);
	function automatic [15:0] sv2v_cast_16;
		input reg [15:0] inp;
		sv2v_cast_16 = inp;
	endfunction
	assign buffet_capacity[0+:16] = (buffet_capacity_log[0+:4] == 4'h0 ? 16'h0000 : 16'h0001 << sv2v_cast_16(buffet_capacity_log[0+:4] + 4'h2));
	assign buffet_capacity[16+:16] = (buffet_capacity_log[4+:4] == 4'h0 ? 16'h0000 : 16'h0001 << sv2v_cast_16(buffet_capacity_log[4+:4] + 4'h2));
	assign buffet_base[0+:16] = 16'h0000;
	assign buffet_base[16+:16] = 16'h0100;
	assign {wr_data_fifo_out_op, wr_data_fifo_out_data} = wr_data_fifo_data_out;
	assign wr_data_ready = ~wr_data_fifo_full;
	assign wr_data_fifo_valid = ~wr_data_fifo_empty;
	assign wr_addr_ready = ~wr_addr_fifo_full;
	assign wr_addr_fifo_valid = ~wr_addr_fifo_empty;
	assign wr_ID_ready = ~wr_ID_fifo_full;
	assign wr_ID_fifo_valid = ~wr_ID_fifo_empty;
	assign rd_op_ready = ~rd_op_fifo_full;
	assign rd_op_fifo_valid = ~rd_op_fifo_empty;
	assign rd_addr_ready = ~rd_addr_fifo_full;
	assign rd_addr_fifo_valid = ~rd_addr_fifo_empty;
	assign rd_ID_ready = ~rd_ID_fifo_full;
	assign rd_ID_fifo_valid = ~rd_ID_fifo_empty;
	assign read_joined = (rd_ID_fifo_valid & rd_op_fifo_valid) & rd_addr_fifo_valid;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			curr_bounds_0 <= 16'hffff;
		else if (clk_en) begin
			if (flush)
				curr_bounds_0 <= 16'hffff;
			else if (en_curr_bounds[0])
				curr_bounds_0 <= wr_addr_fifo_out_data;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			curr_bounds_1 <= 16'hffff;
		else if (clk_en) begin
			if (flush)
				curr_bounds_1 <= 16'hffff;
			else if (en_curr_bounds[1])
				curr_bounds_1 <= wr_addr_fifo_out_data;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			first_base_set_0_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				first_base_set_0_was_high <= 1'h0;
			else if (en_curr_base[0])
				first_base_set_0_was_high <= 1'h1;
		end
	assign first_base_set_0_sticky = first_base_set_0_was_high;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			first_base_set_1_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				first_base_set_1_was_high <= 1'h0;
			else if (en_curr_base[1])
				first_base_set_1_was_high <= 1'h1;
		end
	assign first_base_set_1_sticky = first_base_set_1_was_high;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			curr_base_0 <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				curr_base_0 <= 16'h0000;
			else if (en_curr_base[0])
				curr_base_0 <= curr_base_pre_0;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			curr_base_1 <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				curr_base_1 <= 16'h0000;
			else if (en_curr_base[1])
				curr_base_1 <= curr_base_pre_1;
		end
	assign curr_base_pre_0 = (first_base_set_0_sticky ? ((curr_bounds_0 >> 16'h0002) + 16'h0001) + curr_base_0 : 16'h0000);
	assign curr_base_pre_1 = (first_base_set_1_sticky ? ((curr_bounds_1 >> 16'h0002) + 16'h0001) + curr_base_1 : 16'h0000);
	assign addr_to_mem = addr_to_mem_local[8:0];
	assign tmp_addr_0 = ((sv2v_cast_16(wr_addr_fifo_out_data[15:2]) + curr_base_0) & buffet_capacity_mask[0+:16]) + buffet_base[0+:16];
	assign tmp_addr_1 = ((sv2v_cast_16(wr_addr_fifo_out_data[15:2]) + curr_base_1) & buffet_capacity_mask[16+:16]) + buffet_base[16+:16];
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			write_word_addr_reg_0 <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				write_word_addr_reg_0 <= 16'h0000;
			else if (set_wide_word_addr_0)
				write_word_addr_reg_0 <= tmp_addr_0;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			write_word_addr_reg_1 <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				write_word_addr_reg_1 <= 16'h0000;
			else if (set_wide_word_addr_1)
				write_word_addr_reg_1 <= tmp_addr_1;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			write_word_addr_valid_sticky_0_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				write_word_addr_valid_sticky_0_was_high <= 1'h0;
			else if (set_wide_word_addr_0)
				write_word_addr_valid_sticky_0_was_high <= 1'h1;
		end
	assign write_word_addr_valid_sticky_0_sticky = write_word_addr_valid_sticky_0_was_high;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			write_word_addr_valid_sticky_1_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				write_word_addr_valid_sticky_1_was_high <= 1'h0;
			else if (set_wide_word_addr_1)
				write_word_addr_valid_sticky_1_was_high <= 1'h1;
		end
	assign write_word_addr_valid_sticky_1_sticky = write_word_addr_valid_sticky_1_was_high;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			write_wide_word_mask_reg_strg_0 <= 4'h0;
		else if (clk_en) begin
			if (flush)
				write_wide_word_mask_reg_strg_0 <= 4'h0;
			else if (set_write_wide_word_0 | clr_write_wide_word_0)
				write_wide_word_mask_reg_strg_0 <= write_wide_word_mask_reg_in_0;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			write_wide_word_mask_reg_strg_1 <= 4'h0;
		else if (clk_en) begin
			if (flush)
				write_wide_word_mask_reg_strg_1 <= 4'h0;
			else if (set_write_wide_word_1 | clr_write_wide_word_1)
				write_wide_word_mask_reg_strg_1 <= write_wide_word_mask_reg_in_1;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			write_wide_word_reg_0 <= 64'h0000000000000000;
		else if (clk_en) begin
			if (flush)
				write_wide_word_reg_0 <= 64'h0000000000000000;
			else if (set_write_wide_word_0 | clr_write_wide_word_0)
				write_wide_word_reg_0 <= write_wide_word_comb_in_0;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			write_wide_word_reg_1 <= 64'h0000000000000000;
		else if (clk_en) begin
			if (flush)
				write_wide_word_reg_1 <= 64'h0000000000000000;
			else if (set_write_wide_word_1 | clr_write_wide_word_1)
				write_wide_word_reg_1 <= write_wide_word_comb_in_1;
		end
	assign write_wide_word_comb_out_0[0+:16] = (write_wide_word_mask_reg_out_0[0] ? write_wide_word_reg_0[0+:16] : wr_data_fifo_out_data);
	assign write_wide_word_comb_out_0[16+:16] = (write_wide_word_mask_reg_out_0[1] ? write_wide_word_reg_0[16+:16] : wr_data_fifo_out_data);
	assign write_wide_word_comb_out_0[32+:16] = (write_wide_word_mask_reg_out_0[2] ? write_wide_word_reg_0[32+:16] : wr_data_fifo_out_data);
	assign write_wide_word_comb_out_0[48+:16] = (write_wide_word_mask_reg_out_0[3] ? write_wide_word_reg_0[48+:16] : wr_data_fifo_out_data);
	assign write_wide_word_comb_out_1[0+:16] = (write_wide_word_mask_reg_out_1[0] ? write_wide_word_reg_1[0+:16] : wr_data_fifo_out_data);
	assign write_wide_word_comb_out_1[16+:16] = (write_wide_word_mask_reg_out_1[1] ? write_wide_word_reg_1[16+:16] : wr_data_fifo_out_data);
	assign write_wide_word_comb_out_1[32+:16] = (write_wide_word_mask_reg_out_1[2] ? write_wide_word_reg_1[32+:16] : wr_data_fifo_out_data);
	assign write_wide_word_comb_out_1[48+:16] = (write_wide_word_mask_reg_out_1[3] ? write_wide_word_reg_1[48+:16] : wr_data_fifo_out_data);
	assign write_wide_word_comb_in_0[0+:16] = (write_wide_word_mask_reg_out_0[0] & ~clr_write_wide_word_0 ? write_wide_word_reg_0[0+:16] : wr_data_fifo_out_data);
	assign write_wide_word_comb_in_0[16+:16] = (write_wide_word_mask_reg_out_0[1] & ~clr_write_wide_word_0 ? write_wide_word_reg_0[16+:16] : wr_data_fifo_out_data);
	assign write_wide_word_comb_in_0[32+:16] = (write_wide_word_mask_reg_out_0[2] & ~clr_write_wide_word_0 ? write_wide_word_reg_0[32+:16] : wr_data_fifo_out_data);
	assign write_wide_word_comb_in_0[48+:16] = (write_wide_word_mask_reg_out_0[3] & ~clr_write_wide_word_0 ? write_wide_word_reg_0[48+:16] : wr_data_fifo_out_data);
	assign write_wide_word_comb_in_1[0+:16] = (write_wide_word_mask_reg_out_1[0] & ~clr_write_wide_word_1 ? write_wide_word_reg_1[0+:16] : wr_data_fifo_out_data);
	assign write_wide_word_comb_in_1[16+:16] = (write_wide_word_mask_reg_out_1[1] & ~clr_write_wide_word_1 ? write_wide_word_reg_1[16+:16] : wr_data_fifo_out_data);
	assign write_wide_word_comb_in_1[32+:16] = (write_wide_word_mask_reg_out_1[2] & ~clr_write_wide_word_1 ? write_wide_word_reg_1[32+:16] : wr_data_fifo_out_data);
	assign write_wide_word_comb_in_1[48+:16] = (write_wide_word_mask_reg_out_1[3] & ~clr_write_wide_word_1 ? write_wide_word_reg_1[48+:16] : wr_data_fifo_out_data);
	assign write_wide_word_modified_0[0+:16] = (write_wide_word_mask_reg_out_0[0] ? write_wide_word_reg_0[0+:16] : data_from_mem[0+:16]);
	assign write_wide_word_modified_0[16+:16] = (write_wide_word_mask_reg_out_0[1] ? write_wide_word_reg_0[16+:16] : data_from_mem[16+:16]);
	assign write_wide_word_modified_0[32+:16] = (write_wide_word_mask_reg_out_0[2] ? write_wide_word_reg_0[32+:16] : data_from_mem[32+:16]);
	assign write_wide_word_modified_0[48+:16] = (write_wide_word_mask_reg_out_0[3] ? write_wide_word_reg_0[48+:16] : data_from_mem[48+:16]);
	assign write_wide_word_modified_1[0+:16] = (write_wide_word_mask_reg_out_1[0] ? write_wide_word_reg_1[0+:16] : data_from_mem[0+:16]);
	assign write_wide_word_modified_1[16+:16] = (write_wide_word_mask_reg_out_1[1] ? write_wide_word_reg_1[16+:16] : data_from_mem[16+:16]);
	assign write_wide_word_modified_1[32+:16] = (write_wide_word_mask_reg_out_1[2] ? write_wide_word_reg_1[32+:16] : data_from_mem[32+:16]);
	assign write_wide_word_modified_1[48+:16] = (write_wide_word_mask_reg_out_1[3] ? write_wide_word_reg_1[48+:16] : data_from_mem[48+:16]);
	assign write_wide_word_mask_reg_out_0 = write_wide_word_mask_reg_strg_0;
	assign write_wide_word_mask_reg_out_1 = write_wide_word_mask_reg_strg_1;
	function automatic [1:0] sv2v_cast_2;
		input reg [1:0] inp;
		sv2v_cast_2 = inp;
	endfunction
	function automatic [3:0] sv2v_cast_4;
		input reg [3:0] inp;
		sv2v_cast_4 = inp;
	endfunction
	assign write_wide_word_mask_comb_0 = write_wide_word_mask_reg_out_0 | sv2v_cast_4(sv2v_cast_2(((((tmp_addr_0 == write_word_addr_reg_0) & joined_in_fifo) & (1'h1 == wr_data_fifo_out_op)) & (16'h0000 == wr_ID_fifo_out_data) ? 1'h1 : 1'h0)) << wr_addr_fifo_out_data[1:0]);
	assign write_wide_word_mask_comb_1 = write_wide_word_mask_reg_out_1 | sv2v_cast_4(sv2v_cast_2(((((tmp_addr_1 == write_word_addr_reg_1) & joined_in_fifo) & (1'h1 == wr_data_fifo_out_op)) & (16'h0001 == wr_ID_fifo_out_data) ? 1'h1 : 1'h0)) << wr_addr_fifo_out_data[1:0]);
	assign write_wide_word_mask_reg_in_0 = (clr_write_wide_word_0 ? 4'h0 : write_wide_word_mask_reg_out_0) | (((((clr_write_wide_word_0 & (tmp_addr_0 != write_word_addr_reg_0)) | ((tmp_addr_0 == write_word_addr_reg_0) & (~write_full_word_0 | (write_full_word_0 & ~mem_acq[0])))) & (1'h1 == wr_data_fifo_out_op)) & (16'h0000 == wr_ID_fifo_out_data) ? {3'h0, joined_in_fifo} : 4'h0) << sv2v_cast_4(wr_addr_fifo_out_data[1:0]));
	assign write_wide_word_mask_reg_in_1 = (clr_write_wide_word_1 ? 4'h0 : write_wide_word_mask_reg_out_1) | (((((clr_write_wide_word_1 & (tmp_addr_1 != write_word_addr_reg_1)) | ((tmp_addr_1 == write_word_addr_reg_1) & (~write_full_word_1 | (write_full_word_1 & ~mem_acq[2])))) & (1'h1 == wr_data_fifo_out_op)) & (16'h0001 == wr_ID_fifo_out_data) ? {3'h0, joined_in_fifo} : 4'h0) << sv2v_cast_4(wr_addr_fifo_out_data[1:0]));
	function automatic [2:0] sv2v_cast_3;
		input reg [2:0] inp;
		sv2v_cast_3 = inp;
	endfunction
	always @(*) begin
		num_bits_valid_mask_0_sum = 3'h0;
		num_bits_valid_mask_0_sum = num_bits_valid_mask_0_sum + sv2v_cast_3(write_wide_word_mask_comb_0[0]);
		num_bits_valid_mask_0_sum = num_bits_valid_mask_0_sum + sv2v_cast_3(write_wide_word_mask_comb_0[1]);
		num_bits_valid_mask_0_sum = num_bits_valid_mask_0_sum + sv2v_cast_3(write_wide_word_mask_comb_0[2]);
		num_bits_valid_mask_0_sum = num_bits_valid_mask_0_sum + sv2v_cast_3(write_wide_word_mask_comb_0[3]);
	end
	always @(*) begin
		num_bits_valid_mask_1_sum = 3'h0;
		num_bits_valid_mask_1_sum = num_bits_valid_mask_1_sum + sv2v_cast_3(write_wide_word_mask_comb_1[0]);
		num_bits_valid_mask_1_sum = num_bits_valid_mask_1_sum + sv2v_cast_3(write_wide_word_mask_comb_1[1]);
		num_bits_valid_mask_1_sum = num_bits_valid_mask_1_sum + sv2v_cast_3(write_wide_word_mask_comb_1[2]);
		num_bits_valid_mask_1_sum = num_bits_valid_mask_1_sum + sv2v_cast_3(write_wide_word_mask_comb_1[3]);
	end
	assign write_full_word_0 = 3'h4 == num_bits_valid_mask_0_sum;
	assign write_full_word_1 = 3'h4 == num_bits_valid_mask_1_sum;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			read_wide_word_0 <= 64'h0000000000000000;
		else if (clk_en) begin
			if (flush)
				read_wide_word_0 <= 64'h0000000000000000;
			else if (set_cached_read_0)
				read_wide_word_0 <= data_from_mem;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			read_wide_word_1 <= 64'h0000000000000000;
		else if (clk_en) begin
			if (flush)
				read_wide_word_1 <= 64'h0000000000000000;
			else if (set_cached_read_1)
				read_wide_word_1 <= data_from_mem;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			read_wide_word_valid_sticky_0_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				read_wide_word_valid_sticky_0_was_high <= 1'h0;
			else if (clr_cached_read_0)
				read_wide_word_valid_sticky_0_was_high <= 1'h0;
			else if (set_cached_read_0)
				read_wide_word_valid_sticky_0_was_high <= 1'h1;
		end
	assign read_wide_word_valid_sticky_0_sticky = set_cached_read_0 | read_wide_word_valid_sticky_0_was_high;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			read_wide_word_valid_sticky_1_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				read_wide_word_valid_sticky_1_was_high <= 1'h0;
			else if (clr_cached_read_1)
				read_wide_word_valid_sticky_1_was_high <= 1'h0;
			else if (set_cached_read_1)
				read_wide_word_valid_sticky_1_was_high <= 1'h1;
		end
	assign read_wide_word_valid_sticky_1_sticky = set_cached_read_1 | read_wide_word_valid_sticky_1_was_high;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			last_read_addr <= 2'h0;
		else if (clk_en) begin
			if (flush)
				last_read_addr <= 2'h0;
			else if (ren_to_mem)
				last_read_addr <= rd_addr_fifo_out_addr[1:0];
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			last_read_addr_wide <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				last_read_addr_wide <= 16'h0000;
			else if (ren_to_mem)
				last_read_addr_wide <= addr_to_mem_local;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			last_read_ID <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				last_read_ID <= 16'h0000;
			else if (ren_to_mem)
				last_read_ID <= rd_ID_fifo_out_data;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			cached_read_word_addr_0 <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				cached_read_word_addr_0 <= 16'h0000;
			else if (set_read_word_addr_0)
				cached_read_word_addr_0 <= addr_to_mem_local;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			cached_read_word_addr_1 <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				cached_read_word_addr_1 <= 16'h0000;
			else if (set_read_word_addr_1)
				cached_read_word_addr_1 <= addr_to_mem_local;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			ren_full_delayed_0 <= 1'h0;
		else if (clk_en) begin
			if (flush)
				ren_full_delayed_0 <= 1'h0;
			else
				ren_full_delayed_0 <= ren_full[0];
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			ren_full_delayed_1 <= 1'h0;
		else if (clk_en) begin
			if (flush)
				ren_full_delayed_1 <= 1'h0;
			else
				ren_full_delayed_1 <= ren_full[1];
		end
	assign use_cached_read_0 = read_wide_word_valid_sticky_0_sticky & (valid_from_mem & ren_full_delayed_0 ? (16'h0000 == last_read_ID) & (last_read_addr_wide == cached_read_word_addr_0) : ((((16'h0000 == rd_ID_fifo_out_data) & ((((sv2v_cast_16(rd_addr_fifo_out_addr[15:2]) + blk_base[0+:16]) & buffet_capacity_mask[0+:16]) + buffet_base[0+:16]) == cached_read_word_addr_0)) & (16'h0001 == rd_op_fifo_out_op)) & ~valid_from_mem) & read_joined);
	assign use_cached_read_1 = read_wide_word_valid_sticky_1_sticky & (valid_from_mem & ren_full_delayed_1 ? (16'h0001 == last_read_ID) & (last_read_addr_wide == cached_read_word_addr_1) : ((((16'h0001 == rd_ID_fifo_out_data) & ((((sv2v_cast_16(rd_addr_fifo_out_addr[15:2]) + blk_base[16+:16]) & buffet_capacity_mask[16+:16]) + buffet_base[16+:16]) == cached_read_word_addr_1)) & (16'h0001 == rd_op_fifo_out_op)) & ~valid_from_mem) & read_joined);
	assign chosen_read_0 = ((use_cached_read_0 & read_wide_word_valid_sticky_0_sticky) & ~valid_from_mem ? read_wide_word_0[rd_addr_fifo_out_addr[1:0] * 16+:16] : data_from_mem[last_read_addr[1:0] * 16+:16]);
	assign chosen_read_1 = ((use_cached_read_1 & read_wide_word_valid_sticky_1_sticky) & ~valid_from_mem ? read_wide_word_1[rd_addr_fifo_out_addr[1:0] * 16+:16] : data_from_mem[last_read_addr[1:0] * 16+:16]);
	assign any_sram_lock = |{sram_lock_0, sram_lock_1};
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			read_d1 <= 1'h0;
		else if (clk_en) begin
			if (flush)
				read_d1 <= 1'h0;
			else
				read_d1 <= |{mem_acq[1], mem_acq[3]};
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			read_ID_d1 <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				read_ID_d1 <= 16'h0000;
			else if (ren_to_mem)
				read_ID_d1 <= rd_ID_fifo_out_data;
		end
	assign valid_from_mem = read_d1;
	assign rd_rsp_data[0+:17] = rd_rsp_fifo_data_out;
	assign rd_rsp_data_valid = ~rd_rsp_fifo_empty;
	always @(*) begin
		decode_sel_done_size_request_full_blk_bounds = 1'h0;
		decode_ret_size_request_full_blk_bounds = 16'h0000;
		if (~decode_sel_done_size_request_full_blk_bounds & size_request_full[0]) begin
			decode_ret_size_request_full_blk_bounds = blk_bounds[0+:16];
			decode_sel_done_size_request_full_blk_bounds = 1'h1;
		end
		if (~decode_sel_done_size_request_full_blk_bounds & size_request_full[1]) begin
			decode_ret_size_request_full_blk_bounds = blk_bounds[16+:16];
			decode_sel_done_size_request_full_blk_bounds = 1'h1;
		end
	end
	assign rd_rsp_fifo_in_data[15:0] = (use_cached_read_0 & read_wide_word_valid_sticky_0_sticky ? chosen_read_0 : (use_cached_read_1 & read_wide_word_valid_sticky_1_sticky ? chosen_read_1 : decode_ret_size_request_full_blk_bounds + 16'h0001));
	assign rd_rsp_fifo_in_data[16] = (use_cached_read_0 ? 1'h0 : 1'h1);
	assign rd_rsp_fifo_push = (valid_from_mem | |{use_cached_read_0, use_cached_read_1}) | |size_request_full;
	assign joined_in_fifo = (wr_data_fifo_valid & wr_addr_fifo_valid) & wr_ID_fifo_valid;
	assign {wr_addr_fifo_pop, wr_data_fifo_pop, wr_ID_fifo_pop} = {pop_in_fifos, pop_in_fifos, pop_in_fifos};
	assign pop_in_fifos = |pop_in_full;
	assign {rd_ID_fifo_pop, rd_op_fifo_pop, rd_addr_fifo_pop} = {read_pop, read_pop, read_pop};
	assign read_pop = |read_pop_full;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			curr_capacity_pre[0+:16] <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				curr_capacity_pre[0+:16] <= 16'h0000;
			else if (push_blk[0] || pop_blk[0])
				curr_capacity_pre[0+:16] <= (curr_capacity_pre[0+:16] + (push_blk[0] ? blk_bounds[0+:16] : 16'h0000)) - (pop_blk[0] ? blk_bounds[0+:16] : 16'h0000);
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			curr_capacity_pre[16+:16] <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				curr_capacity_pre[16+:16] <= 16'h0000;
			else if (push_blk[1] || pop_blk[1])
				curr_capacity_pre[16+:16] <= (curr_capacity_pre[16+:16] + (push_blk[1] ? blk_bounds[16+:16] : 16'h0000)) - (pop_blk[1] ? blk_bounds[16+:16] : 16'h0000);
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			PREVIOUS_WR_OP <= 1'h0;
		else if (clk_en) begin
			if (flush)
				PREVIOUS_WR_OP <= 1'h0;
			else
				PREVIOUS_WR_OP <= wr_data_fifo_out_op;
		end
	assign blk_fifo_0_data_in = {curr_base_0, curr_bounds_0};
	assign {blk_base[0+:16], blk_bounds[0+:16]} = blk_fifo_0_data_out;
	assign blk_full[0] = blk_fifo_0_full;
	assign blk_valid[0] = ~blk_fifo_0_empty;
	assign blk_fifo_1_data_in = {curr_base_1, curr_bounds_1};
	assign {blk_base[16+:16], blk_bounds[16+:16]} = blk_fifo_1_data_out;
	assign blk_full[1] = blk_fifo_1_full;
	assign blk_valid[1] = ~blk_fifo_1_empty;
	always @(posedge clk or negedge rst_n)
		if (!rst_n)
			read_fsm_0_current_state <= 1'h0;
		else if (clk_en) begin
			if (flush)
				read_fsm_0_current_state <= 1'h0;
			else
				read_fsm_0_current_state <= read_fsm_0_next_state;
		end
	always @(*) begin
		read_fsm_0_next_state = read_fsm_0_current_state;
		case (read_fsm_0_current_state)
			1'h0: read_fsm_0_next_state = 1'h0;
			default:
				;
		endcase
	end
	always @(*)
		case (read_fsm_0_current_state)
			1'h0: begin : read_fsm_0_RD_START_0_Output
				pop_blk[0] = ((rd_op_fifo_out_op == 16'h0000) & read_joined) & (16'h0000 == rd_ID_fifo_out_data);
				ren_full[0] = ((((((rd_op_fifo_out_op == 16'h0001) & ~use_cached_read_0) & read_joined) & ~rd_rsp_fifo_almost_full) & blk_valid[0]) & ((((sv2v_cast_16(rd_addr_fifo_out_addr[15:2]) + blk_base[0+:16]) + buffet_base[0+:16]) != cached_read_word_addr_0) | ~read_wide_word_valid_sticky_0_sticky)) & (16'h0000 == rd_ID_fifo_out_data);
				read_pop_full[0] = ((rd_op_fifo_out_op == 16'h0002 ? ~valid_from_mem & blk_valid[0] : (rd_op_fifo_out_op == 16'h0001 ? (mem_acq[1] | (use_cached_read_0 & ~valid_from_mem)) & ~rd_rsp_fifo_full : 1'h1)) & read_joined) & (16'h0000 == rd_ID_fifo_out_data);
				size_request_full[0] = ((blk_valid[0] & (rd_op_fifo_out_op == 16'h0002)) & read_joined) & (16'h0000 == rd_ID_fifo_out_data);
				set_cached_read_0 = valid_from_mem & (16'h0000 == read_ID_d1);
				clr_cached_read_0 = ((rd_op_fifo_out_op == 16'h0000) & read_joined) & (16'h0000 == rd_ID_fifo_out_data);
				set_read_word_addr_0 = ((ren_full[0] & mem_acq[1]) & (addr_to_mem_local != cached_read_word_addr_0)) & (16'h0000 == rd_ID_fifo_out_data);
			end
			default:
				;
		endcase
	always @(posedge clk or negedge rst_n)
		if (!rst_n)
			read_fsm_1_current_state <= 1'h0;
		else if (clk_en) begin
			if (flush)
				read_fsm_1_current_state <= 1'h0;
			else
				read_fsm_1_current_state <= read_fsm_1_next_state;
		end
	always @(*) begin
		read_fsm_1_next_state = read_fsm_1_current_state;
		case (read_fsm_1_current_state)
			1'h0: read_fsm_1_next_state = 1'h0;
			default:
				;
		endcase
	end
	always @(*)
		case (read_fsm_1_current_state)
			1'h0: begin : read_fsm_1_RD_START_1_Output
				pop_blk[1] = ((rd_op_fifo_out_op == 16'h0000) & read_joined) & (16'h0001 == rd_ID_fifo_out_data);
				ren_full[1] = ((((((rd_op_fifo_out_op == 16'h0001) & ~use_cached_read_1) & read_joined) & ~rd_rsp_fifo_almost_full) & blk_valid[1]) & ((((sv2v_cast_16(rd_addr_fifo_out_addr[15:2]) + blk_base[16+:16]) + buffet_base[16+:16]) != cached_read_word_addr_1) | ~read_wide_word_valid_sticky_1_sticky)) & (16'h0001 == rd_ID_fifo_out_data);
				read_pop_full[1] = ((rd_op_fifo_out_op == 16'h0002 ? ~valid_from_mem & blk_valid[1] : (rd_op_fifo_out_op == 16'h0001 ? (mem_acq[3] | (use_cached_read_1 & ~valid_from_mem)) & ~rd_rsp_fifo_full : 1'h1)) & read_joined) & (16'h0001 == rd_ID_fifo_out_data);
				size_request_full[1] = ((blk_valid[1] & (rd_op_fifo_out_op == 16'h0002)) & read_joined) & (16'h0001 == rd_ID_fifo_out_data);
				set_cached_read_1 = valid_from_mem & (16'h0001 == read_ID_d1);
				clr_cached_read_1 = ((rd_op_fifo_out_op == 16'h0000) & read_joined) & (16'h0001 == rd_ID_fifo_out_data);
				set_read_word_addr_1 = ((ren_full[1] & mem_acq[3]) & (addr_to_mem_local != cached_read_word_addr_1)) & (16'h0001 == rd_ID_fifo_out_data);
			end
			default:
				;
		endcase
	always @(posedge clk or negedge rst_n)
		if (!rst_n)
			write_fsm_0_current_state <= 2'h2;
		else if (clk_en) begin
			if (flush)
				write_fsm_0_current_state <= 2'h2;
			else
				write_fsm_0_current_state <= write_fsm_0_next_state;
		end
	always @(*) begin
		write_fsm_0_next_state = write_fsm_0_current_state;
		case (write_fsm_0_current_state)
			2'h0:
				if (1'h1 == PREVIOUS_WR_OP)
					write_fsm_0_next_state = 2'h1;
				else if ((1'h0 == PREVIOUS_WR_OP) & ~blk_full[0])
					write_fsm_0_next_state = 2'h2;
				else
					write_fsm_0_next_state = 2'h0;
			2'h1:
				if ((((joined_in_fifo & (wr_data_fifo_out_op == 1'h0)) & ~blk_full[0]) & ((write_full_word_0 & mem_acq[0]) | (num_bits_valid_mask_0_sum == 3'h0))) & (16'h0000 == wr_ID_fifo_out_data))
					write_fsm_0_next_state = 2'h2;
				else if (((((joined_in_fifo & (16'h0000 == wr_ID_fifo_out_data)) & mem_acq[0]) & ((1'h0 == wr_data_fifo_out_op) | (((tmp_addr_0 != write_word_addr_reg_0) & write_word_addr_valid_sticky_0_sticky) & (1'h1 == wr_data_fifo_out_op)))) & (num_bits_valid_mask_0_sum > 3'h0)) & ~write_full_word_0)
					write_fsm_0_next_state = 2'h0;
				else
					write_fsm_0_next_state = 2'h1;
			2'h2:
				if (((joined_in_fifo & (wr_data_fifo_out_op == 1'h0)) & (16'h0000 == wr_ID_fifo_out_data)) & tile_en)
					write_fsm_0_next_state = 2'h1;
				else
					write_fsm_0_next_state = 2'h2;
			default: write_fsm_0_next_state = write_fsm_0_current_state;
		endcase
	end
	always @(*)
		case (write_fsm_0_current_state)
			2'h0: begin : write_fsm_0_MODIFY_0_Output
				push_blk[0] = (1'h0 == PREVIOUS_WR_OP) & ~blk_full[0];
				en_curr_base[0] = (1'h0 == PREVIOUS_WR_OP) & ~blk_full[0];
				en_curr_bounds[0] = 1'h0;
				wen_full[0] = ~blk_full[0];
				pop_in_full[0] = ~blk_full[0];
				set_write_wide_word_0 = 1'h0;
				clr_write_wide_word_0 = ~blk_full[0];
				write_to_sram_0 = ~blk_full[0];
				read_from_sram_write_side_0 = 1'h0;
				set_wide_word_addr_0 = 1'h0;
				sram_lock_0 = ~blk_full[0];
			end
			2'h1: begin : write_fsm_0_WRITING_0_Output
				push_blk[0] = (((joined_in_fifo & (wr_data_fifo_out_op == 1'h0)) & ~blk_full[0]) & ((write_full_word_0 & mem_acq[0]) | (num_bits_valid_mask_0_sum == 3'h0))) & (16'h0000 == wr_ID_fifo_out_data);
				en_curr_base[0] = (((joined_in_fifo & (wr_data_fifo_out_op == 1'h0)) & ~blk_full[0]) & ((write_full_word_0 & mem_acq[0]) | (num_bits_valid_mask_0_sum == 3'h0))) & (16'h0000 == wr_ID_fifo_out_data);
				set_write_wide_word_0 = ((((tmp_addr_0 == write_word_addr_reg_0) & write_word_addr_valid_sticky_0_sticky) & joined_in_fifo) & (wr_data_fifo_out_op == 1'h1)) & (16'h0000 == wr_ID_fifo_out_data);
				en_curr_bounds[0] = (((mem_acq[0] | set_write_wide_word_0) & joined_in_fifo) & (wr_data_fifo_out_op == 1'h1)) & (16'h0000 == wr_ID_fifo_out_data);
				wen_full[0] = ((joined_in_fifo & (wr_data_fifo_out_op == 1'h1)) & ((buffet_capacity[0+:16] - curr_capacity_pre[0+:16]) > wr_addr_fifo_out_data)) & (16'h0000 == wr_ID_fifo_out_data);
				clr_write_wide_word_0 = ((((((tmp_addr_0 != write_word_addr_reg_0) | ~write_word_addr_valid_sticky_0_sticky) | (((tmp_addr_0 == write_word_addr_reg_0) & write_word_addr_valid_sticky_0_sticky) & write_full_word_0)) & joined_in_fifo) & (wr_data_fifo_out_op == 1'h1)) & mem_acq[0]) & (16'h0000 == wr_ID_fifo_out_data);
				write_to_sram_0 = ((write_full_word_0 & joined_in_fifo) & ((buffet_capacity[0+:16] - curr_capacity_pre[0+:16]) > wr_addr_fifo_out_data)) & (16'h0000 == wr_ID_fifo_out_data);
				set_wide_word_addr_0 = ((((tmp_addr_0 != write_word_addr_reg_0) | ~write_word_addr_valid_sticky_0_sticky) & joined_in_fifo) & (wr_data_fifo_out_op == 1'h1)) & (16'h0000 == wr_ID_fifo_out_data);
				sram_lock_0 = 1'h0;
				read_from_sram_write_side_0 = (((((joined_in_fifo & (16'h0000 == wr_ID_fifo_out_data)) & ~any_sram_lock) & ((buffet_capacity[0+:16] - curr_capacity_pre[0+:16]) > wr_addr_fifo_out_data)) & ((1'h0 == wr_data_fifo_out_op) | (((tmp_addr_0 != write_word_addr_reg_0) & write_word_addr_valid_sticky_0_sticky) & (1'h1 == wr_data_fifo_out_op)))) & (num_bits_valid_mask_0_sum > 3'h0)) & ~write_full_word_0;
				pop_in_full[0] = (((((mem_acq[0] | set_write_wide_word_0) & joined_in_fifo) & (wr_data_fifo_out_op == 1'h1)) & ((buffet_capacity[0+:16] - curr_capacity_pre[0+:16]) > wr_addr_fifo_out_data)) & (16'h0000 == wr_ID_fifo_out_data)) | ((((joined_in_fifo & (wr_data_fifo_out_op == 1'h0)) & ~blk_full[0]) & ((write_full_word_0 & mem_acq[0]) | (num_bits_valid_mask_0_sum == 3'h0))) & (16'h0000 == wr_ID_fifo_out_data));
			end
			2'h2: begin : write_fsm_0_WR_START_0_Output
				push_blk[0] = 1'h0;
				en_curr_base[0] = 1'h0;
				en_curr_bounds[0] = 1'h0;
				wen_full[0] = 1'h0;
				pop_in_full[0] = (wr_data_fifo_out_op == 1'h0) & (16'h0000 == wr_ID_fifo_out_data);
				set_write_wide_word_0 = 1'h0;
				clr_write_wide_word_0 = 1'h0;
				write_to_sram_0 = 1'h0;
				set_wide_word_addr_0 = 1'h0;
				sram_lock_0 = 1'h0;
				read_from_sram_write_side_0 = 1'h0;
			end
			default: begin : write_fsm_0_default_Output
				push_blk[0] = 1'h0;
				en_curr_base[0] = 1'h0;
				en_curr_bounds[0] = 1'h0;
				wen_full[0] = 1'h0;
				pop_in_full[0] = (wr_data_fifo_out_op == 1'h0) & (16'h0000 == wr_ID_fifo_out_data);
				set_write_wide_word_0 = 1'h0;
				clr_write_wide_word_0 = 1'h0;
				write_to_sram_0 = 1'h0;
				set_wide_word_addr_0 = 1'h0;
				sram_lock_0 = 1'h0;
				read_from_sram_write_side_0 = 1'h0;
			end
		endcase
	always @(posedge clk or negedge rst_n)
		if (!rst_n)
			write_fsm_1_current_state <= 2'h2;
		else if (clk_en) begin
			if (flush)
				write_fsm_1_current_state <= 2'h2;
			else
				write_fsm_1_current_state <= write_fsm_1_next_state;
		end
	always @(*) begin
		write_fsm_1_next_state = write_fsm_1_current_state;
		case (write_fsm_1_current_state)
			2'h0:
				if (1'h1 == PREVIOUS_WR_OP)
					write_fsm_1_next_state = 2'h1;
				else if ((1'h0 == PREVIOUS_WR_OP) & ~blk_full[1])
					write_fsm_1_next_state = 2'h2;
				else
					write_fsm_1_next_state = 2'h0;
			2'h1:
				if ((((joined_in_fifo & (wr_data_fifo_out_op == 1'h0)) & ~blk_full[1]) & ((write_full_word_1 & mem_acq[2]) | (num_bits_valid_mask_1_sum == 3'h0))) & (16'h0001 == wr_ID_fifo_out_data))
					write_fsm_1_next_state = 2'h2;
				else if (((((joined_in_fifo & (16'h0001 == wr_ID_fifo_out_data)) & mem_acq[2]) & ((1'h0 == wr_data_fifo_out_op) | (((tmp_addr_1 != write_word_addr_reg_1) & write_word_addr_valid_sticky_1_sticky) & (1'h1 == wr_data_fifo_out_op)))) & (num_bits_valid_mask_1_sum > 3'h0)) & ~write_full_word_1)
					write_fsm_1_next_state = 2'h0;
				else
					write_fsm_1_next_state = 2'h1;
			2'h2:
				if (((joined_in_fifo & (wr_data_fifo_out_op == 1'h0)) & (16'h0001 == wr_ID_fifo_out_data)) & tile_en)
					write_fsm_1_next_state = 2'h1;
				else
					write_fsm_1_next_state = 2'h2;
			default: write_fsm_1_next_state = write_fsm_1_current_state;
		endcase
	end
	always @(*)
		case (write_fsm_1_current_state)
			2'h0: begin : write_fsm_1_MODIFY_1_Output
				push_blk[1] = (1'h0 == PREVIOUS_WR_OP) & ~blk_full[1];
				en_curr_base[1] = (1'h0 == PREVIOUS_WR_OP) & ~blk_full[1];
				en_curr_bounds[1] = 1'h0;
				wen_full[1] = ~blk_full[1];
				pop_in_full[1] = ~blk_full[1];
				set_write_wide_word_1 = 1'h0;
				clr_write_wide_word_1 = ~blk_full[1];
				write_to_sram_1 = ~blk_full[1];
				read_from_sram_write_side_1 = 1'h0;
				set_wide_word_addr_1 = 1'h0;
				sram_lock_1 = ~blk_full[1];
			end
			2'h1: begin : write_fsm_1_WRITING_1_Output
				push_blk[1] = (((joined_in_fifo & (wr_data_fifo_out_op == 1'h0)) & ~blk_full[1]) & ((write_full_word_1 & mem_acq[2]) | (num_bits_valid_mask_1_sum == 3'h0))) & (16'h0001 == wr_ID_fifo_out_data);
				en_curr_base[1] = (((joined_in_fifo & (wr_data_fifo_out_op == 1'h0)) & ~blk_full[1]) & ((write_full_word_1 & mem_acq[2]) | (num_bits_valid_mask_1_sum == 3'h0))) & (16'h0001 == wr_ID_fifo_out_data);
				set_write_wide_word_1 = ((((tmp_addr_1 == write_word_addr_reg_1) & write_word_addr_valid_sticky_1_sticky) & joined_in_fifo) & (wr_data_fifo_out_op == 1'h1)) & (16'h0001 == wr_ID_fifo_out_data);
				en_curr_bounds[1] = (((mem_acq[2] | set_write_wide_word_1) & joined_in_fifo) & (wr_data_fifo_out_op == 1'h1)) & (16'h0001 == wr_ID_fifo_out_data);
				wen_full[1] = ((joined_in_fifo & (wr_data_fifo_out_op == 1'h1)) & ((buffet_capacity[16+:16] - curr_capacity_pre[16+:16]) > wr_addr_fifo_out_data)) & (16'h0001 == wr_ID_fifo_out_data);
				clr_write_wide_word_1 = ((((((tmp_addr_1 != write_word_addr_reg_1) | ~write_word_addr_valid_sticky_1_sticky) | (((tmp_addr_1 == write_word_addr_reg_1) & write_word_addr_valid_sticky_1_sticky) & write_full_word_1)) & joined_in_fifo) & (wr_data_fifo_out_op == 1'h1)) & mem_acq[2]) & (16'h0001 == wr_ID_fifo_out_data);
				write_to_sram_1 = ((write_full_word_1 & joined_in_fifo) & ((buffet_capacity[16+:16] - curr_capacity_pre[16+:16]) > wr_addr_fifo_out_data)) & (16'h0001 == wr_ID_fifo_out_data);
				set_wide_word_addr_1 = ((((tmp_addr_1 != write_word_addr_reg_1) | ~write_word_addr_valid_sticky_1_sticky) & joined_in_fifo) & (wr_data_fifo_out_op == 1'h1)) & (16'h0001 == wr_ID_fifo_out_data);
				sram_lock_1 = 1'h0;
				read_from_sram_write_side_1 = (((((joined_in_fifo & (16'h0001 == wr_ID_fifo_out_data)) & ~any_sram_lock) & ((buffet_capacity[16+:16] - curr_capacity_pre[16+:16]) > wr_addr_fifo_out_data)) & ((1'h0 == wr_data_fifo_out_op) | (((tmp_addr_1 != write_word_addr_reg_1) & write_word_addr_valid_sticky_1_sticky) & (1'h1 == wr_data_fifo_out_op)))) & (num_bits_valid_mask_1_sum > 3'h0)) & ~write_full_word_1;
				pop_in_full[1] = (((((mem_acq[2] | set_write_wide_word_1) & joined_in_fifo) & (wr_data_fifo_out_op == 1'h1)) & ((buffet_capacity[16+:16] - curr_capacity_pre[16+:16]) > wr_addr_fifo_out_data)) & (16'h0001 == wr_ID_fifo_out_data)) | ((((joined_in_fifo & (wr_data_fifo_out_op == 1'h0)) & ~blk_full[1]) & ((write_full_word_1 & mem_acq[2]) | (num_bits_valid_mask_1_sum == 3'h0))) & (16'h0001 == wr_ID_fifo_out_data));
			end
			2'h2: begin : write_fsm_1_WR_START_1_Output
				push_blk[1] = 1'h0;
				en_curr_base[1] = 1'h0;
				en_curr_bounds[1] = 1'h0;
				wen_full[1] = 1'h0;
				pop_in_full[1] = (wr_data_fifo_out_op == 1'h0) & (16'h0001 == wr_ID_fifo_out_data);
				set_write_wide_word_1 = 1'h0;
				clr_write_wide_word_1 = 1'h0;
				write_to_sram_1 = 1'h0;
				set_wide_word_addr_1 = 1'h0;
				sram_lock_1 = 1'h0;
				read_from_sram_write_side_1 = 1'h0;
			end
			default: begin : write_fsm_1_default_Output
				push_blk[1] = 1'h0;
				en_curr_base[1] = 1'h0;
				en_curr_bounds[1] = 1'h0;
				wen_full[1] = 1'h0;
				pop_in_full[1] = (wr_data_fifo_out_op == 1'h0) & (16'h0001 == wr_ID_fifo_out_data);
				set_write_wide_word_1 = 1'h0;
				clr_write_wide_word_1 = 1'h0;
				write_to_sram_1 = 1'h0;
				set_wide_word_addr_1 = 1'h0;
				sram_lock_1 = 1'h0;
				read_from_sram_write_side_1 = 1'h0;
			end
		endcase
	assign base_rr = {ren_full[1], write_to_sram_1 | read_from_sram_write_side_1, ren_full[0], write_to_sram_0 | read_from_sram_write_side_0};
	assign rr_arbiter_resource_ready = ~any_sram_lock;
	assign ren_to_mem = |{mem_acq[1] & ren_full[0], mem_acq[3] & ren_full[1]} | |{read_from_sram_write_side_0, read_from_sram_write_side_1};
	assign wen_to_mem = |({mem_acq[0] & write_to_sram_0, mem_acq[2] & write_to_sram_1} | {sram_lock_0, sram_lock_1});
	assign tmp_wr_base = (mem_acq[2] & write_to_sram_1 ? curr_base_1 + buffet_base[16+:16] : (mem_acq[0] & write_to_sram_0 ? curr_base_0 + buffet_base[0+:16] : 16'h0000));
	assign tmp_rd_base = (mem_acq[3] & ren_full[1] ? blk_base[16+:16] + buffet_base[16+:16] : (mem_acq[1] & ren_full[0] ? blk_base[0+:16] + buffet_base[0+:16] : 16'h0000));
	assign data_to_mem = (mem_acq[0] & write_to_sram_0 ? write_wide_word_comb_out_0 : (mem_acq[2] & write_to_sram_1 ? write_wide_word_comb_out_1 : (sram_lock_0 ? write_wide_word_modified_0 : (sram_lock_1 ? write_wide_word_modified_1 : 64'h0000000000000000))));
	assign addr_to_mem_local = ((wen_to_mem | mem_acq[0]) | mem_acq[2] ? (mem_acq[0] | sram_lock_0 ? write_word_addr_reg_0 : write_word_addr_reg_1) : (mem_acq[1] & ren_full[0] ? ((sv2v_cast_16(rd_addr_fifo_out_addr[15:2]) + blk_base[0+:16]) & buffet_capacity_mask[0+:16]) + buffet_base[0+:16] : ((sv2v_cast_16(rd_addr_fifo_out_addr[15:2]) + blk_base[16+:16]) & buffet_capacity_mask[16+:16]) + buffet_base[16+:16]));
	reg_fifo_depth_2_w_17_afd_2 wr_data_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(wr_data),
		.flush(flush),
		.pop(wr_data_fifo_pop),
		.push(wr_data_valid),
		.rst_n(rst_n),
		.data_out(wr_data_fifo_data_out),
		.empty(wr_data_fifo_empty),
		.full(wr_data_fifo_full)
	);
	reg_fifo_depth_2_w_16_afd_2 wr_addr_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(wr_addr[15-:16]),
		.flush(flush),
		.pop(wr_addr_fifo_pop),
		.push(wr_addr_valid),
		.rst_n(rst_n),
		.data_out(wr_addr_fifo_out_data),
		.empty(wr_addr_fifo_empty),
		.full(wr_addr_fifo_full)
	);
	reg_fifo_depth_2_w_16_afd_2 wr_ID_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(wr_ID[15-:16]),
		.flush(flush),
		.pop(wr_ID_fifo_pop),
		.push(wr_ID_valid),
		.rst_n(rst_n),
		.data_out(wr_ID_fifo_out_data),
		.empty(wr_ID_fifo_empty),
		.full(wr_ID_fifo_full)
	);
	reg_fifo_depth_2_w_16_afd_2 rd_op_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(rd_op[15-:16]),
		.flush(flush),
		.pop(rd_op_fifo_pop),
		.push(rd_op_valid),
		.rst_n(rst_n),
		.data_out(rd_op_fifo_out_op),
		.empty(rd_op_fifo_empty),
		.full(rd_op_fifo_full)
	);
	reg_fifo_depth_2_w_16_afd_2 rd_addr_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(rd_addr[15-:16]),
		.flush(flush),
		.pop(rd_addr_fifo_pop),
		.push(rd_addr_valid),
		.rst_n(rst_n),
		.data_out(rd_addr_fifo_out_addr),
		.empty(rd_addr_fifo_empty),
		.full(rd_addr_fifo_full)
	);
	reg_fifo_depth_2_w_16_afd_2 rd_ID_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(rd_ID[15-:16]),
		.flush(flush),
		.pop(rd_ID_fifo_pop),
		.push(rd_ID_valid),
		.rst_n(rst_n),
		.data_out(rd_ID_fifo_out_data),
		.empty(rd_ID_fifo_empty),
		.full(rd_ID_fifo_full)
	);
	reg_fifo_depth_2_w_17_afd_1 rd_rsp_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(rd_rsp_fifo_in_data),
		.flush(flush),
		.pop(rd_rsp_data_ready),
		.push(rd_rsp_fifo_push),
		.rst_n(rst_n),
		.almost_full(rd_rsp_fifo_almost_full),
		.data_out(rd_rsp_fifo_data_out),
		.empty(rd_rsp_fifo_empty),
		.full(rd_rsp_fifo_full)
	);
	reg_fifo_depth_2_w_32_afd_2 blk_fifo_0(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(blk_fifo_0_data_in),
		.flush(flush),
		.pop(pop_blk[0]),
		.push(push_blk[0]),
		.rst_n(rst_n),
		.data_out(blk_fifo_0_data_out),
		.empty(blk_fifo_0_empty),
		.full(blk_fifo_0_full)
	);
	reg_fifo_depth_2_w_32_afd_2 blk_fifo_1(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(blk_fifo_1_data_in),
		.flush(flush),
		.pop(pop_blk[1]),
		.push(push_blk[1]),
		.rst_n(rst_n),
		.data_out(blk_fifo_1_data_out),
		.empty(blk_fifo_1_empty),
		.full(blk_fifo_1_full)
	);
	arbiter_4_in_RR_algo rr_arbiter(
		.clk(gclk),
		.clk_en(clk_en),
		.flush(flush),
		.request_in(base_rr),
		.resource_ready(rr_arbiter_resource_ready),
		.rst_n(rst_n),
		.grant_out(mem_acq)
	);
endmodule
module fiber_access_16 (
	buffet_buffet_capacity_log,
	buffet_data_from_mem_lifted,
	buffet_tile_en,
	clk,
	clk_en,
	flush,
	read_scanner_block_mode,
	read_scanner_block_rd_out_ready,
	read_scanner_coord_out_ready,
	read_scanner_dense,
	read_scanner_dim_size,
	read_scanner_do_repeat,
	read_scanner_inner_dim_offset,
	read_scanner_lookup,
	read_scanner_pos_out_ready,
	read_scanner_repeat_factor,
	read_scanner_repeat_outer_inner_n,
	read_scanner_root,
	read_scanner_spacc_mode,
	read_scanner_stop_lvl,
	read_scanner_tile_en,
	read_scanner_us_pos_in,
	read_scanner_us_pos_in_valid,
	rst_n,
	tile_en,
	write_scanner_addr_in,
	write_scanner_addr_in_valid,
	write_scanner_block_mode,
	write_scanner_block_wr_in,
	write_scanner_block_wr_in_valid,
	write_scanner_compressed,
	write_scanner_data_in,
	write_scanner_data_in_valid,
	write_scanner_init_blank,
	write_scanner_lowest_level,
	write_scanner_spacc_mode,
	write_scanner_stop_lvl,
	write_scanner_tile_en,
	buffet_addr_to_mem_lifted,
	buffet_data_to_mem_lifted,
	buffet_ren_to_mem_lifted,
	buffet_wen_to_mem_lifted,
	read_scanner_block_rd_out,
	read_scanner_block_rd_out_valid,
	read_scanner_coord_out,
	read_scanner_coord_out_valid,
	read_scanner_pos_out,
	read_scanner_pos_out_valid,
	read_scanner_us_pos_in_ready,
	write_scanner_addr_in_ready,
	write_scanner_block_wr_in_ready,
	write_scanner_data_in_ready
);
	input wire [7:0] buffet_buffet_capacity_log;
	input wire [63:0] buffet_data_from_mem_lifted;
	input wire buffet_tile_en;
	input wire clk;
	input wire clk_en;
	input wire flush;
	input wire read_scanner_block_mode;
	input wire read_scanner_block_rd_out_ready;
	input wire read_scanner_coord_out_ready;
	input wire read_scanner_dense;
	input wire [15:0] read_scanner_dim_size;
	input wire read_scanner_do_repeat;
	input wire [15:0] read_scanner_inner_dim_offset;
	input wire read_scanner_lookup;
	input wire read_scanner_pos_out_ready;
	input wire [15:0] read_scanner_repeat_factor;
	input wire read_scanner_repeat_outer_inner_n;
	input wire read_scanner_root;
	input wire read_scanner_spacc_mode;
	input wire [15:0] read_scanner_stop_lvl;
	input wire read_scanner_tile_en;
	input wire [16:0] read_scanner_us_pos_in;
	input wire read_scanner_us_pos_in_valid;
	input wire rst_n;
	input wire tile_en;
	input wire [16:0] write_scanner_addr_in;
	input wire write_scanner_addr_in_valid;
	input wire write_scanner_block_mode;
	input wire [16:0] write_scanner_block_wr_in;
	input wire write_scanner_block_wr_in_valid;
	input wire write_scanner_compressed;
	input wire [16:0] write_scanner_data_in;
	input wire write_scanner_data_in_valid;
	input wire write_scanner_init_blank;
	input wire write_scanner_lowest_level;
	input wire write_scanner_spacc_mode;
	input wire [15:0] write_scanner_stop_lvl;
	input wire write_scanner_tile_en;
	output wire [8:0] buffet_addr_to_mem_lifted;
	output wire [63:0] buffet_data_to_mem_lifted;
	output wire buffet_ren_to_mem_lifted;
	output wire buffet_wen_to_mem_lifted;
	output wire [16:0] read_scanner_block_rd_out;
	output wire read_scanner_block_rd_out_valid;
	output wire [16:0] read_scanner_coord_out;
	output wire read_scanner_coord_out_valid;
	output wire [16:0] read_scanner_pos_out;
	output wire read_scanner_pos_out_valid;
	output wire read_scanner_us_pos_in_ready;
	output wire write_scanner_addr_in_ready;
	output wire write_scanner_block_wr_in_ready;
	output wire write_scanner_data_in_ready;
	wire [16:0] buffet_rd_ID;
	wire buffet_rd_ID_ready;
	wire buffet_rd_ID_valid;
	wire [16:0] buffet_rd_addr;
	wire buffet_rd_addr_ready;
	wire buffet_rd_addr_valid;
	wire [16:0] buffet_rd_op;
	wire buffet_rd_op_ready;
	wire buffet_rd_op_valid;
	wire [16:0] buffet_rd_rsp_data;
	wire buffet_rd_rsp_data_ready;
	wire buffet_rd_rsp_data_valid;
	wire [16:0] buffet_wr_ID;
	wire buffet_wr_ID_ready;
	wire buffet_wr_ID_valid;
	wire [16:0] buffet_wr_addr;
	wire buffet_wr_addr_ready;
	wire buffet_wr_addr_valid;
	wire [16:0] buffet_wr_data;
	wire buffet_wr_data_ready;
	wire buffet_wr_data_valid;
	wire gclk;
	assign gclk = clk & tile_en;
	buffet_like_16 buffet(
		.buffet_capacity_log(buffet_buffet_capacity_log),
		.clk(gclk),
		.clk_en(clk_en),
		.data_from_mem(buffet_data_from_mem_lifted),
		.flush(flush),
		.rd_ID(buffet_rd_ID),
		.rd_ID_valid(buffet_rd_ID_valid),
		.rd_addr(buffet_rd_addr),
		.rd_addr_valid(buffet_rd_addr_valid),
		.rd_op(buffet_rd_op),
		.rd_op_valid(buffet_rd_op_valid),
		.rd_rsp_data_ready(buffet_rd_rsp_data_ready),
		.rst_n(rst_n),
		.tile_en(buffet_tile_en),
		.wr_ID(buffet_wr_ID),
		.wr_ID_valid(buffet_wr_ID_valid),
		.wr_addr(buffet_wr_addr),
		.wr_addr_valid(buffet_wr_addr_valid),
		.wr_data(buffet_wr_data),
		.wr_data_valid(buffet_wr_data_valid),
		.addr_to_mem(buffet_addr_to_mem_lifted),
		.data_to_mem(buffet_data_to_mem_lifted),
		.rd_ID_ready(buffet_rd_ID_ready),
		.rd_addr_ready(buffet_rd_addr_ready),
		.rd_op_ready(buffet_rd_op_ready),
		.rd_rsp_data(buffet_rd_rsp_data),
		.rd_rsp_data_valid(buffet_rd_rsp_data_valid),
		.ren_to_mem(buffet_ren_to_mem_lifted),
		.wen_to_mem(buffet_wen_to_mem_lifted),
		.wr_ID_ready(buffet_wr_ID_ready),
		.wr_addr_ready(buffet_wr_addr_ready),
		.wr_data_ready(buffet_wr_data_ready)
	);
	write_scanner write_scanner(
		.ID_out_ready(buffet_wr_ID_ready),
		.addr_in(write_scanner_addr_in),
		.addr_in_valid(write_scanner_addr_in_valid),
		.addr_out_ready(buffet_wr_addr_ready),
		.block_mode(write_scanner_block_mode),
		.block_wr_in(write_scanner_block_wr_in),
		.block_wr_in_valid(write_scanner_block_wr_in_valid),
		.clk(gclk),
		.clk_en(clk_en),
		.compressed(write_scanner_compressed),
		.data_in(write_scanner_data_in),
		.data_in_valid(write_scanner_data_in_valid),
		.data_out_ready(buffet_wr_data_ready),
		.flush(flush),
		.init_blank(write_scanner_init_blank),
		.lowest_level(write_scanner_lowest_level),
		.rst_n(rst_n),
		.spacc_mode(write_scanner_spacc_mode),
		.stop_lvl(write_scanner_stop_lvl),
		.tile_en(write_scanner_tile_en),
		.ID_out(buffet_wr_ID),
		.ID_out_valid(buffet_wr_ID_valid),
		.addr_in_ready(write_scanner_addr_in_ready),
		.addr_out(buffet_wr_addr),
		.addr_out_valid(buffet_wr_addr_valid),
		.block_wr_in_ready(write_scanner_block_wr_in_ready),
		.data_in_ready(write_scanner_data_in_ready),
		.data_out(buffet_wr_data),
		.data_out_valid(buffet_wr_data_valid)
	);
	scanner_pipe read_scanner(
		.ID_out_ready(buffet_rd_ID_ready),
		.addr_out_ready(buffet_rd_addr_ready),
		.block_mode(read_scanner_block_mode),
		.block_rd_out_ready(read_scanner_block_rd_out_ready),
		.clk(gclk),
		.clk_en(clk_en),
		.coord_out_ready(read_scanner_coord_out_ready),
		.dense(read_scanner_dense),
		.dim_size(read_scanner_dim_size),
		.do_repeat(read_scanner_do_repeat),
		.flush(flush),
		.inner_dim_offset(read_scanner_inner_dim_offset),
		.lookup(read_scanner_lookup),
		.op_out_ready(buffet_rd_op_ready),
		.pos_out_ready(read_scanner_pos_out_ready),
		.rd_rsp_data_in(buffet_rd_rsp_data),
		.rd_rsp_data_in_valid(buffet_rd_rsp_data_valid),
		.repeat_factor(read_scanner_repeat_factor),
		.repeat_outer_inner_n(read_scanner_repeat_outer_inner_n),
		.root(read_scanner_root),
		.rst_n(rst_n),
		.spacc_mode(read_scanner_spacc_mode),
		.stop_lvl(read_scanner_stop_lvl),
		.tile_en(read_scanner_tile_en),
		.us_pos_in(read_scanner_us_pos_in),
		.us_pos_in_valid(read_scanner_us_pos_in_valid),
		.ID_out(buffet_rd_ID),
		.ID_out_valid(buffet_rd_ID_valid),
		.addr_out(buffet_rd_addr),
		.addr_out_valid(buffet_rd_addr_valid),
		.block_rd_out(read_scanner_block_rd_out),
		.block_rd_out_valid(read_scanner_block_rd_out_valid),
		.coord_out(read_scanner_coord_out),
		.coord_out_valid(read_scanner_coord_out_valid),
		.op_out(buffet_rd_op),
		.op_out_valid(buffet_rd_op_valid),
		.pos_out(read_scanner_pos_out),
		.pos_out_valid(read_scanner_pos_out_valid),
		.rd_rsp_data_in_ready(buffet_rd_rsp_data_ready),
		.us_pos_in_ready(read_scanner_us_pos_in_ready)
	);
endmodule
module fiber_access_16_flat (
	clk,
	clk_en,
	fiber_access_16_inst_buffet_buffet_capacity_log_0,
	fiber_access_16_inst_buffet_buffet_capacity_log_1,
	fiber_access_16_inst_buffet_data_from_mem_lifted_lifted,
	fiber_access_16_inst_buffet_tile_en,
	fiber_access_16_inst_read_scanner_block_mode,
	fiber_access_16_inst_read_scanner_dense,
	fiber_access_16_inst_read_scanner_dim_size,
	fiber_access_16_inst_read_scanner_do_repeat,
	fiber_access_16_inst_read_scanner_inner_dim_offset,
	fiber_access_16_inst_read_scanner_lookup,
	fiber_access_16_inst_read_scanner_repeat_factor,
	fiber_access_16_inst_read_scanner_repeat_outer_inner_n,
	fiber_access_16_inst_read_scanner_root,
	fiber_access_16_inst_read_scanner_spacc_mode,
	fiber_access_16_inst_read_scanner_stop_lvl,
	fiber_access_16_inst_read_scanner_tile_en,
	fiber_access_16_inst_tile_en,
	fiber_access_16_inst_write_scanner_block_mode,
	fiber_access_16_inst_write_scanner_compressed,
	fiber_access_16_inst_write_scanner_init_blank,
	fiber_access_16_inst_write_scanner_lowest_level,
	fiber_access_16_inst_write_scanner_spacc_mode,
	fiber_access_16_inst_write_scanner_stop_lvl,
	fiber_access_16_inst_write_scanner_tile_en,
	flush,
	read_scanner_block_rd_out_ready_f_,
	read_scanner_coord_out_ready_f_,
	read_scanner_pos_out_ready_f_,
	read_scanner_us_pos_in_f_,
	read_scanner_us_pos_in_valid_f_,
	rst_n,
	write_scanner_addr_in_f_,
	write_scanner_addr_in_valid_f_,
	write_scanner_block_wr_in_f_,
	write_scanner_block_wr_in_valid_f_,
	write_scanner_data_in_f_,
	write_scanner_data_in_valid_f_,
	fiber_access_16_inst_buffet_addr_to_mem_lifted_lifted,
	fiber_access_16_inst_buffet_data_to_mem_lifted_lifted,
	fiber_access_16_inst_buffet_ren_to_mem_lifted_lifted,
	fiber_access_16_inst_buffet_wen_to_mem_lifted_lifted,
	read_scanner_block_rd_out_f_,
	read_scanner_block_rd_out_valid_f_,
	read_scanner_coord_out_f_,
	read_scanner_coord_out_valid_f_,
	read_scanner_pos_out_f_,
	read_scanner_pos_out_valid_f_,
	read_scanner_us_pos_in_ready_f_,
	write_scanner_addr_in_ready_f_,
	write_scanner_block_wr_in_ready_f_,
	write_scanner_data_in_ready_f_
);
	input wire clk;
	input wire clk_en;
	input wire [3:0] fiber_access_16_inst_buffet_buffet_capacity_log_0;
	input wire [3:0] fiber_access_16_inst_buffet_buffet_capacity_log_1;
	input wire [63:0] fiber_access_16_inst_buffet_data_from_mem_lifted_lifted;
	input wire fiber_access_16_inst_buffet_tile_en;
	input wire fiber_access_16_inst_read_scanner_block_mode;
	input wire fiber_access_16_inst_read_scanner_dense;
	input wire [15:0] fiber_access_16_inst_read_scanner_dim_size;
	input wire fiber_access_16_inst_read_scanner_do_repeat;
	input wire [15:0] fiber_access_16_inst_read_scanner_inner_dim_offset;
	input wire fiber_access_16_inst_read_scanner_lookup;
	input wire [15:0] fiber_access_16_inst_read_scanner_repeat_factor;
	input wire fiber_access_16_inst_read_scanner_repeat_outer_inner_n;
	input wire fiber_access_16_inst_read_scanner_root;
	input wire fiber_access_16_inst_read_scanner_spacc_mode;
	input wire [15:0] fiber_access_16_inst_read_scanner_stop_lvl;
	input wire fiber_access_16_inst_read_scanner_tile_en;
	input wire fiber_access_16_inst_tile_en;
	input wire fiber_access_16_inst_write_scanner_block_mode;
	input wire fiber_access_16_inst_write_scanner_compressed;
	input wire fiber_access_16_inst_write_scanner_init_blank;
	input wire fiber_access_16_inst_write_scanner_lowest_level;
	input wire fiber_access_16_inst_write_scanner_spacc_mode;
	input wire [15:0] fiber_access_16_inst_write_scanner_stop_lvl;
	input wire fiber_access_16_inst_write_scanner_tile_en;
	input wire flush;
	input wire read_scanner_block_rd_out_ready_f_;
	input wire read_scanner_coord_out_ready_f_;
	input wire read_scanner_pos_out_ready_f_;
	input wire [16:0] read_scanner_us_pos_in_f_;
	input wire read_scanner_us_pos_in_valid_f_;
	input wire rst_n;
	input wire [16:0] write_scanner_addr_in_f_;
	input wire write_scanner_addr_in_valid_f_;
	input wire [16:0] write_scanner_block_wr_in_f_;
	input wire write_scanner_block_wr_in_valid_f_;
	input wire [16:0] write_scanner_data_in_f_;
	input wire write_scanner_data_in_valid_f_;
	output wire [8:0] fiber_access_16_inst_buffet_addr_to_mem_lifted_lifted;
	output wire [63:0] fiber_access_16_inst_buffet_data_to_mem_lifted_lifted;
	output wire fiber_access_16_inst_buffet_ren_to_mem_lifted_lifted;
	output wire fiber_access_16_inst_buffet_wen_to_mem_lifted_lifted;
	output wire [16:0] read_scanner_block_rd_out_f_;
	output wire read_scanner_block_rd_out_valid_f_;
	output wire [16:0] read_scanner_coord_out_f_;
	output wire read_scanner_coord_out_valid_f_;
	output wire [16:0] read_scanner_pos_out_f_;
	output wire read_scanner_pos_out_valid_f_;
	output wire read_scanner_us_pos_in_ready_f_;
	output wire write_scanner_addr_in_ready_f_;
	output wire write_scanner_block_wr_in_ready_f_;
	output wire write_scanner_data_in_ready_f_;
	wire [7:0] fiber_access_16_inst_buffet_buffet_capacity_log;
	assign fiber_access_16_inst_buffet_buffet_capacity_log[0+:4] = fiber_access_16_inst_buffet_buffet_capacity_log_0;
	assign fiber_access_16_inst_buffet_buffet_capacity_log[4+:4] = fiber_access_16_inst_buffet_buffet_capacity_log_1;
	fiber_access_16 fiber_access_16_inst(
		.buffet_buffet_capacity_log(fiber_access_16_inst_buffet_buffet_capacity_log),
		.buffet_data_from_mem_lifted(fiber_access_16_inst_buffet_data_from_mem_lifted_lifted),
		.buffet_tile_en(fiber_access_16_inst_buffet_tile_en),
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.read_scanner_block_mode(fiber_access_16_inst_read_scanner_block_mode),
		.read_scanner_block_rd_out_ready(read_scanner_block_rd_out_ready_f_),
		.read_scanner_coord_out_ready(read_scanner_coord_out_ready_f_),
		.read_scanner_dense(fiber_access_16_inst_read_scanner_dense),
		.read_scanner_dim_size(fiber_access_16_inst_read_scanner_dim_size),
		.read_scanner_do_repeat(fiber_access_16_inst_read_scanner_do_repeat),
		.read_scanner_inner_dim_offset(fiber_access_16_inst_read_scanner_inner_dim_offset),
		.read_scanner_lookup(fiber_access_16_inst_read_scanner_lookup),
		.read_scanner_pos_out_ready(read_scanner_pos_out_ready_f_),
		.read_scanner_repeat_factor(fiber_access_16_inst_read_scanner_repeat_factor),
		.read_scanner_repeat_outer_inner_n(fiber_access_16_inst_read_scanner_repeat_outer_inner_n),
		.read_scanner_root(fiber_access_16_inst_read_scanner_root),
		.read_scanner_spacc_mode(fiber_access_16_inst_read_scanner_spacc_mode),
		.read_scanner_stop_lvl(fiber_access_16_inst_read_scanner_stop_lvl),
		.read_scanner_tile_en(fiber_access_16_inst_read_scanner_tile_en),
		.read_scanner_us_pos_in(read_scanner_us_pos_in_f_),
		.read_scanner_us_pos_in_valid(read_scanner_us_pos_in_valid_f_),
		.rst_n(rst_n),
		.tile_en(fiber_access_16_inst_tile_en),
		.write_scanner_addr_in(write_scanner_addr_in_f_),
		.write_scanner_addr_in_valid(write_scanner_addr_in_valid_f_),
		.write_scanner_block_mode(fiber_access_16_inst_write_scanner_block_mode),
		.write_scanner_block_wr_in(write_scanner_block_wr_in_f_),
		.write_scanner_block_wr_in_valid(write_scanner_block_wr_in_valid_f_),
		.write_scanner_compressed(fiber_access_16_inst_write_scanner_compressed),
		.write_scanner_data_in(write_scanner_data_in_f_),
		.write_scanner_data_in_valid(write_scanner_data_in_valid_f_),
		.write_scanner_init_blank(fiber_access_16_inst_write_scanner_init_blank),
		.write_scanner_lowest_level(fiber_access_16_inst_write_scanner_lowest_level),
		.write_scanner_spacc_mode(fiber_access_16_inst_write_scanner_spacc_mode),
		.write_scanner_stop_lvl(fiber_access_16_inst_write_scanner_stop_lvl),
		.write_scanner_tile_en(fiber_access_16_inst_write_scanner_tile_en),
		.buffet_addr_to_mem_lifted(fiber_access_16_inst_buffet_addr_to_mem_lifted_lifted),
		.buffet_data_to_mem_lifted(fiber_access_16_inst_buffet_data_to_mem_lifted_lifted),
		.buffet_ren_to_mem_lifted(fiber_access_16_inst_buffet_ren_to_mem_lifted_lifted),
		.buffet_wen_to_mem_lifted(fiber_access_16_inst_buffet_wen_to_mem_lifted_lifted),
		.read_scanner_block_rd_out(read_scanner_block_rd_out_f_),
		.read_scanner_block_rd_out_valid(read_scanner_block_rd_out_valid_f_),
		.read_scanner_coord_out(read_scanner_coord_out_f_),
		.read_scanner_coord_out_valid(read_scanner_coord_out_valid_f_),
		.read_scanner_pos_out(read_scanner_pos_out_f_),
		.read_scanner_pos_out_valid(read_scanner_pos_out_valid_f_),
		.read_scanner_us_pos_in_ready(read_scanner_us_pos_in_ready_f_),
		.write_scanner_addr_in_ready(write_scanner_addr_in_ready_f_),
		.write_scanner_block_wr_in_ready(write_scanner_block_wr_in_ready_f_),
		.write_scanner_data_in_ready(write_scanner_data_in_ready_f_)
	);
endmodule
module for_loop_3_11 (
	clk,
	clk_en,
	dimensionality,
	flush,
	ranges,
	rst_n,
	step,
	mux_sel_out,
	restart
);
	parameter CONFIG_WIDTH = 5'h0b;
	parameter ITERATOR_SUPPORT = 3'h3;
	parameter ITERATOR_SUPPORT2 = 2'h2;
	input wire clk;
	input wire clk_en;
	input wire [2:0] dimensionality;
	input wire flush;
	input wire [32:0] ranges;
	input wire rst_n;
	input wire step;
	output wire [1:0] mux_sel_out;
	output wire restart;
	reg [2:0] clear;
	reg [32:0] dim_counter;
	reg done;
	reg [2:0] inc;
	wire [10:0] inced_cnt;
	reg [2:0] max_value;
	wire maxed_value;
	reg [1:0] mux_sel;
	assign mux_sel_out = mux_sel;
	assign inced_cnt = dim_counter[mux_sel * 11+:11] + 11'h001;
	assign maxed_value = (dim_counter[mux_sel * 11+:11] == ranges[mux_sel * 11+:11]) & inc[mux_sel];
	always @(*) begin
		mux_sel = 2'h0;
		done = 1'h0;
		if (~done) begin
			if (~max_value[0] & (dimensionality > 3'h0)) begin
				mux_sel = 2'h0;
				done = 1'h1;
			end
		end
		if (~done) begin
			if (~max_value[1] & (dimensionality > 3'h1)) begin
				mux_sel = 2'h1;
				done = 1'h1;
			end
		end
		if (~done) begin
			if (~max_value[2] & (dimensionality > 3'h2)) begin
				mux_sel = 2'h2;
				done = 1'h1;
			end
		end
	end
	always @(*) begin
		clear[0] = 1'h0;
		if (((mux_sel > 2'h0) | ~done) & step)
			clear[0] = 1'h1;
	end
	always @(*) begin
		inc[0] = 1'h0;
		if ((1'd1 & step) & (dimensionality > 3'h0))
			inc[0] = 1'h1;
		else if (((mux_sel == 2'h0) & step) & (dimensionality > 3'h0))
			inc[0] = 1'h1;
	end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			dim_counter[0+:11] <= 11'h000;
		else if (clk_en) begin
			if (flush)
				dim_counter[0+:11] <= 11'h000;
			else if (clear[0])
				dim_counter[0+:11] <= 11'h000;
			else if (inc[0])
				dim_counter[0+:11] <= inced_cnt;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			max_value[0] <= 1'h0;
		else if (clk_en) begin
			if (flush)
				max_value[0] <= 1'h0;
			else if (clear[0])
				max_value[0] <= 1'h0;
			else if (inc[0])
				max_value[0] <= maxed_value;
		end
	always @(*) begin
		clear[1] = 1'h0;
		if (((mux_sel > 2'h1) | ~done) & step)
			clear[1] = 1'h1;
	end
	always @(*) begin
		inc[1] = 1'h0;
		if ((1'd0 & step) & (dimensionality > 3'h1))
			inc[1] = 1'h1;
		else if (((mux_sel == 2'h1) & step) & (dimensionality > 3'h1))
			inc[1] = 1'h1;
	end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			dim_counter[11+:11] <= 11'h000;
		else if (clk_en) begin
			if (flush)
				dim_counter[11+:11] <= 11'h000;
			else if (clear[1])
				dim_counter[11+:11] <= 11'h000;
			else if (inc[1])
				dim_counter[11+:11] <= inced_cnt;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			max_value[1] <= 1'h0;
		else if (clk_en) begin
			if (flush)
				max_value[1] <= 1'h0;
			else if (clear[1])
				max_value[1] <= 1'h0;
			else if (inc[1])
				max_value[1] <= maxed_value;
		end
	always @(*) begin
		clear[2] = 1'h0;
		if (((mux_sel > 2'h2) | ~done) & step)
			clear[2] = 1'h1;
	end
	always @(*) begin
		inc[2] = 1'h0;
		if ((1'd0 & step) & (dimensionality > 3'h2))
			inc[2] = 1'h1;
		else if (((mux_sel == 2'h2) & step) & (dimensionality > 3'h2))
			inc[2] = 1'h1;
	end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			dim_counter[22+:11] <= 11'h000;
		else if (clk_en) begin
			if (flush)
				dim_counter[22+:11] <= 11'h000;
			else if (clear[2])
				dim_counter[22+:11] <= 11'h000;
			else if (inc[2])
				dim_counter[22+:11] <= inced_cnt;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			max_value[2] <= 1'h0;
		else if (clk_en) begin
			if (flush)
				max_value[2] <= 1'h0;
			else if (clear[2])
				max_value[2] <= 1'h0;
			else if (inc[2])
				max_value[2] <= maxed_value;
		end
	assign restart = step & ~done;
endmodule
module for_loop_6_11 (
	clk,
	clk_en,
	dimensionality,
	flush,
	ranges,
	rst_n,
	step,
	mux_sel_out,
	restart
);
	parameter CONFIG_WIDTH = 5'h0b;
	parameter ITERATOR_SUPPORT = 4'h6;
	parameter ITERATOR_SUPPORT2 = 2'h2;
	input wire clk;
	input wire clk_en;
	input wire [3:0] dimensionality;
	input wire flush;
	input wire [65:0] ranges;
	input wire rst_n;
	input wire step;
	output wire [2:0] mux_sel_out;
	output wire restart;
	reg [5:0] clear;
	reg [65:0] dim_counter;
	reg done;
	reg [5:0] inc;
	wire [10:0] inced_cnt;
	reg [5:0] max_value;
	wire maxed_value;
	reg [2:0] mux_sel;
	assign mux_sel_out = mux_sel;
	assign inced_cnt = dim_counter[mux_sel * 11+:11] + 11'h001;
	assign maxed_value = (dim_counter[mux_sel * 11+:11] == ranges[mux_sel * 11+:11]) & inc[mux_sel];
	always @(*) begin
		mux_sel = 3'h0;
		done = 1'h0;
		if (~done) begin
			if (~max_value[0] & (dimensionality > 4'h0)) begin
				mux_sel = 3'h0;
				done = 1'h1;
			end
		end
		if (~done) begin
			if (~max_value[1] & (dimensionality > 4'h1)) begin
				mux_sel = 3'h1;
				done = 1'h1;
			end
		end
		if (~done) begin
			if (~max_value[2] & (dimensionality > 4'h2)) begin
				mux_sel = 3'h2;
				done = 1'h1;
			end
		end
		if (~done) begin
			if (~max_value[3] & (dimensionality > 4'h3)) begin
				mux_sel = 3'h3;
				done = 1'h1;
			end
		end
		if (~done) begin
			if (~max_value[4] & (dimensionality > 4'h4)) begin
				mux_sel = 3'h4;
				done = 1'h1;
			end
		end
		if (~done) begin
			if (~max_value[5] & (dimensionality > 4'h5)) begin
				mux_sel = 3'h5;
				done = 1'h1;
			end
		end
	end
	always @(*) begin
		clear[0] = 1'h0;
		if (((mux_sel > 3'h0) | ~done) & step)
			clear[0] = 1'h1;
	end
	always @(*) begin
		inc[0] = 1'h0;
		if ((1'd1 & step) & (dimensionality > 4'h0))
			inc[0] = 1'h1;
		else if (((mux_sel == 3'h0) & step) & (dimensionality > 4'h0))
			inc[0] = 1'h1;
	end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			dim_counter[0+:11] <= 11'h000;
		else if (clk_en) begin
			if (flush)
				dim_counter[0+:11] <= 11'h000;
			else if (clear[0])
				dim_counter[0+:11] <= 11'h000;
			else if (inc[0])
				dim_counter[0+:11] <= inced_cnt;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			max_value[0] <= 1'h0;
		else if (clk_en) begin
			if (flush)
				max_value[0] <= 1'h0;
			else if (clear[0])
				max_value[0] <= 1'h0;
			else if (inc[0])
				max_value[0] <= maxed_value;
		end
	always @(*) begin
		clear[1] = 1'h0;
		if (((mux_sel > 3'h1) | ~done) & step)
			clear[1] = 1'h1;
	end
	always @(*) begin
		inc[1] = 1'h0;
		if ((1'd0 & step) & (dimensionality > 4'h1))
			inc[1] = 1'h1;
		else if (((mux_sel == 3'h1) & step) & (dimensionality > 4'h1))
			inc[1] = 1'h1;
	end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			dim_counter[11+:11] <= 11'h000;
		else if (clk_en) begin
			if (flush)
				dim_counter[11+:11] <= 11'h000;
			else if (clear[1])
				dim_counter[11+:11] <= 11'h000;
			else if (inc[1])
				dim_counter[11+:11] <= inced_cnt;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			max_value[1] <= 1'h0;
		else if (clk_en) begin
			if (flush)
				max_value[1] <= 1'h0;
			else if (clear[1])
				max_value[1] <= 1'h0;
			else if (inc[1])
				max_value[1] <= maxed_value;
		end
	always @(*) begin
		clear[2] = 1'h0;
		if (((mux_sel > 3'h2) | ~done) & step)
			clear[2] = 1'h1;
	end
	always @(*) begin
		inc[2] = 1'h0;
		if ((1'd0 & step) & (dimensionality > 4'h2))
			inc[2] = 1'h1;
		else if (((mux_sel == 3'h2) & step) & (dimensionality > 4'h2))
			inc[2] = 1'h1;
	end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			dim_counter[22+:11] <= 11'h000;
		else if (clk_en) begin
			if (flush)
				dim_counter[22+:11] <= 11'h000;
			else if (clear[2])
				dim_counter[22+:11] <= 11'h000;
			else if (inc[2])
				dim_counter[22+:11] <= inced_cnt;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			max_value[2] <= 1'h0;
		else if (clk_en) begin
			if (flush)
				max_value[2] <= 1'h0;
			else if (clear[2])
				max_value[2] <= 1'h0;
			else if (inc[2])
				max_value[2] <= maxed_value;
		end
	always @(*) begin
		clear[3] = 1'h0;
		if (((mux_sel > 3'h3) | ~done) & step)
			clear[3] = 1'h1;
	end
	always @(*) begin
		inc[3] = 1'h0;
		if ((1'd0 & step) & (dimensionality > 4'h3))
			inc[3] = 1'h1;
		else if (((mux_sel == 3'h3) & step) & (dimensionality > 4'h3))
			inc[3] = 1'h1;
	end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			dim_counter[33+:11] <= 11'h000;
		else if (clk_en) begin
			if (flush)
				dim_counter[33+:11] <= 11'h000;
			else if (clear[3])
				dim_counter[33+:11] <= 11'h000;
			else if (inc[3])
				dim_counter[33+:11] <= inced_cnt;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			max_value[3] <= 1'h0;
		else if (clk_en) begin
			if (flush)
				max_value[3] <= 1'h0;
			else if (clear[3])
				max_value[3] <= 1'h0;
			else if (inc[3])
				max_value[3] <= maxed_value;
		end
	always @(*) begin
		clear[4] = 1'h0;
		if (((mux_sel > 3'h4) | ~done) & step)
			clear[4] = 1'h1;
	end
	always @(*) begin
		inc[4] = 1'h0;
		if ((1'd0 & step) & (dimensionality > 4'h4))
			inc[4] = 1'h1;
		else if (((mux_sel == 3'h4) & step) & (dimensionality > 4'h4))
			inc[4] = 1'h1;
	end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			dim_counter[44+:11] <= 11'h000;
		else if (clk_en) begin
			if (flush)
				dim_counter[44+:11] <= 11'h000;
			else if (clear[4])
				dim_counter[44+:11] <= 11'h000;
			else if (inc[4])
				dim_counter[44+:11] <= inced_cnt;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			max_value[4] <= 1'h0;
		else if (clk_en) begin
			if (flush)
				max_value[4] <= 1'h0;
			else if (clear[4])
				max_value[4] <= 1'h0;
			else if (inc[4])
				max_value[4] <= maxed_value;
		end
	always @(*) begin
		clear[5] = 1'h0;
		if (((mux_sel > 3'h5) | ~done) & step)
			clear[5] = 1'h1;
	end
	always @(*) begin
		inc[5] = 1'h0;
		if ((1'd0 & step) & (dimensionality > 4'h5))
			inc[5] = 1'h1;
		else if (((mux_sel == 3'h5) & step) & (dimensionality > 4'h5))
			inc[5] = 1'h1;
	end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			dim_counter[55+:11] <= 11'h000;
		else if (clk_en) begin
			if (flush)
				dim_counter[55+:11] <= 11'h000;
			else if (clear[5])
				dim_counter[55+:11] <= 11'h000;
			else if (inc[5])
				dim_counter[55+:11] <= inced_cnt;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			max_value[5] <= 1'h0;
		else if (clk_en) begin
			if (flush)
				max_value[5] <= 1'h0;
			else if (clear[5])
				max_value[5] <= 1'h0;
			else if (inc[5])
				max_value[5] <= maxed_value;
		end
	assign restart = step & ~done;
endmodule
module reg_fifo_depth_0_w_16_afd_2 (
	clk,
	clk_en,
	data_in,
	flush,
	pop,
	push,
	rst_n,
	almost_full,
	data_out,
	empty,
	full,
	valid
);
	input wire clk;
	input wire clk_en;
	input wire [15:0] data_in;
	input wire flush;
	input wire pop;
	input wire push;
	input wire rst_n;
	output wire almost_full;
	output wire [15:0] data_out;
	output wire empty;
	output wire full;
	output wire valid;
	assign data_out = data_in;
	assign valid = push;
	assign empty = ~push;
	assign full = ~pop;
	assign almost_full = ~pop;
endmodule
module reg_fifo_depth_2_w_16_afd_2 (
	clk,
	clk_en,
	data_in,
	flush,
	pop,
	push,
	rst_n,
	almost_full,
	data_out,
	empty,
	full,
	valid
);
	input wire clk;
	input wire clk_en;
	input wire [15:0] data_in;
	input wire flush;
	input wire pop;
	input wire push;
	input wire rst_n;
	output wire almost_full;
	output reg [15:0] data_out;
	output wire empty;
	output wire full;
	output reg valid;
	reg [1:0] num_items;
	wire passthru;
	reg rd_ptr;
	wire read;
	reg [31:0] reg_array;
	reg wr_ptr;
	wire write;
	assign full = num_items == 2'h2;
	assign almost_full = num_items >= 2'h0;
	assign empty = num_items == 2'h0;
	assign read = (pop & ~passthru) & ~empty;
	assign passthru = 1'h0;
	assign write = (push & ~passthru) & ~full;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			num_items <= 2'h0;
		else if (flush)
			num_items <= 2'h0;
		else if (clk_en) begin
			if (write & ~read)
				num_items <= num_items + 2'h1;
			else if (~write & read)
				num_items <= num_items - 2'h1;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			reg_array <= 32'h00000000;
		else if (flush)
			reg_array <= 32'h00000000;
		else if (clk_en) begin
			if (write)
				reg_array[16 * wr_ptr+:16] <= data_in;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			wr_ptr <= 1'h0;
		else if (flush)
			wr_ptr <= 1'h0;
		else if (clk_en) begin
			if (write) begin
				if (wr_ptr == 1'h1)
					wr_ptr <= 1'h0;
				else
					wr_ptr <= wr_ptr + 1'h1;
			end
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			rd_ptr <= 1'h0;
		else if (flush)
			rd_ptr <= 1'h0;
		else if (clk_en) begin
			if (read)
				rd_ptr <= rd_ptr + 1'h1;
		end
	always @(*)
		if (passthru)
			data_out = data_in;
		else
			data_out = reg_array[16 * rd_ptr+:16];
	always @(*) valid = ~empty | passthru;
endmodule
module reg_fifo_depth_2_w_17_afd_1 (
	clk,
	clk_en,
	data_in,
	flush,
	pop,
	push,
	rst_n,
	almost_full,
	data_out,
	empty,
	full,
	valid
);
	input wire clk;
	input wire clk_en;
	input wire [16:0] data_in;
	input wire flush;
	input wire pop;
	input wire push;
	input wire rst_n;
	output wire almost_full;
	output reg [16:0] data_out;
	output wire empty;
	output wire full;
	output reg valid;
	reg [1:0] num_items;
	wire passthru;
	reg rd_ptr;
	wire read;
	reg [33:0] reg_array;
	reg wr_ptr;
	wire write;
	assign full = num_items == 2'h2;
	assign almost_full = num_items >= 2'h1;
	assign empty = num_items == 2'h0;
	assign read = (pop & ~passthru) & ~empty;
	assign passthru = 1'h0;
	assign write = (push & ~passthru) & ~full;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			num_items <= 2'h0;
		else if (flush)
			num_items <= 2'h0;
		else if (clk_en) begin
			if (write & ~read)
				num_items <= num_items + 2'h1;
			else if (~write & read)
				num_items <= num_items - 2'h1;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			reg_array <= 34'h000000000;
		else if (flush)
			reg_array <= 34'h000000000;
		else if (clk_en) begin
			if (write)
				reg_array[17 * wr_ptr+:17] <= data_in;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			wr_ptr <= 1'h0;
		else if (flush)
			wr_ptr <= 1'h0;
		else if (clk_en) begin
			if (write) begin
				if (wr_ptr == 1'h1)
					wr_ptr <= 1'h0;
				else
					wr_ptr <= wr_ptr + 1'h1;
			end
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			rd_ptr <= 1'h0;
		else if (flush)
			rd_ptr <= 1'h0;
		else if (clk_en) begin
			if (read)
				rd_ptr <= rd_ptr + 1'h1;
		end
	always @(*)
		if (passthru)
			data_out = data_in;
		else
			data_out = reg_array[17 * rd_ptr+:17];
	always @(*) valid = ~empty | passthru;
endmodule
module reg_fifo_depth_2_w_32_afd_2 (
	clk,
	clk_en,
	data_in,
	flush,
	pop,
	push,
	rst_n,
	almost_full,
	data_out,
	empty,
	full,
	valid
);
	input wire clk;
	input wire clk_en;
	input wire [31:0] data_in;
	input wire flush;
	input wire pop;
	input wire push;
	input wire rst_n;
	output wire almost_full;
	output reg [31:0] data_out;
	output wire empty;
	output wire full;
	output reg valid;
	reg [1:0] num_items;
	wire passthru;
	reg rd_ptr;
	wire read;
	reg [63:0] reg_array;
	reg wr_ptr;
	wire write;
	assign full = num_items == 2'h2;
	assign almost_full = num_items >= 2'h0;
	assign empty = num_items == 2'h0;
	assign read = (pop & ~passthru) & ~empty;
	assign passthru = 1'h0;
	assign write = (push & ~passthru) & ~full;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			num_items <= 2'h0;
		else if (flush)
			num_items <= 2'h0;
		else if (clk_en) begin
			if (clk_en) begin
				if (clk_en) begin
					if (write & ~read)
						num_items <= num_items + 2'h1;
					else if (~write & read)
						num_items <= num_items - 2'h1;
				end
			end
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			reg_array <= 64'h0000000000000000;
		else if (flush)
			reg_array <= 64'h0000000000000000;
		else if (clk_en) begin
			if (clk_en) begin
				if (clk_en) begin
					if (write)
						reg_array[32 * wr_ptr+:32] <= data_in;
				end
			end
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			wr_ptr <= 1'h0;
		else if (flush)
			wr_ptr <= 1'h0;
		else if (clk_en) begin
			if (clk_en) begin
				if (clk_en) begin
					if (write) begin
						if (wr_ptr == 1'h1)
							wr_ptr <= 1'h0;
						else
							wr_ptr <= wr_ptr + 1'h1;
					end
				end
			end
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			rd_ptr <= 1'h0;
		else if (flush)
			rd_ptr <= 1'h0;
		else if (clk_en) begin
			if (clk_en) begin
				if (clk_en) begin
					if (read)
						rd_ptr <= rd_ptr + 1'h1;
				end
			end
		end
	always @(*)
		if (passthru)
			data_out = data_in;
		else
			data_out = reg_array[32 * rd_ptr+:32];
	always @(*) valid = ~empty | passthru;
endmodule
module reservation_fifo_depth_8_w_17_num_per_1 (
	clk,
	clk_en,
	data_in_0,
	fill_data_in,
	flush,
	pop,
	push_alloc,
	push_fill,
	push_reserve,
	rst_n,
	data_out_0,
	empty,
	full,
	valid
);
	input wire clk;
	input wire clk_en;
	input wire [16:0] data_in_0;
	input wire [16:0] fill_data_in;
	input wire flush;
	input wire pop;
	input wire push_alloc;
	input wire push_fill;
	input wire push_reserve;
	input wire rst_n;
	output wire [16:0] data_out_0;
	output wire empty;
	output wire full;
	output reg valid;
	wire clr_item_ptr;
	wire clr_read_ptr;
	wire clr_write_ptr;
	wire [16:0] data_in_packed;
	reg [16:0] data_out;
	wire enable_reserve_ptr;
	wire inc_item_ptr;
	wire inc_read_ptr;
	wire inc_reserve_count;
	wire inc_write_ptr;
	wire item_ptr;
	wire jump_next_0;
	wire [2:0] next_0_valid;
	reg [2:0] next_0_valid_d1;
	reg [2:0] next_0_valid_high;
	reg next_0_valid_high_done;
	reg next_0_valid_high_found;
	reg [2:0] next_0_valid_low;
	reg next_0_valid_low_done;
	reg next_0_valid_low_found;
	reg [3:0] num_items;
	wire read;
	reg [2:0] read_ptr_addr;
	reg [135:0] reg_array;
	reg [15:0] reserve_count;
	wire [2:0] reserve_ptr_val;
	reg [7:0] valid_mask;
	wire write_alloc;
	wire write_fill;
	reg [2:0] write_ptr_addr;
	wire write_reserve;
	wire write_reserve_final;
	assign data_in_packed[0+:17] = data_in_0;
	assign data_out_0 = data_out[0+:17];
	assign item_ptr = 1'h0;
	assign inc_item_ptr = push_reserve;
	assign clr_item_ptr = push_reserve & (item_ptr == 1'h0);
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			read_ptr_addr <= 3'h0;
		else if (flush)
			read_ptr_addr <= 3'h0;
		else if (clk_en) begin
			if (clk_en) begin
				if (clr_read_ptr)
					read_ptr_addr <= 3'h0;
				else if (inc_read_ptr)
					read_ptr_addr <= read_ptr_addr + 3'h1;
			end
		end
	assign inc_read_ptr = read;
	assign clr_read_ptr = 1'h0;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			write_ptr_addr <= 3'h0;
		else if (flush)
			write_ptr_addr <= 3'h0;
		else if (clk_en) begin
			if (clk_en) begin
				if (clr_write_ptr)
					write_ptr_addr <= 3'h0;
				else if (inc_write_ptr)
					write_ptr_addr <= write_ptr_addr + 3'h1;
			end
		end
	assign inc_write_ptr = write_alloc | write_fill;
	assign clr_write_ptr = 1'h0;
	assign jump_next_0 = next_0_valid_high_found | next_0_valid_low_found;
	assign enable_reserve_ptr = write_reserve_final | (write_fill & (reserve_ptr_val == write_ptr_addr));
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			next_0_valid_d1 <= 3'h0;
		else if (flush)
			next_0_valid_d1 <= 3'h0;
		else if (clk_en) begin
			if (clk_en) begin
				if (enable_reserve_ptr)
					next_0_valid_d1 <= next_0_valid;
			end
		end
	assign reserve_ptr_val = next_0_valid_d1;
	assign next_0_valid = (write_fill & (((next_0_valid_d1 == write_ptr_addr) | (~next_0_valid_high_found & ~next_0_valid_low_found)) | (next_0_valid_high_found ? next_0_valid_high == write_ptr_addr : next_0_valid_low == write_ptr_addr)) ? write_ptr_addr + 3'h1 : (~next_0_valid_high_found & ~next_0_valid_low_found ? write_ptr_addr : (next_0_valid_high_found ? next_0_valid_high : next_0_valid_low)));
	assign full = num_items == 4'h8;
	assign empty = num_items == 4'h0;
	assign write_fill = (push_fill & push_alloc) & ~full;
	assign write_alloc = push_alloc & ~full;
	assign write_reserve = inc_item_ptr;
	assign write_reserve_final = clr_item_ptr;
	assign read = pop & valid_mask[read_ptr_addr];
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			num_items <= 4'h0;
		else if (flush)
			num_items <= 4'h0;
		else if (clk_en) begin
			if (clk_en) begin
				if (write_alloc & ~read)
					num_items <= num_items + 4'h1;
				else if (~write_alloc & read)
					num_items <= num_items - 4'h1;
			end
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			reg_array <= 136'h0000000000000000000000000000000000;
		else if (flush)
			reg_array <= 136'h0000000000000000000000000000000000;
		else if (clk_en) begin
			if (clk_en) begin
				if (write_fill)
					reg_array[17 * write_ptr_addr+:17] <= fill_data_in;
				if (write_reserve)
					reg_array[17 * next_0_valid_d1+:17] <= data_in_packed;
			end
		end
	always @(*) data_out = reg_array[17 * read_ptr_addr+:17];
	always @(*) valid = valid_mask[read_ptr_addr];
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			valid_mask <= 8'h00;
		else if (flush)
			valid_mask <= 8'h00;
		else if (clk_en) begin
			if (clk_en) begin
				if (write_fill)
					valid_mask[write_ptr_addr] <= 1'h1;
				if (write_reserve_final)
					valid_mask[next_0_valid_d1] <= 1'h1;
				if (read)
					valid_mask[read_ptr_addr] <= 1'h0;
			end
		end
	always @(*) begin
		next_0_valid_high_found = 1'h0;
		next_0_valid_high = 3'h0;
		next_0_valid_high_done = 1'h0;
		if (~next_0_valid_high_done) begin
			if (next_0_valid_d1 < 3'h0) begin
				if (valid_mask[0] == 1'h0) begin
					next_0_valid_high_found = 1'h1;
					next_0_valid_high = 3'h0;
					next_0_valid_high_done = 1'h1;
				end
			end
		end
		if (~next_0_valid_high_done) begin
			if (next_0_valid_d1 < 3'h1) begin
				if (valid_mask[1] == 1'h0) begin
					next_0_valid_high_found = 1'h1;
					next_0_valid_high = 3'h1;
					next_0_valid_high_done = 1'h1;
				end
			end
		end
		if (~next_0_valid_high_done) begin
			if (next_0_valid_d1 < 3'h2) begin
				if (valid_mask[2] == 1'h0) begin
					next_0_valid_high_found = 1'h1;
					next_0_valid_high = 3'h2;
					next_0_valid_high_done = 1'h1;
				end
			end
		end
		if (~next_0_valid_high_done) begin
			if (next_0_valid_d1 < 3'h3) begin
				if (valid_mask[3] == 1'h0) begin
					next_0_valid_high_found = 1'h1;
					next_0_valid_high = 3'h3;
					next_0_valid_high_done = 1'h1;
				end
			end
		end
		if (~next_0_valid_high_done) begin
			if (next_0_valid_d1 < 3'h4) begin
				if (valid_mask[4] == 1'h0) begin
					next_0_valid_high_found = 1'h1;
					next_0_valid_high = 3'h4;
					next_0_valid_high_done = 1'h1;
				end
			end
		end
		if (~next_0_valid_high_done) begin
			if (next_0_valid_d1 < 3'h5) begin
				if (valid_mask[5] == 1'h0) begin
					next_0_valid_high_found = 1'h1;
					next_0_valid_high = 3'h5;
					next_0_valid_high_done = 1'h1;
				end
			end
		end
		if (~next_0_valid_high_done) begin
			if (next_0_valid_d1 < 3'h6) begin
				if (valid_mask[6] == 1'h0) begin
					next_0_valid_high_found = 1'h1;
					next_0_valid_high = 3'h6;
					next_0_valid_high_done = 1'h1;
				end
			end
		end
		if (~next_0_valid_high_done) begin
			if (next_0_valid_d1 < 3'h7) begin
				if (valid_mask[7] == 1'h0) begin
					next_0_valid_high_found = 1'h1;
					next_0_valid_high = 3'h7;
					next_0_valid_high_done = 1'h1;
				end
			end
		end
	end
	always @(*) begin
		next_0_valid_low_found = 1'h0;
		next_0_valid_low = 3'h0;
		next_0_valid_low_done = 1'h0;
		if (~next_0_valid_low_done) begin
			if (next_0_valid_d1 > 3'h0) begin
				if (valid_mask[0] == 1'h0) begin
					next_0_valid_low_found = 1'h1;
					next_0_valid_low = 3'h0;
					next_0_valid_low_done = 1'h1;
				end
			end
		end
		if (~next_0_valid_low_done) begin
			if (next_0_valid_d1 > 3'h1) begin
				if (valid_mask[1] == 1'h0) begin
					next_0_valid_low_found = 1'h1;
					next_0_valid_low = 3'h1;
					next_0_valid_low_done = 1'h1;
				end
			end
		end
		if (~next_0_valid_low_done) begin
			if (next_0_valid_d1 > 3'h2) begin
				if (valid_mask[2] == 1'h0) begin
					next_0_valid_low_found = 1'h1;
					next_0_valid_low = 3'h2;
					next_0_valid_low_done = 1'h1;
				end
			end
		end
		if (~next_0_valid_low_done) begin
			if (next_0_valid_d1 > 3'h3) begin
				if (valid_mask[3] == 1'h0) begin
					next_0_valid_low_found = 1'h1;
					next_0_valid_low = 3'h3;
					next_0_valid_low_done = 1'h1;
				end
			end
		end
		if (~next_0_valid_low_done) begin
			if (next_0_valid_d1 > 3'h4) begin
				if (valid_mask[4] == 1'h0) begin
					next_0_valid_low_found = 1'h1;
					next_0_valid_low = 3'h4;
					next_0_valid_low_done = 1'h1;
				end
			end
		end
		if (~next_0_valid_low_done) begin
			if (next_0_valid_d1 > 3'h5) begin
				if (valid_mask[5] == 1'h0) begin
					next_0_valid_low_found = 1'h1;
					next_0_valid_low = 3'h5;
					next_0_valid_low_done = 1'h1;
				end
			end
		end
		if (~next_0_valid_low_done) begin
			if (next_0_valid_d1 > 3'h6) begin
				if (valid_mask[6] == 1'h0) begin
					next_0_valid_low_found = 1'h1;
					next_0_valid_low = 3'h6;
					next_0_valid_low_done = 1'h1;
				end
			end
		end
		if (~next_0_valid_low_done) begin
			if (next_0_valid_d1 > 3'h7) begin
				if (valid_mask[7] == 1'h0) begin
					next_0_valid_low_found = 1'h1;
					next_0_valid_low = 3'h7;
					next_0_valid_low_done = 1'h1;
				end
			end
		end
	end
	assign inc_reserve_count = write_alloc & ~write_fill;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			reserve_count <= 16'h0000;
		else if (flush)
			reserve_count <= 16'h0000;
		else if (clk_en) begin
			if (clk_en) begin
				if (inc_reserve_count)
					reserve_count <= reserve_count + 16'h0001;
			end
		end
endmodule
module reservation_fifo_depth_8_w_17_num_per_2 (
	clk,
	clk_en,
	data_in_0,
	data_in_1,
	fill_data_in,
	flush,
	pop,
	push_alloc,
	push_fill,
	push_reserve,
	rst_n,
	data_out_0,
	data_out_1,
	empty,
	full,
	valid
);
	input wire clk;
	input wire clk_en;
	input wire [16:0] data_in_0;
	input wire [16:0] data_in_1;
	input wire [16:0] fill_data_in;
	input wire flush;
	input wire pop;
	input wire push_alloc;
	input wire push_fill;
	input wire push_reserve;
	input wire rst_n;
	output wire [16:0] data_out_0;
	output wire [16:0] data_out_1;
	output wire empty;
	output wire full;
	output reg valid;
	wire clr_item_ptr;
	wire clr_read_ptr;
	wire clr_write_ptr;
	wire [33:0] data_in_packed;
	reg [33:0] data_out;
	wire enable_reserve_ptr;
	wire inc_item_ptr;
	wire inc_read_ptr;
	wire inc_reserve_count;
	wire inc_write_ptr;
	reg item_ptr_addr;
	wire jump_next_0;
	wire [2:0] next_0_valid;
	reg [2:0] next_0_valid_d1;
	reg [2:0] next_0_valid_high;
	reg next_0_valid_high_done;
	reg next_0_valid_high_found;
	reg [2:0] next_0_valid_low;
	reg next_0_valid_low_done;
	reg next_0_valid_low_found;
	reg [3:0] num_items;
	wire read;
	reg [2:0] read_ptr_addr;
	reg [271:0] reg_array;
	reg [15:0] reserve_count;
	wire [2:0] reserve_ptr_val;
	reg [7:0] valid_mask;
	wire write_alloc;
	wire write_fill;
	reg [2:0] write_ptr_addr;
	wire write_reserve;
	wire write_reserve_final;
	assign data_in_packed[0+:17] = data_in_0;
	assign data_in_packed[17+:17] = data_in_1;
	assign data_out_0 = data_out[0+:17];
	assign data_out_1 = data_out[17+:17];
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			item_ptr_addr <= 1'h0;
		else if (flush)
			item_ptr_addr <= 1'h0;
		else if (clk_en) begin
			if (clk_en) begin
				if (clr_item_ptr)
					item_ptr_addr <= 1'h0;
				else if (inc_item_ptr)
					item_ptr_addr <= item_ptr_addr + 1'h1;
			end
		end
	assign inc_item_ptr = push_reserve;
	assign clr_item_ptr = push_reserve & (item_ptr_addr == 1'h1);
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			read_ptr_addr <= 3'h0;
		else if (flush)
			read_ptr_addr <= 3'h0;
		else if (clk_en) begin
			if (clk_en) begin
				if (clr_read_ptr)
					read_ptr_addr <= 3'h0;
				else if (inc_read_ptr)
					read_ptr_addr <= read_ptr_addr + 3'h1;
			end
		end
	assign inc_read_ptr = read;
	assign clr_read_ptr = 1'h0;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			write_ptr_addr <= 3'h0;
		else if (flush)
			write_ptr_addr <= 3'h0;
		else if (clk_en) begin
			if (clk_en) begin
				if (clr_write_ptr)
					write_ptr_addr <= 3'h0;
				else if (inc_write_ptr)
					write_ptr_addr <= write_ptr_addr + 3'h1;
			end
		end
	assign inc_write_ptr = write_alloc | write_fill;
	assign clr_write_ptr = 1'h0;
	assign jump_next_0 = next_0_valid_high_found | next_0_valid_low_found;
	assign enable_reserve_ptr = write_reserve_final | (write_fill & (reserve_ptr_val == write_ptr_addr));
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			next_0_valid_d1 <= 3'h0;
		else if (flush)
			next_0_valid_d1 <= 3'h0;
		else if (clk_en) begin
			if (clk_en) begin
				if (enable_reserve_ptr)
					next_0_valid_d1 <= next_0_valid;
			end
		end
	assign reserve_ptr_val = next_0_valid_d1;
	assign next_0_valid = (write_fill & (((next_0_valid_d1 == write_ptr_addr) | (~next_0_valid_high_found & ~next_0_valid_low_found)) | (next_0_valid_high_found ? next_0_valid_high == write_ptr_addr : next_0_valid_low == write_ptr_addr)) ? write_ptr_addr + 3'h1 : (~next_0_valid_high_found & ~next_0_valid_low_found ? write_ptr_addr : (next_0_valid_high_found ? next_0_valid_high : next_0_valid_low)));
	assign full = num_items == 4'h8;
	assign empty = num_items == 4'h0;
	assign write_fill = (push_fill & push_alloc) & ~full;
	assign write_alloc = push_alloc & ~full;
	assign write_reserve = inc_item_ptr;
	assign write_reserve_final = clr_item_ptr;
	assign read = pop & valid_mask[read_ptr_addr];
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			num_items <= 4'h0;
		else if (flush)
			num_items <= 4'h0;
		else if (clk_en) begin
			if (clk_en) begin
				if (write_alloc & ~read)
					num_items <= num_items + 4'h1;
				else if (~write_alloc & read)
					num_items <= num_items - 4'h1;
			end
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			reg_array <= 272'h0;
		else if (flush)
			reg_array <= 272'h0;
		else if (clk_en) begin
			if (clk_en) begin
				if (write_fill)
					reg_array[(write_ptr_addr * 2) * 17+:17] <= fill_data_in;
				if (write_reserve)
					reg_array[((next_0_valid_d1 * 2) + item_ptr_addr) * 17+:17] <= data_in_packed[item_ptr_addr * 17+:17];
			end
		end
	always @(*) data_out = reg_array[17 * (read_ptr_addr * 2)+:34];
	always @(*) valid = valid_mask[read_ptr_addr];
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			valid_mask <= 8'h00;
		else if (flush)
			valid_mask <= 8'h00;
		else if (clk_en) begin
			if (clk_en) begin
				if (write_fill)
					valid_mask[write_ptr_addr] <= 1'h1;
				if (write_reserve_final)
					valid_mask[next_0_valid_d1] <= 1'h1;
				if (read)
					valid_mask[read_ptr_addr] <= 1'h0;
			end
		end
	always @(*) begin
		next_0_valid_high_found = 1'h0;
		next_0_valid_high = 3'h0;
		next_0_valid_high_done = 1'h0;
		if (~next_0_valid_high_done) begin
			if (next_0_valid_d1 < 3'h0) begin
				if (valid_mask[0] == 1'h0) begin
					next_0_valid_high_found = 1'h1;
					next_0_valid_high = 3'h0;
					next_0_valid_high_done = 1'h1;
				end
			end
		end
		if (~next_0_valid_high_done) begin
			if (next_0_valid_d1 < 3'h1) begin
				if (valid_mask[1] == 1'h0) begin
					next_0_valid_high_found = 1'h1;
					next_0_valid_high = 3'h1;
					next_0_valid_high_done = 1'h1;
				end
			end
		end
		if (~next_0_valid_high_done) begin
			if (next_0_valid_d1 < 3'h2) begin
				if (valid_mask[2] == 1'h0) begin
					next_0_valid_high_found = 1'h1;
					next_0_valid_high = 3'h2;
					next_0_valid_high_done = 1'h1;
				end
			end
		end
		if (~next_0_valid_high_done) begin
			if (next_0_valid_d1 < 3'h3) begin
				if (valid_mask[3] == 1'h0) begin
					next_0_valid_high_found = 1'h1;
					next_0_valid_high = 3'h3;
					next_0_valid_high_done = 1'h1;
				end
			end
		end
		if (~next_0_valid_high_done) begin
			if (next_0_valid_d1 < 3'h4) begin
				if (valid_mask[4] == 1'h0) begin
					next_0_valid_high_found = 1'h1;
					next_0_valid_high = 3'h4;
					next_0_valid_high_done = 1'h1;
				end
			end
		end
		if (~next_0_valid_high_done) begin
			if (next_0_valid_d1 < 3'h5) begin
				if (valid_mask[5] == 1'h0) begin
					next_0_valid_high_found = 1'h1;
					next_0_valid_high = 3'h5;
					next_0_valid_high_done = 1'h1;
				end
			end
		end
		if (~next_0_valid_high_done) begin
			if (next_0_valid_d1 < 3'h6) begin
				if (valid_mask[6] == 1'h0) begin
					next_0_valid_high_found = 1'h1;
					next_0_valid_high = 3'h6;
					next_0_valid_high_done = 1'h1;
				end
			end
		end
		if (~next_0_valid_high_done) begin
			if (next_0_valid_d1 < 3'h7) begin
				if (valid_mask[7] == 1'h0) begin
					next_0_valid_high_found = 1'h1;
					next_0_valid_high = 3'h7;
					next_0_valid_high_done = 1'h1;
				end
			end
		end
	end
	always @(*) begin
		next_0_valid_low_found = 1'h0;
		next_0_valid_low = 3'h0;
		next_0_valid_low_done = 1'h0;
		if (~next_0_valid_low_done) begin
			if (next_0_valid_d1 > 3'h0) begin
				if (valid_mask[0] == 1'h0) begin
					next_0_valid_low_found = 1'h1;
					next_0_valid_low = 3'h0;
					next_0_valid_low_done = 1'h1;
				end
			end
		end
		if (~next_0_valid_low_done) begin
			if (next_0_valid_d1 > 3'h1) begin
				if (valid_mask[1] == 1'h0) begin
					next_0_valid_low_found = 1'h1;
					next_0_valid_low = 3'h1;
					next_0_valid_low_done = 1'h1;
				end
			end
		end
		if (~next_0_valid_low_done) begin
			if (next_0_valid_d1 > 3'h2) begin
				if (valid_mask[2] == 1'h0) begin
					next_0_valid_low_found = 1'h1;
					next_0_valid_low = 3'h2;
					next_0_valid_low_done = 1'h1;
				end
			end
		end
		if (~next_0_valid_low_done) begin
			if (next_0_valid_d1 > 3'h3) begin
				if (valid_mask[3] == 1'h0) begin
					next_0_valid_low_found = 1'h1;
					next_0_valid_low = 3'h3;
					next_0_valid_low_done = 1'h1;
				end
			end
		end
		if (~next_0_valid_low_done) begin
			if (next_0_valid_d1 > 3'h4) begin
				if (valid_mask[4] == 1'h0) begin
					next_0_valid_low_found = 1'h1;
					next_0_valid_low = 3'h4;
					next_0_valid_low_done = 1'h1;
				end
			end
		end
		if (~next_0_valid_low_done) begin
			if (next_0_valid_d1 > 3'h5) begin
				if (valid_mask[5] == 1'h0) begin
					next_0_valid_low_found = 1'h1;
					next_0_valid_low = 3'h5;
					next_0_valid_low_done = 1'h1;
				end
			end
		end
		if (~next_0_valid_low_done) begin
			if (next_0_valid_d1 > 3'h6) begin
				if (valid_mask[6] == 1'h0) begin
					next_0_valid_low_found = 1'h1;
					next_0_valid_low = 3'h6;
					next_0_valid_low_done = 1'h1;
				end
			end
		end
		if (~next_0_valid_low_done) begin
			if (next_0_valid_d1 > 3'h7) begin
				if (valid_mask[7] == 1'h0) begin
					next_0_valid_low_found = 1'h1;
					next_0_valid_low = 3'h7;
					next_0_valid_low_done = 1'h1;
				end
			end
		end
	end
	assign inc_reserve_count = write_alloc & ~write_fill;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			reserve_count <= 16'h0000;
		else if (flush)
			reserve_count <= 16'h0000;
		else if (clk_en) begin
			if (clk_en) begin
				if (inc_reserve_count)
					reserve_count <= reserve_count + 16'h0001;
			end
		end
endmodule
module scanner_pipe (
	ID_out_ready,
	addr_out_ready,
	block_mode,
	block_rd_out_ready,
	clk,
	clk_en,
	coord_out_ready,
	dense,
	dim_size,
	do_repeat,
	flush,
	inner_dim_offset,
	lookup,
	op_out_ready,
	pos_out_ready,
	rd_rsp_data_in,
	rd_rsp_data_in_valid,
	repeat_factor,
	repeat_outer_inner_n,
	root,
	rst_n,
	spacc_mode,
	stop_lvl,
	tile_en,
	us_pos_in,
	us_pos_in_valid,
	ID_out,
	ID_out_valid,
	addr_out,
	addr_out_valid,
	block_rd_out,
	block_rd_out_valid,
	coord_out,
	coord_out_valid,
	op_out,
	op_out_valid,
	pos_out,
	pos_out_valid,
	rd_rsp_data_in_ready,
	us_pos_in_ready
);
	input wire ID_out_ready;
	input wire addr_out_ready;
	input wire block_mode;
	input wire block_rd_out_ready;
	input wire clk;
	input wire clk_en;
	input wire coord_out_ready;
	input wire dense;
	input wire [15:0] dim_size;
	input wire do_repeat;
	input wire flush;
	input wire [15:0] inner_dim_offset;
	input wire lookup;
	input wire op_out_ready;
	input wire pos_out_ready;
	input wire [16:0] rd_rsp_data_in;
	input wire rd_rsp_data_in_valid;
	input wire [15:0] repeat_factor;
	input wire repeat_outer_inner_n;
	input wire root;
	input wire rst_n;
	input wire spacc_mode;
	input wire [15:0] stop_lvl;
	input wire tile_en;
	input wire [16:0] us_pos_in;
	input wire us_pos_in_valid;
	output wire [16:0] ID_out;
	output wire ID_out_valid;
	output wire [16:0] addr_out;
	output wire addr_out_valid;
	output wire [16:0] block_rd_out;
	output wire block_rd_out_valid;
	output wire [16:0] coord_out;
	output wire coord_out_valid;
	output wire [16:0] op_out;
	output wire op_out_valid;
	output wire [16:0] pos_out;
	output wire pos_out_valid;
	output wire rd_rsp_data_in_ready;
	output wire us_pos_in_ready;
	wire [16:0] ID_out_fifo_data_in;
	wire ID_out_fifo_empty;
	wire ID_out_fifo_full;
	wire ID_out_fifo_push;
	wire [15:0] ID_out_to_fifo;
	reg [15:0] READS_MADE;
	reg [15:0] READS_REC_CRD_READ;
	wire [16:0] addr_out_fifo_data_in;
	wire addr_out_fifo_empty;
	wire addr_out_fifo_full;
	wire addr_out_fifo_push;
	wire [15:0] addr_out_to_fifo;
	wire [1:0] base_rr;
	wire block_rd_fifo_empty;
	wire block_rd_fifo_full;
	wire block_rd_fifo_push;
	wire clr_fiber_addr;
	wire clr_final_pushed_done;
	wire clr_pop_infifo_sticky;
	reg clr_pushed_done_crd;
	reg clr_pushed_done_seg;
	reg clr_readout_loop_crd;
	reg clr_readout_loop_seg;
	wire clr_rep;
	reg clr_req_made_crd;
	reg clr_req_made_seg;
	reg clr_req_rec_crd;
	reg clr_req_rec_seg;
	wire clr_seen_root_eos;
	wire clr_used_data;
	wire [16:0] coord_fifo_in_packed;
	wire [16:0] coord_fifo_out_packed;
	wire coordinate_fifo_empty;
	wire coordinate_fifo_full;
	wire coordinate_fifo_push;
	reg [15:0] crd_ID_out_to_fifo;
	reg [15:0] crd_addr_out_to_fifo;
	wire crd_grant_push;
	reg crd_in_done_state;
	reg [15:0] crd_op_out_to_fifo;
	reg [16:0] crd_out_to_fifo;
	reg crd_pop_infifo;
	reg crd_rd_rsp_fifo_pop;
	reg crd_req_push;
	wire [16:0] crd_res_fifo_data_in_0;
	wire [16:0] crd_res_fifo_data_out;
	wire [16:0] crd_res_fifo_fill_data_in;
	wire crd_res_fifo_full;
	wire crd_res_fifo_pop;
	reg crd_res_fifo_push_alloc;
	wire crd_res_fifo_push_alloc_0;
	reg crd_res_fifo_push_fill;
	wire crd_res_fifo_push_fill_0;
	wire crd_res_fifo_push_reserve_0;
	wire crd_res_fifo_valid;
	wire crd_stop_lvl_geq;
	wire done_in;
	reg en_reg_data_in;
	wire eos_in;
	wire [15:0] fiber_addr;
	reg [15:0] fiber_addr_pre;
	reg [15:0] fiber_addr_pre_d1;
	reg [15:0] fiber_addr_pre_d1_d1;
	wire fifo_full;
	wire [1:0] fifo_full_pre;
	wire [16:0] fifo_out_us_packed;
	wire fifo_us_full;
	wire [16:0] fifo_us_in_packed;
	wire final_pushed_done_sticky_sticky;
	reg final_pushed_done_sticky_was_high;
	wire gclk;
	wire go_to_readout_sticky_sticky;
	reg go_to_readout_sticky_was_high;
	wire inc_fiber_addr;
	wire inc_rep;
	reg inc_req_made_crd;
	reg inc_req_made_seg;
	reg inc_req_rec_crd;
	reg inc_req_rec_seg;
	wire inc_requests_REC_CRD_READ;
	wire inc_requests_made_CRDDD_READ;
	wire infifo_eos_in;
	wire [15:0] infifo_pos_in;
	wire infifo_valid_in;
	wire [16:0] input_fifo_data_out;
	wire input_fifo_empty;
	wire iter_finish_sticky;
	reg iter_finish_was_high;
	wire last_stop_done;
	reg [16:0] last_stop_token;
	wire last_valid_accepting;
	wire maybe_in;
	wire [15:0] next_seq_addr;
	wire [15:0] next_seq_length;
	wire no_outfifo_full;
	reg [15:0] num_reps;
	reg [15:0] num_req_made_crd;
	reg [15:0] num_req_made_seg;
	reg [15:0] num_req_rec_crd;
	reg [15:0] num_req_rec_seg;
	wire [16:0] op_out_fifo_data_in;
	wire op_out_fifo_empty;
	wire op_out_fifo_full;
	wire op_out_fifo_push;
	wire [15:0] op_out_to_fifo;
	reg [15:0] payload_ptr;
	wire pop_infifo;
	wire pop_infifo_sticky_sticky;
	reg pop_infifo_sticky_was_high;
	wire [15:0] pos_addr;
	wire pos_fifo_empty;
	wire pos_fifo_full;
	wire [16:0] pos_fifo_in_packed;
	wire [16:0] pos_fifo_out_packed;
	reg pos_out_fifo_push;
	reg [16:0] pos_out_to_fifo;
	wire [15:0] ptr_in;
	reg [15:0] ptr_in_d1;
	reg ptr_reg_en;
	wire pushed_done_sticky_sticky;
	reg pushed_done_sticky_was_high;
	wire rd_rsp_fifo_empty;
	wire rd_rsp_fifo_full;
	wire [16:0] rd_rsp_fifo_out_data;
	reg [16:0] rd_rsp_fifo_out_data_d1;
	wire rd_rsp_fifo_valid;
	wire readout_dst_crd;
	wire readout_dst_seg;
	wire readout_loop_sticky_sticky;
	reg readout_loop_sticky_was_high;
	wire rep_finish_sticky;
	reg rep_finish_was_high;
	wire [1:0] rr_arbiter_grant_out;
	reg [3:0] scan_seq_crd_current_state;
	reg [3:0] scan_seq_crd_next_state;
	reg [3:0] scan_seq_seg_current_state;
	reg [3:0] scan_seq_seg_next_state;
	wire seen_root_eos_sticky;
	reg seen_root_eos_was_high;
	reg [15:0] seg_ID_out_to_fifo;
	reg [15:0] seg_addr_out_to_fifo;
	wire seg_grant_push;
	reg seg_in_done_state;
	reg seg_in_start_state;
	reg [15:0] seg_op_out_to_fifo;
	reg seg_pop_infifo;
	reg seg_rd_rsp_fifo_pop;
	reg seg_req_push;
	wire [16:0] seg_res_fifo_data_out_0;
	wire [16:0] seg_res_fifo_data_out_1;
	wire seg_res_fifo_done_out;
	reg [16:0] seg_res_fifo_fill_data_in;
	wire seg_res_fifo_full;
	reg seg_res_fifo_pop;
	wire seg_res_fifo_pop_0;
	reg seg_res_fifo_push_alloc;
	wire seg_res_fifo_push_alloc_0;
	reg seg_res_fifo_push_fill;
	wire seg_res_fifo_push_fill_0;
	wire seg_res_fifo_push_reserve_0;
	wire seg_res_fifo_valid;
	wire seg_stop_lvl_geq;
	wire seg_stop_lvl_geq_p1;
	reg [15:0] seq_addr;
	reg [15:0] seq_length;
	wire [15:0] seq_length_ptr_math;
	wire set_final_pushed_done;
	reg set_pushed_done_crd;
	reg set_pushed_done_seg;
	reg set_readout_loop_crd;
	reg set_readout_loop_seg;
	wire update_seq_state;
	reg [15:0] us_fifo_inject_data;
	reg us_fifo_inject_eos;
	reg us_fifo_inject_push;
	wire us_fifo_push;
	wire use_data_sticky_sticky;
	reg use_data_sticky_was_high;
	reg [15:0] valid_cnt;
	wire valid_inc;
	wire valid_rst;
	assign gclk = clk & tile_en;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			fiber_addr_pre <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				fiber_addr_pre <= 16'h0000;
			else if (clr_fiber_addr)
				fiber_addr_pre <= 16'h0000;
			else if (inc_fiber_addr)
				fiber_addr_pre <= fiber_addr_pre + 16'h0001;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			num_reps <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				num_reps <= 16'h0000;
			else if (clr_rep)
				num_reps <= 16'h0000;
			else if (inc_rep)
				num_reps <= num_reps + 16'h0001;
		end
	assign us_fifo_push = (root ? us_fifo_inject_push : us_pos_in_valid);
	assign fifo_us_in_packed[16] = (root ? us_fifo_inject_eos : us_pos_in[16]);
	assign fifo_us_in_packed[15:0] = (root ? us_fifo_inject_data : us_pos_in[15:0]);
	assign infifo_eos_in = fifo_out_us_packed[16];
	assign infifo_pos_in = fifo_out_us_packed[15:0];
	assign pop_infifo = seg_pop_infifo | crd_pop_infifo;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			pop_infifo_sticky_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				pop_infifo_sticky_was_high <= 1'h0;
			else if (clr_pop_infifo_sticky)
				pop_infifo_sticky_was_high <= 1'h0;
			else if (pop_infifo)
				pop_infifo_sticky_was_high <= 1'h1;
		end
	assign pop_infifo_sticky_sticky = pop_infifo_sticky_was_high;
	assign fifo_out_us_packed = input_fifo_data_out;
	assign us_pos_in_ready = ~fifo_us_full;
	assign infifo_valid_in = ~input_fifo_empty;
	assign rd_rsp_data_in_ready = ~rd_rsp_fifo_full;
	assign rd_rsp_fifo_valid = ~rd_rsp_fifo_empty;
	assign base_rr = {crd_req_push, seg_req_push};
	assign {crd_grant_push, seg_grant_push} = rr_arbiter_grant_out;
	assign addr_out_to_fifo = (crd_grant_push ? crd_addr_out_to_fifo : seg_addr_out_to_fifo);
	assign op_out_to_fifo = (crd_grant_push ? crd_op_out_to_fifo : seg_op_out_to_fifo);
	assign ID_out_to_fifo = (crd_grant_push ? crd_ID_out_to_fifo : seg_ID_out_to_fifo);
	assign addr_out_fifo_push = seg_grant_push | crd_grant_push;
	assign addr_out_fifo_data_in = {1'h0, addr_out_to_fifo};
	assign addr_out_valid = ~addr_out_fifo_empty;
	assign op_out_fifo_push = seg_grant_push | crd_grant_push;
	assign op_out_fifo_data_in = {1'h0, op_out_to_fifo};
	assign op_out_valid = ~op_out_fifo_empty;
	assign ID_out_fifo_push = seg_grant_push | crd_grant_push;
	assign ID_out_fifo_data_in = {1'h0, ID_out_to_fifo};
	assign ID_out_valid = ~ID_out_fifo_empty;
	assign no_outfifo_full = ~((ID_out_fifo_full | op_out_fifo_full) | addr_out_fifo_full);
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			pushed_done_sticky_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				pushed_done_sticky_was_high <= 1'h0;
			else if (clr_pushed_done_seg | clr_pushed_done_crd)
				pushed_done_sticky_was_high <= 1'h0;
			else if (set_pushed_done_seg | set_pushed_done_crd)
				pushed_done_sticky_was_high <= 1'h1;
		end
	assign pushed_done_sticky_sticky = pushed_done_sticky_was_high;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			readout_loop_sticky_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				readout_loop_sticky_was_high <= 1'h0;
			else if (clr_readout_loop_seg | clr_readout_loop_crd)
				readout_loop_sticky_was_high <= 1'h0;
			else if (set_readout_loop_seg | set_readout_loop_crd)
				readout_loop_sticky_was_high <= 1'h1;
		end
	assign readout_loop_sticky_sticky = readout_loop_sticky_was_high;
	assign seg_res_fifo_push_alloc_0 = seg_res_fifo_push_alloc & ~lookup;
	assign seg_res_fifo_push_reserve_0 = ((rd_rsp_fifo_valid & (rd_rsp_fifo_out_data[16] == 1'h0)) & ~block_mode) & ~lookup;
	assign seg_res_fifo_push_fill_0 = seg_res_fifo_push_fill & ~lookup;
	assign seg_res_fifo_pop_0 = seg_res_fifo_pop & ~lookup;
	assign crd_res_fifo_data_in_0 = {1'h0, rd_rsp_fifo_out_data[15:0]};
	assign crd_res_fifo_fill_data_in = (lookup ? seg_res_fifo_fill_data_in : (dense ? crd_out_to_fifo : seg_res_fifo_data_out_0));
	assign crd_res_fifo_push_alloc_0 = (lookup ? seg_res_fifo_push_alloc : crd_res_fifo_push_alloc);
	assign crd_res_fifo_push_reserve_0 = rd_rsp_fifo_valid & (((rd_rsp_fifo_out_data[16] == 1'h1) | block_mode) | lookup);
	assign crd_res_fifo_push_fill_0 = (lookup ? seg_res_fifo_push_fill : crd_res_fifo_push_fill);
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			last_stop_token <= 17'h00000;
		else if (clk_en) begin
			if (flush)
				last_stop_token <= 17'h00000;
			else if ((seg_in_start_state ? 1'h0 : (((seg_res_fifo_push_fill & seg_res_fifo_push_alloc) & (lookup ? ~crd_res_fifo_full : ~seg_res_fifo_full)) & seg_res_fifo_fill_data_in[16]) & (seg_res_fifo_fill_data_in[9:8] == 2'h0)))
				last_stop_token <= (seg_in_start_state ? input_fifo_data_out + 17'h00001 : seg_res_fifo_fill_data_in);
		end
	assign last_stop_done = last_stop_token[15:0] == (stop_lvl + 16'h0002);
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			use_data_sticky_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				use_data_sticky_was_high <= 1'h0;
			else if (clr_used_data)
				use_data_sticky_was_high <= 1'h0;
			else if (infifo_valid_in & ~infifo_eos_in)
				use_data_sticky_was_high <= 1'h1;
		end
	assign use_data_sticky_sticky = use_data_sticky_was_high;
	assign clr_used_data = readout_loop_sticky_sticky & spacc_mode;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			valid_cnt <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				valid_cnt <= 16'h0000;
			else if (valid_rst)
				valid_cnt <= 16'h0000;
			else if (valid_inc)
				valid_cnt <= valid_cnt + 16'h0001;
		end
	assign ptr_in = rd_rsp_fifo_out_data[15:0];
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			ptr_in_d1 <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				ptr_in_d1 <= 16'h0000;
			else if (ptr_reg_en)
				ptr_in_d1 <= ptr_in;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			fiber_addr_pre_d1 <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				fiber_addr_pre_d1 <= 16'h0000;
			else
				fiber_addr_pre_d1 <= fiber_addr_pre;
		end
	assign seq_length_ptr_math = seg_res_fifo_data_out_1 - seg_res_fifo_data_out_0[15:0];
	assign pos_addr = (root ? 16'h0000 : infifo_pos_in);
	assign next_seq_addr = ptr_in_d1 + inner_dim_offset;
	always @(posedge clk or negedge rst_n)
		if (~rst_n) begin
			seq_length <= 16'h0000;
			seq_addr <= 16'h0000;
			payload_ptr <= 16'h0000;
		end
		else if (clk_en) begin
			if (flush) begin
				seq_length <= 16'h0000;
				seq_addr <= 16'h0000;
				payload_ptr <= 16'h0000;
			end
			else if (update_seq_state) begin
				seq_length <= next_seq_length;
				seq_addr <= next_seq_addr;
				payload_ptr <= ptr_in_d1;
			end
		end
	assign fiber_addr = fiber_addr_pre + seq_addr;
	assign fifo_full = |fifo_full_pre;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			iter_finish_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				iter_finish_was_high <= 1'h0;
			else if (clr_fiber_addr)
				iter_finish_was_high <= 1'h0;
			else if (last_valid_accepting)
				iter_finish_was_high <= 1'h1;
		end
	assign iter_finish_sticky = last_valid_accepting | iter_finish_was_high;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			rep_finish_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				rep_finish_was_high <= 1'h0;
			else if (clr_rep)
				rep_finish_was_high <= 1'h0;
			else if (((repeat_factor - 16'h0001) == num_reps) & inc_rep)
				rep_finish_was_high <= 1'h1;
		end
	assign rep_finish_sticky = (((repeat_factor - 16'h0001) == num_reps) & inc_rep) | rep_finish_was_high;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			seen_root_eos_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				seen_root_eos_was_high <= 1'h0;
			else if (clr_seen_root_eos)
				seen_root_eos_was_high <= 1'h0;
			else if (infifo_eos_in & (infifo_pos_in == 16'h0000))
				seen_root_eos_was_high <= 1'h1;
		end
	assign seen_root_eos_sticky = (infifo_eos_in & (infifo_pos_in == 16'h0000)) | seen_root_eos_was_high;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			rd_rsp_fifo_out_data_d1 <= 17'h00000;
		else if (clk_en) begin
			if (flush)
				rd_rsp_fifo_out_data_d1 <= 17'h00000;
			else if (en_reg_data_in)
				rd_rsp_fifo_out_data_d1 <= rd_rsp_fifo_out_data;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			fiber_addr_pre_d1_d1 <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				fiber_addr_pre_d1_d1 <= 16'h0000;
			else if (en_reg_data_in)
				fiber_addr_pre_d1_d1 <= fiber_addr_pre_d1;
		end
	assign done_in = (infifo_eos_in & infifo_valid_in) & (infifo_pos_in[9:8] == 2'h1);
	assign eos_in = (infifo_eos_in & infifo_valid_in) & (infifo_pos_in[9:8] == 2'h0);
	assign maybe_in = (infifo_eos_in & infifo_valid_in) & (infifo_pos_in[9:8] == 2'h2);
	assign seg_stop_lvl_geq = (seg_res_fifo_fill_data_in[16] & (seg_res_fifo_fill_data_in[9:8] == 2'h0)) & (seg_res_fifo_fill_data_in[7:0] >= stop_lvl[7:0]);
	assign seg_stop_lvl_geq_p1 = (seg_res_fifo_fill_data_in[16] & (seg_res_fifo_fill_data_in[9:8] == 2'h0)) & (seg_res_fifo_fill_data_in[7:0] >= (stop_lvl[7:0] + 8'h01));
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			go_to_readout_sticky_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				go_to_readout_sticky_was_high <= 1'h0;
			else if (clr_readout_loop_seg)
				go_to_readout_sticky_was_high <= 1'h0;
			else if ((seg_stop_lvl_geq_p1 & seg_res_fifo_push_alloc) & seg_res_fifo_push_fill)
				go_to_readout_sticky_was_high <= 1'h1;
		end
	assign go_to_readout_sticky_sticky = ((seg_stop_lvl_geq_p1 & seg_res_fifo_push_alloc) & seg_res_fifo_push_fill) | go_to_readout_sticky_was_high;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			num_req_made_seg <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				num_req_made_seg <= 16'h0000;
			else if (clr_req_made_seg)
				num_req_made_seg <= 16'h0000;
			else if (inc_req_made_seg)
				num_req_made_seg <= num_req_made_seg + 16'h0001;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			num_req_rec_seg <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				num_req_rec_seg <= 16'h0000;
			else if (clr_req_rec_seg)
				num_req_rec_seg <= 16'h0000;
			else if (inc_req_rec_seg)
				num_req_rec_seg <= num_req_rec_seg + 16'h0001;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			num_req_made_crd <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				num_req_made_crd <= 16'h0000;
			else if (clr_req_made_crd)
				num_req_made_crd <= 16'h0000;
			else if (inc_req_made_crd)
				num_req_made_crd <= num_req_made_crd + 16'h0001;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			num_req_rec_crd <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				num_req_rec_crd <= 16'h0000;
			else if (clr_req_rec_crd)
				num_req_rec_crd <= 16'h0000;
			else if (inc_req_rec_crd)
				num_req_rec_crd <= num_req_rec_crd + 16'h0001;
		end
	assign seg_res_fifo_done_out = (seg_res_fifo_valid & seg_res_fifo_data_out_0[16]) & (seg_res_fifo_data_out_0[9:8] == 2'h1);
	assign crd_stop_lvl_geq = ((seg_res_fifo_valid & seg_res_fifo_data_out_0[16]) & (seg_res_fifo_data_out_0[9:8] == 2'h0)) & (seg_res_fifo_data_out_0[7:0] >= stop_lvl[7:0]);
	assign readout_dst_crd = readout_loop_sticky_sticky;
	assign readout_dst_seg = readout_loop_sticky_sticky;
	assign inc_requests_made_CRDDD_READ = crd_grant_push;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			READS_MADE <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				READS_MADE <= 16'h0000;
			else if (inc_requests_made_CRDDD_READ)
				READS_MADE <= READS_MADE + 16'h0001;
		end
	assign inc_requests_REC_CRD_READ = rd_rsp_fifo_valid & (rd_rsp_fifo_out_data[16] == 1'h1);
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			READS_REC_CRD_READ <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				READS_REC_CRD_READ <= 16'h0000;
			else if (inc_requests_REC_CRD_READ)
				READS_REC_CRD_READ <= READS_REC_CRD_READ + 16'h0001;
		end
	assign coord_fifo_in_packed = crd_res_fifo_data_out;
	assign coord_out[16] = coord_fifo_out_packed[16];
	assign coord_out[15:0] = coord_fifo_out_packed[15:0];
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			final_pushed_done_sticky_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				final_pushed_done_sticky_was_high <= 1'h0;
			else if (clr_final_pushed_done)
				final_pushed_done_sticky_was_high <= 1'h0;
			else if (set_final_pushed_done)
				final_pushed_done_sticky_was_high <= 1'h1;
		end
	assign final_pushed_done_sticky_sticky = final_pushed_done_sticky_was_high;
	assign set_final_pushed_done = (((((crd_res_fifo_valid & ~block_mode) & crd_res_fifo_data_out[16]) & crd_res_fifo_valid) & (crd_res_fifo_data_out[9:8] == 2'h3)) & spacc_mode) & crd_res_fifo_data_out[0];
	assign clr_final_pushed_done = (((((crd_res_fifo_valid & ~block_mode) & crd_res_fifo_data_out[16]) & crd_res_fifo_valid) & (crd_res_fifo_data_out[9:8] == 2'h3)) & spacc_mode) & ~crd_res_fifo_data_out[0];
	assign coordinate_fifo_push = ((crd_res_fifo_valid & ~block_mode) & ~(spacc_mode & final_pushed_done_sticky_sticky)) & ~((crd_res_fifo_data_out[16] & crd_res_fifo_valid) & (crd_res_fifo_data_out[9:8] == 2'h3));
	assign coord_out_valid = ~coordinate_fifo_empty;
	assign fifo_full_pre[0] = coordinate_fifo_full;
	assign crd_res_fifo_pop = (block_mode ? ~block_rd_fifo_full : (spacc_mode ? ((crd_res_fifo_data_out[16] & crd_res_fifo_valid) & (crd_res_fifo_data_out[9:8] == 2'h3) ? 1'h1 : (final_pushed_done_sticky_sticky ? ~block_rd_fifo_full : ~coordinate_fifo_full)) : ~coordinate_fifo_full));
	assign pos_fifo_in_packed = pos_out_to_fifo;
	assign pos_out[16] = pos_fifo_out_packed[16];
	assign pos_out[15:0] = pos_fifo_out_packed[15:0];
	assign pos_out_valid = ~pos_fifo_empty;
	assign fifo_full_pre[1] = pos_fifo_full;
	assign block_rd_fifo_push = (crd_res_fifo_valid & (block_mode | (spacc_mode & final_pushed_done_sticky_sticky))) & ~((crd_res_fifo_data_out[16] & crd_res_fifo_valid) & (crd_res_fifo_data_out[9:8] == 2'h3));
	assign block_rd_out_valid = ~block_rd_fifo_empty;
	always @(posedge clk or negedge rst_n)
		if (!rst_n)
			scan_seq_crd_current_state <= 4'hd;
		else if (clk_en) begin
			if (flush)
				scan_seq_crd_current_state <= 4'hd;
			else
				scan_seq_crd_current_state <= scan_seq_crd_next_state;
		end
	always @(*) begin
		scan_seq_crd_next_state = scan_seq_crd_current_state;
		case (scan_seq_crd_current_state)
			4'h0:
				if ((num_req_rec_crd == ptr_in_d1) & ~lookup)
					scan_seq_crd_next_state = 4'h5;
				else if ((num_req_rec_crd == ptr_in_d1) & lookup)
					scan_seq_crd_next_state = 4'h8;
				else
					scan_seq_crd_next_state = 4'h0;
			4'h1:
				if (rd_rsp_fifo_valid)
					scan_seq_crd_next_state = 4'h0;
				else
					scan_seq_crd_next_state = 4'h1;
			4'h2:
				if (crd_grant_push)
					scan_seq_crd_next_state = 4'h1;
				else
					scan_seq_crd_next_state = 4'h2;
			4'h3:
				if (num_req_rec_crd == ptr_in_d1)
					scan_seq_crd_next_state = 4'h8;
				else
					scan_seq_crd_next_state = 4'h3;
			4'h4:
				if (rd_rsp_fifo_valid)
					scan_seq_crd_next_state = 4'h3;
				else
					scan_seq_crd_next_state = 4'h4;
			4'h5:
				if (crd_grant_push)
					scan_seq_crd_next_state = 4'h4;
				else
					scan_seq_crd_next_state = 4'h5;
			4'h6: scan_seq_crd_next_state = 4'h6;
			4'h7:
				if (~spacc_mode | (spacc_mode & seg_in_done_state))
					scan_seq_crd_next_state = 4'hd;
			4'h8:
				if ((crd_grant_push & block_mode) & ~lookup)
					scan_seq_crd_next_state = 4'h9;
				else if ((crd_grant_push & pushed_done_sticky_sticky) & spacc_mode)
					scan_seq_crd_next_state = 4'ha;
				else if (crd_grant_push & (~spacc_mode | ~pushed_done_sticky_sticky))
					scan_seq_crd_next_state = 4'h7;
				else
					scan_seq_crd_next_state = 4'h8;
			4'h9:
				if (crd_grant_push)
					scan_seq_crd_next_state = 4'h7;
				else
					scan_seq_crd_next_state = 4'h9;
			4'ha:
				if (~crd_res_fifo_full & ~pos_fifo_full)
					scan_seq_crd_next_state = 4'h7;
			4'hb: scan_seq_crd_next_state = 4'h7;
			4'hc:
				if (((seg_res_fifo_done_out | (spacc_mode & crd_stop_lvl_geq)) & ~crd_res_fifo_full) & ~pos_fifo_full)
					scan_seq_crd_next_state = 4'h8;
			4'hd:
				if (block_mode & tile_en)
					scan_seq_crd_next_state = 4'h2;
				else if ((dense & ~lookup) & tile_en)
					scan_seq_crd_next_state = 4'h6;
				else if ((~dense & ~lookup) & tile_en)
					scan_seq_crd_next_state = 4'hc;
			default: scan_seq_crd_next_state = scan_seq_crd_current_state;
		endcase
	end
	function automatic [16:0] sv2v_cast_17;
		input reg [16:0] inp;
		sv2v_cast_17 = inp;
	endfunction
	always @(*)
		case (scan_seq_crd_current_state)
			4'h0: begin : scan_seq_crd_BLOCK_1_RD_Output
				crd_addr_out_to_fifo = num_req_made_crd;
				crd_op_out_to_fifo = 16'h0001;
				crd_ID_out_to_fifo = 16'h0000;
				crd_req_push = (num_req_made_crd < ptr_in_d1) & ~crd_res_fifo_full;
				crd_rd_rsp_fifo_pop = num_req_rec_crd < ptr_in_d1;
				pos_out_fifo_push = 1'h0;
				crd_pop_infifo = 1'h0;
				en_reg_data_in = 1'h0;
				pos_out_to_fifo = 17'h00000;
				crd_out_to_fifo = 17'h00000;
				inc_req_made_crd = ((num_req_made_crd < ptr_in_d1) & crd_grant_push) & ~crd_res_fifo_full;
				clr_req_made_crd = 1'h0;
				inc_req_rec_crd = (num_req_rec_crd < ptr_in_d1) & rd_rsp_fifo_valid;
				clr_req_rec_crd = 1'h0;
				crd_res_fifo_push_alloc = ((num_req_made_crd < ptr_in_d1) & crd_grant_push) & ~crd_res_fifo_full;
				crd_res_fifo_push_fill = 1'h0;
				ptr_reg_en = 1'h0;
				seg_res_fifo_pop = 1'h0;
				clr_readout_loop_crd = 1'h0;
				set_readout_loop_crd = 1'h0;
				clr_pushed_done_crd = 1'h0;
				crd_in_done_state = 1'h0;
				set_pushed_done_crd = 1'h0;
			end
			4'h1: begin : scan_seq_crd_BLOCK_1_SIZE_REC_Output
				crd_addr_out_to_fifo = 16'h0000;
				crd_op_out_to_fifo = 16'h0000;
				crd_ID_out_to_fifo = 16'h0000;
				crd_req_push = 1'h0;
				crd_rd_rsp_fifo_pop = 1'h1;
				pos_out_fifo_push = 1'h0;
				crd_pop_infifo = 1'h0;
				en_reg_data_in = 1'h0;
				pos_out_to_fifo = 17'h00000;
				crd_out_to_fifo = 17'h00000;
				inc_req_made_crd = 1'h0;
				clr_req_made_crd = 1'h1;
				inc_req_rec_crd = 1'h0;
				clr_req_rec_crd = 1'h0;
				crd_res_fifo_push_alloc = 1'h0;
				crd_res_fifo_push_fill = 1'h0;
				ptr_reg_en = rd_rsp_fifo_valid;
				seg_res_fifo_pop = 1'h0;
				clr_readout_loop_crd = 1'h0;
				set_readout_loop_crd = 1'h0;
				clr_pushed_done_crd = 1'h0;
				crd_in_done_state = 1'h0;
				set_pushed_done_crd = 1'h0;
			end
			4'h2: begin : scan_seq_crd_BLOCK_1_SIZE_REQ_Output
				crd_addr_out_to_fifo = 16'h0000;
				crd_op_out_to_fifo = 16'h0002;
				crd_ID_out_to_fifo = 16'h0000;
				crd_req_push = ~crd_res_fifo_full;
				crd_rd_rsp_fifo_pop = 1'h0;
				pos_out_fifo_push = 1'h0;
				crd_pop_infifo = 1'h0;
				en_reg_data_in = 1'h0;
				pos_out_to_fifo = 17'h00000;
				crd_out_to_fifo = 17'h00000;
				inc_req_made_crd = 1'h0;
				clr_req_made_crd = 1'h0;
				inc_req_rec_crd = 1'h0;
				clr_req_rec_crd = 1'h0;
				crd_res_fifo_push_alloc = ~crd_res_fifo_full & crd_grant_push;
				crd_res_fifo_push_fill = 1'h0;
				ptr_reg_en = 1'h0;
				seg_res_fifo_pop = 1'h0;
				clr_readout_loop_crd = 1'h0;
				set_readout_loop_crd = 1'h0;
				clr_pushed_done_crd = 1'h0;
				crd_in_done_state = 1'h0;
				set_pushed_done_crd = 1'h0;
			end
			4'h3: begin : scan_seq_crd_BLOCK_2_RD_Output
				crd_addr_out_to_fifo = num_req_made_crd;
				crd_op_out_to_fifo = 16'h0001;
				crd_ID_out_to_fifo = 16'h0001;
				crd_req_push = (num_req_made_crd < ptr_in_d1) & ~crd_res_fifo_full;
				crd_rd_rsp_fifo_pop = num_req_rec_crd < ptr_in_d1;
				pos_out_fifo_push = 1'h0;
				crd_pop_infifo = 1'h0;
				en_reg_data_in = 1'h0;
				pos_out_to_fifo = 17'h00000;
				crd_out_to_fifo = 17'h00000;
				inc_req_made_crd = ((num_req_made_crd < ptr_in_d1) & crd_grant_push) & ~crd_res_fifo_full;
				clr_req_made_crd = 1'h0;
				inc_req_rec_crd = (num_req_rec_crd < ptr_in_d1) & rd_rsp_fifo_valid;
				clr_req_rec_crd = 1'h0;
				crd_res_fifo_push_alloc = ((num_req_made_crd < ptr_in_d1) & crd_grant_push) & ~crd_res_fifo_full;
				crd_res_fifo_push_fill = 1'h0;
				ptr_reg_en = 1'h0;
				seg_res_fifo_pop = 1'h0;
				clr_readout_loop_crd = 1'h0;
				set_readout_loop_crd = 1'h0;
				clr_pushed_done_crd = 1'h0;
				crd_in_done_state = 1'h0;
				set_pushed_done_crd = 1'h0;
			end
			4'h4: begin : scan_seq_crd_BLOCK_2_SIZE_REC_Output
				crd_addr_out_to_fifo = 16'h0000;
				crd_op_out_to_fifo = 16'h0000;
				crd_ID_out_to_fifo = 16'h0000;
				crd_req_push = 1'h0;
				crd_rd_rsp_fifo_pop = 1'h1;
				pos_out_fifo_push = 1'h0;
				crd_pop_infifo = 1'h0;
				en_reg_data_in = 1'h0;
				pos_out_to_fifo = 17'h00000;
				crd_out_to_fifo = 17'h00000;
				inc_req_made_crd = 1'h0;
				clr_req_made_crd = 1'h1;
				inc_req_rec_crd = 1'h0;
				clr_req_rec_crd = 1'h1;
				crd_res_fifo_push_alloc = 1'h0;
				crd_res_fifo_push_fill = 1'h0;
				ptr_reg_en = rd_rsp_fifo_valid;
				seg_res_fifo_pop = 1'h0;
				clr_readout_loop_crd = 1'h0;
				set_readout_loop_crd = 1'h0;
				clr_pushed_done_crd = 1'h0;
				crd_in_done_state = 1'h0;
				set_pushed_done_crd = 1'h0;
			end
			4'h5: begin : scan_seq_crd_BLOCK_2_SIZE_REQ_Output
				crd_addr_out_to_fifo = 16'h0000;
				crd_op_out_to_fifo = 16'h0002;
				crd_ID_out_to_fifo = 16'h0001;
				crd_req_push = ~crd_res_fifo_full;
				crd_rd_rsp_fifo_pop = 1'h0;
				pos_out_fifo_push = 1'h0;
				crd_pop_infifo = 1'h0;
				en_reg_data_in = 1'h0;
				pos_out_to_fifo = 17'h00000;
				crd_out_to_fifo = 17'h00000;
				inc_req_made_crd = 1'h0;
				clr_req_made_crd = 1'h0;
				inc_req_rec_crd = 1'h0;
				clr_req_rec_crd = 1'h0;
				crd_res_fifo_push_alloc = ~crd_res_fifo_full & crd_grant_push;
				crd_res_fifo_push_fill = 1'h0;
				ptr_reg_en = 1'h0;
				seg_res_fifo_pop = 1'h0;
				clr_readout_loop_crd = 1'h0;
				set_readout_loop_crd = 1'h0;
				clr_pushed_done_crd = 1'h0;
				crd_in_done_state = 1'h0;
				set_pushed_done_crd = 1'h0;
			end
			4'h6: begin : scan_seq_crd_DENSE_STRM_Output
				crd_addr_out_to_fifo = 16'h0000;
				crd_op_out_to_fifo = 16'h0000;
				crd_ID_out_to_fifo = 16'h0000;
				crd_req_push = 1'h0;
				crd_rd_rsp_fifo_pop = 1'h0;
				pos_out_fifo_push = ((seg_res_fifo_valid & ~pos_fifo_full) & ~crd_res_fifo_full) & (seg_res_fifo_data_out_0[16] ? 1'h1 : dim_size > num_req_made_crd);
				crd_pop_infifo = 1'h0;
				en_reg_data_in = 1'h0;
				pos_out_to_fifo = (seg_res_fifo_data_out_0[16] ? seg_res_fifo_data_out_0 : sv2v_cast_17((seg_res_fifo_data_out_0[15:0] * dim_size) + num_req_made_crd));
				crd_out_to_fifo = (seg_res_fifo_data_out_0[16] ? seg_res_fifo_data_out_0 : sv2v_cast_17(num_req_made_crd));
				inc_req_made_crd = (((seg_res_fifo_valid & (dim_size > num_req_made_crd)) & ~seg_res_fifo_data_out_0[16]) & ~pos_fifo_full) & ~crd_res_fifo_full;
				clr_req_made_crd = seg_res_fifo_valid & seg_res_fifo_data_out_0[16];
				inc_req_rec_crd = 1'h0;
				clr_req_rec_crd = 1'h0;
				crd_res_fifo_push_alloc = ((seg_res_fifo_valid & ~pos_fifo_full) & ~crd_res_fifo_full) & (seg_res_fifo_data_out_0[16] ? 1'h1 : dim_size > num_req_made_crd);
				crd_res_fifo_push_fill = ((seg_res_fifo_valid & ~pos_fifo_full) & ~crd_res_fifo_full) & (seg_res_fifo_data_out_0[16] ? 1'h1 : dim_size > num_req_made_crd);
				ptr_reg_en = 1'h0;
				seg_res_fifo_pop = ((seg_res_fifo_valid & ~pos_fifo_full) & ~crd_res_fifo_full) & (seg_res_fifo_data_out_0[16] ? 1'h1 : ((dim_size - 16'h0001) == num_req_made_crd) & inc_req_made_crd);
				clr_readout_loop_crd = 1'h0;
				set_readout_loop_crd = 1'h0;
				clr_pushed_done_crd = 1'h0;
				crd_in_done_state = 1'h0;
				set_pushed_done_crd = 1'h0;
			end
			4'h7: begin : scan_seq_crd_DONE_CRD_Output
				crd_addr_out_to_fifo = 16'h0000;
				crd_op_out_to_fifo = 16'h0000;
				crd_ID_out_to_fifo = 16'h0000;
				crd_req_push = 1'h0;
				crd_rd_rsp_fifo_pop = 1'h0;
				pos_out_fifo_push = 1'h0;
				crd_pop_infifo = 1'h0;
				en_reg_data_in = 1'h0;
				pos_out_to_fifo = 17'h00000;
				crd_out_to_fifo = 17'h00000;
				inc_req_made_crd = 1'h0;
				clr_req_made_crd = 1'h1;
				inc_req_rec_crd = 1'h0;
				clr_req_rec_crd = 1'h1;
				crd_res_fifo_push_alloc = 1'h0;
				crd_res_fifo_push_fill = 1'h0;
				ptr_reg_en = 1'h0;
				seg_res_fifo_pop = 1'h0;
				crd_in_done_state = 1'h1;
				set_readout_loop_crd = 1'h0;
				clr_readout_loop_crd = 1'h0;
				clr_pushed_done_crd = 1'h0;
				set_pushed_done_crd = 1'h0;
			end
			4'h8: begin : scan_seq_crd_FREE_CRD_Output
				crd_addr_out_to_fifo = 16'h0000;
				crd_op_out_to_fifo = 16'h0000;
				crd_ID_out_to_fifo = (block_mode ? 16'h0000 : 16'h0001);
				crd_req_push = 1'h1;
				crd_rd_rsp_fifo_pop = 1'h0;
				pos_out_fifo_push = 1'h0;
				crd_pop_infifo = 1'h0;
				en_reg_data_in = 1'h0;
				pos_out_to_fifo = 17'h00000;
				crd_out_to_fifo = 17'h00000;
				inc_req_made_crd = 1'h0;
				clr_req_made_crd = 1'h1;
				inc_req_rec_crd = 1'h0;
				clr_req_rec_crd = 1'h1;
				crd_res_fifo_push_alloc = 1'h0;
				crd_res_fifo_push_fill = 1'h0;
				ptr_reg_en = 1'h0;
				seg_res_fifo_pop = 1'h0;
				clr_readout_loop_crd = 1'h0;
				set_readout_loop_crd = 1'h0;
				clr_pushed_done_crd = 1'h0;
				crd_in_done_state = 1'h0;
				set_pushed_done_crd = 1'h0;
			end
			4'h9: begin : scan_seq_crd_FREE_CRD2_Output
				crd_addr_out_to_fifo = 16'h0000;
				crd_op_out_to_fifo = 16'h0000;
				crd_ID_out_to_fifo = 16'h0001;
				crd_req_push = 1'h1;
				crd_rd_rsp_fifo_pop = 1'h0;
				pos_out_fifo_push = 1'h0;
				crd_pop_infifo = 1'h0;
				en_reg_data_in = 1'h0;
				pos_out_to_fifo = 17'h00000;
				crd_out_to_fifo = 17'h00000;
				inc_req_made_crd = 1'h0;
				clr_req_made_crd = 1'h1;
				inc_req_rec_crd = 1'h0;
				clr_req_rec_crd = 1'h1;
				crd_res_fifo_push_alloc = 1'h0;
				crd_res_fifo_push_fill = 1'h0;
				ptr_reg_en = 1'h0;
				seg_res_fifo_pop = 1'h0;
				clr_readout_loop_crd = 1'h0;
				set_readout_loop_crd = 1'h0;
				clr_pushed_done_crd = 1'h0;
				crd_in_done_state = 1'h0;
				set_pushed_done_crd = 1'h0;
			end
			4'ha: begin : scan_seq_crd_PASS_DONE_CRD_Output
				crd_addr_out_to_fifo = 16'h0000;
				crd_op_out_to_fifo = 16'h0000;
				crd_ID_out_to_fifo = 16'h0000;
				crd_req_push = 1'h0;
				crd_rd_rsp_fifo_pop = 1'h0;
				pos_out_fifo_push = ((~pos_fifo_full & ~crd_res_fifo_full) & seg_res_fifo_done_out) & seg_res_fifo_valid;
				crd_pop_infifo = 1'h0;
				en_reg_data_in = 1'h0;
				pos_out_to_fifo = 17'h10100;
				crd_out_to_fifo = 17'h00000;
				inc_req_made_crd = 1'h0;
				clr_req_made_crd = 1'h0;
				inc_req_rec_crd = 1'h0;
				clr_req_rec_crd = 1'h0;
				crd_res_fifo_push_alloc = ((~pos_fifo_full & ~crd_res_fifo_full) & seg_res_fifo_done_out) & seg_res_fifo_valid;
				crd_res_fifo_push_fill = ((~pos_fifo_full & ~crd_res_fifo_full) & seg_res_fifo_done_out) & seg_res_fifo_valid;
				ptr_reg_en = 1'h0;
				seg_res_fifo_pop = ((~pos_fifo_full & ~crd_res_fifo_full) & seg_res_fifo_done_out) & seg_res_fifo_valid;
				clr_pushed_done_crd = 1'h0;
				clr_readout_loop_crd = 1'h0;
				set_readout_loop_crd = 1'h0;
				crd_in_done_state = 1'h0;
				set_pushed_done_crd = 1'h0;
			end
			4'hb: begin : scan_seq_crd_READOUT_SYNC_LOCK_Output
				crd_addr_out_to_fifo = 16'h0000;
				crd_op_out_to_fifo = 16'h0000;
				crd_ID_out_to_fifo = 16'h0000;
				crd_req_push = 1'h0;
				crd_rd_rsp_fifo_pop = 1'h0;
				pos_out_fifo_push = 1'h0;
				crd_pop_infifo = 1'h0;
				en_reg_data_in = 1'h0;
				pos_out_to_fifo = 17'h00000;
				crd_out_to_fifo = 17'h00000;
				inc_req_made_crd = 1'h0;
				clr_req_made_crd = 1'h0;
				inc_req_rec_crd = 1'h0;
				clr_req_rec_crd = 1'h0;
				crd_res_fifo_push_alloc = 1'h0;
				crd_res_fifo_push_fill = 1'h0;
				ptr_reg_en = 1'h0;
				seg_res_fifo_pop = 1'h0;
				clr_pushed_done_crd = 1'h1;
				clr_readout_loop_crd = 1'h1;
				set_readout_loop_crd = 1'h0;
				crd_in_done_state = 1'h0;
				set_pushed_done_crd = 1'h0;
			end
			4'hc: begin : scan_seq_crd_SEQ_STRM_Output
				crd_addr_out_to_fifo = num_req_made_crd + seg_res_fifo_data_out_0[15:0];
				crd_op_out_to_fifo = 16'h0001;
				crd_ID_out_to_fifo = 16'h0001;
				crd_req_push = (((seg_res_fifo_valid & ~seg_res_fifo_data_out_0[16]) & ~crd_res_fifo_full) & (num_req_made_crd < seq_length_ptr_math)) & ~pos_fifo_full;
				crd_rd_rsp_fifo_pop = 1'h1;
				pos_out_fifo_push = (seg_res_fifo_data_out_0[16] ? (~pos_fifo_full & ~crd_res_fifo_full) & seg_res_fifo_valid : (((crd_grant_push & (num_req_made_crd < seq_length_ptr_math)) & ~pos_fifo_full) & ~crd_res_fifo_full) & seg_res_fifo_valid);
				crd_pop_infifo = 1'h0;
				en_reg_data_in = 1'h0;
				pos_out_to_fifo = (seg_res_fifo_data_out_0[16] ? seg_res_fifo_data_out_0 : {1'h0, num_req_made_crd + seg_res_fifo_data_out_0[15:0]});
				crd_out_to_fifo = 17'h00000;
				inc_req_made_crd = (((crd_grant_push & (num_req_made_crd < seq_length_ptr_math)) & ~pos_fifo_full) & ~crd_res_fifo_full) & seg_res_fifo_valid;
				clr_req_made_crd = ((((crd_grant_push & ((seq_length_ptr_math - 16'h0001) == num_req_made_crd)) | (seq_length_ptr_math == 16'h0000)) & ~pos_fifo_full) & ~crd_res_fifo_full) & seg_res_fifo_valid;
				inc_req_rec_crd = 1'h0;
				clr_req_rec_crd = 1'h0;
				crd_res_fifo_push_alloc = (seg_res_fifo_data_out_0[16] ? (~pos_fifo_full & ~crd_res_fifo_full) & seg_res_fifo_valid : (((crd_grant_push & (num_req_made_crd < seq_length_ptr_math)) & ~pos_fifo_full) & ~crd_res_fifo_full) & seg_res_fifo_valid);
				crd_res_fifo_push_fill = ((seg_res_fifo_valid & seg_res_fifo_data_out_0[16]) & ~pos_fifo_full) & ~crd_res_fifo_full;
				ptr_reg_en = 1'h0;
				seg_res_fifo_pop = clr_req_made_crd | (((seg_res_fifo_valid & seg_res_fifo_data_out_0[16]) & ~pos_fifo_full) & ~crd_res_fifo_full);
				clr_readout_loop_crd = 1'h0;
				set_readout_loop_crd = 1'h0;
				clr_pushed_done_crd = 1'h0;
				crd_in_done_state = 1'h0;
				set_pushed_done_crd = 1'h0;
			end
			4'hd: begin : scan_seq_crd_START_CRD_Output
				crd_addr_out_to_fifo = 16'h0000;
				crd_op_out_to_fifo = 16'h0000;
				crd_ID_out_to_fifo = 16'h0000;
				crd_req_push = 1'h0;
				crd_rd_rsp_fifo_pop = 1'h0;
				pos_out_fifo_push = 1'h0;
				crd_pop_infifo = 1'h0;
				en_reg_data_in = 1'h0;
				pos_out_to_fifo = 17'h00000;
				crd_out_to_fifo = 17'h00000;
				inc_req_made_crd = 1'h0;
				clr_req_made_crd = 1'h0;
				inc_req_rec_crd = 1'h0;
				clr_req_rec_crd = 1'h0;
				crd_res_fifo_push_alloc = 1'h0;
				crd_res_fifo_push_fill = 1'h0;
				ptr_reg_en = 1'h0;
				seg_res_fifo_pop = 1'h0;
				clr_readout_loop_crd = 1'h0;
				set_readout_loop_crd = 1'h0;
				clr_pushed_done_crd = 1'h0;
				crd_in_done_state = 1'h0;
				set_pushed_done_crd = 1'h0;
			end
			default: begin : scan_seq_crd_default_Output
				crd_addr_out_to_fifo = 16'h0000;
				crd_op_out_to_fifo = 16'h0000;
				crd_ID_out_to_fifo = 16'h0000;
				crd_req_push = 1'h0;
				crd_rd_rsp_fifo_pop = 1'h0;
				pos_out_fifo_push = 1'h0;
				crd_pop_infifo = 1'h0;
				en_reg_data_in = 1'h0;
				pos_out_to_fifo = 17'h00000;
				crd_out_to_fifo = 17'h00000;
				inc_req_made_crd = 1'h0;
				clr_req_made_crd = 1'h0;
				inc_req_rec_crd = 1'h0;
				clr_req_rec_crd = 1'h0;
				crd_res_fifo_push_alloc = 1'h0;
				crd_res_fifo_push_fill = 1'h0;
				ptr_reg_en = 1'h0;
				seg_res_fifo_pop = 1'h0;
				clr_readout_loop_crd = 1'h0;
				set_readout_loop_crd = 1'h0;
				clr_pushed_done_crd = 1'h0;
				crd_in_done_state = 1'h0;
				set_pushed_done_crd = 1'h0;
			end
		endcase
	always @(posedge clk or negedge rst_n)
		if (!rst_n)
			scan_seq_seg_current_state <= 4'ha;
		else if (clk_en) begin
			if (flush)
				scan_seq_seg_current_state <= 4'ha;
			else
				scan_seq_seg_current_state <= scan_seq_seg_next_state;
		end
	always @(*) begin
		scan_seq_seg_next_state = scan_seq_seg_current_state;
		case (scan_seq_seg_current_state)
			4'h0:
				if ((lookup ? 1'h1 : ~dense & crd_in_done_state))
					scan_seq_seg_next_state = 4'ha;
			4'h1:
				if (seg_grant_push)
					scan_seq_seg_next_state = 4'h0;
			4'h2: scan_seq_seg_next_state = 4'h3;
			4'h3: scan_seq_seg_next_state = 4'h8;
			4'h4:
				if (~seg_res_fifo_full)
					scan_seq_seg_next_state = 4'h8;
			4'h5:
				if (((done_in & ~spacc_mode) | (((spacc_mode & seg_stop_lvl_geq) & infifo_valid_in) & ~pushed_done_sticky_sticky)) & ~crd_res_fifo_full)
					scan_seq_seg_next_state = 4'h1;
				else
					scan_seq_seg_next_state = 4'h5;
			4'h6:
				if (((readout_loop_sticky_sticky & (~pushed_done_sticky_sticky | ~seg_res_fifo_full)) | ~last_stop_done) | ~seg_res_fifo_full)
					scan_seq_seg_next_state = 4'h1;
			4'h7:
				if (((((infifo_valid_in & ~lookup) & spacc_mode) & seg_stop_lvl_geq) | readout_loop_sticky_sticky) & ~seg_res_fifo_full)
					scan_seq_seg_next_state = 4'h6;
				else if ((infifo_valid_in & ~lookup) & ~seg_res_fifo_full)
					scan_seq_seg_next_state = 4'h8;
				else
					scan_seq_seg_next_state = 4'h7;
			4'h8:
				if ((maybe_in | (((dense & ~done_in) & ~seg_res_fifo_full) & infifo_valid_in)) | ((((~spacc_mode | ~readout_loop_sticky_sticky) & ~dense) & eos_in) & (~spacc_mode | ~use_data_sticky_sticky)))
					scan_seq_seg_next_state = 4'h7;
				else if (seg_grant_push & ~seg_res_fifo_full)
					scan_seq_seg_next_state = 4'h9;
				else if (done_in & ~seg_res_fifo_full)
					scan_seq_seg_next_state = 4'h1;
				else
					scan_seq_seg_next_state = 4'h8;
			4'h9:
				if (seg_grant_push & ~seg_res_fifo_full)
					scan_seq_seg_next_state = 4'h7;
				else
					scan_seq_seg_next_state = 4'h9;
			4'ha:
				if (block_mode)
					scan_seq_seg_next_state = 4'ha;
				else if ((((~root & ~lookup) & ~block_mode) & ~spacc_mode) & tile_en)
					scan_seq_seg_next_state = 4'h8;
				else if (((((~root & ~lookup) & ~block_mode) & (infifo_valid_in | readout_loop_sticky_sticky)) & spacc_mode) & tile_en)
					scan_seq_seg_next_state = 4'h4;
				else if (((root & ~lookup) & ~block_mode) & tile_en)
					scan_seq_seg_next_state = 4'h2;
				else if (((~root & lookup) & ~block_mode) & tile_en)
					scan_seq_seg_next_state = 4'h5;
			default: scan_seq_seg_next_state = scan_seq_seg_current_state;
		endcase
	end
	always @(*)
		case (scan_seq_seg_current_state)
			4'h0: begin : scan_seq_seg_DONE_SEG_Output
				seg_addr_out_to_fifo = 16'h0000;
				seg_op_out_to_fifo = 16'h0000;
				seg_ID_out_to_fifo = 16'h0000;
				seg_req_push = 1'h0;
				seg_rd_rsp_fifo_pop = 1'h1;
				seg_pop_infifo = 1'h0;
				inc_req_made_seg = 1'h0;
				clr_req_made_seg = 1'h0;
				inc_req_rec_seg = 1'h0;
				clr_req_rec_seg = 1'h0;
				us_fifo_inject_data = 16'h0000;
				us_fifo_inject_eos = 1'h0;
				us_fifo_inject_push = 1'h0;
				seg_res_fifo_push_alloc = 1'h0;
				seg_res_fifo_push_fill = 1'h0;
				seg_res_fifo_fill_data_in = 17'h00000;
				set_readout_loop_seg = ((go_to_readout_sticky_sticky & ~readout_loop_sticky_sticky) & spacc_mode) & (crd_in_done_state | lookup);
				clr_readout_loop_seg = (readout_loop_sticky_sticky & spacc_mode) & (crd_in_done_state | lookup);
				seg_in_done_state = 1'h1;
				seg_in_start_state = 1'h0;
				set_pushed_done_seg = 1'h0;
				clr_pushed_done_seg = 1'h0;
			end
			4'h1: begin : scan_seq_seg_FREE_SEG_Output
				seg_addr_out_to_fifo = 16'h0000;
				seg_op_out_to_fifo = 16'h0000;
				seg_ID_out_to_fifo = 16'h0000;
				seg_req_push = 1'h1;
				seg_rd_rsp_fifo_pop = 1'h1;
				seg_pop_infifo = 1'h0;
				inc_req_made_seg = 1'h0;
				clr_req_made_seg = 1'h0;
				inc_req_rec_seg = 1'h0;
				clr_req_rec_seg = 1'h0;
				us_fifo_inject_data = 16'h0000;
				us_fifo_inject_eos = 1'h0;
				us_fifo_inject_push = 1'h0;
				seg_res_fifo_push_alloc = 1'h0;
				seg_res_fifo_push_fill = 1'h0;
				seg_res_fifo_fill_data_in = 17'h00000;
				seg_in_start_state = 1'h0;
				set_readout_loop_seg = 1'h0;
				set_pushed_done_seg = 1'h0;
				clr_pushed_done_seg = 1'h0;
				clr_readout_loop_seg = 1'h0;
				seg_in_done_state = 1'h0;
			end
			4'h2: begin : scan_seq_seg_INJECT_0_Output
				seg_addr_out_to_fifo = 16'h0000;
				seg_op_out_to_fifo = 16'h0000;
				seg_ID_out_to_fifo = 16'h0000;
				seg_req_push = 1'h0;
				seg_rd_rsp_fifo_pop = 1'h0;
				seg_pop_infifo = 1'h0;
				inc_req_made_seg = 1'h0;
				clr_req_made_seg = 1'h0;
				inc_req_rec_seg = 1'h0;
				clr_req_rec_seg = 1'h0;
				us_fifo_inject_data = 16'h0000;
				us_fifo_inject_eos = 1'h0;
				us_fifo_inject_push = 1'h1;
				seg_res_fifo_push_alloc = 1'h0;
				seg_res_fifo_push_fill = 1'h0;
				seg_res_fifo_fill_data_in = 17'h00000;
				seg_in_start_state = 1'h0;
				set_readout_loop_seg = 1'h0;
				set_pushed_done_seg = 1'h0;
				clr_pushed_done_seg = 1'h0;
				clr_readout_loop_seg = 1'h0;
				seg_in_done_state = 1'h0;
			end
			4'h3: begin : scan_seq_seg_INJECT_DONE_Output
				seg_addr_out_to_fifo = 16'h0000;
				seg_op_out_to_fifo = 16'h0000;
				seg_ID_out_to_fifo = 16'h0000;
				seg_req_push = 1'h0;
				seg_rd_rsp_fifo_pop = 1'h0;
				seg_pop_infifo = 1'h0;
				inc_req_made_seg = 1'h0;
				clr_req_made_seg = 1'h0;
				inc_req_rec_seg = 1'h0;
				clr_req_rec_seg = 1'h0;
				us_fifo_inject_data = 16'h0100;
				us_fifo_inject_eos = 1'h1;
				us_fifo_inject_push = 1'h1;
				seg_res_fifo_push_alloc = 1'h0;
				seg_res_fifo_push_fill = 1'h0;
				seg_res_fifo_fill_data_in = 17'h00000;
				seg_in_start_state = 1'h0;
				set_readout_loop_seg = 1'h0;
				set_pushed_done_seg = 1'h0;
				clr_pushed_done_seg = 1'h0;
				clr_readout_loop_seg = 1'h0;
				seg_in_done_state = 1'h0;
			end
			4'h4: begin : scan_seq_seg_INJECT_ROUTING_Output
				seg_addr_out_to_fifo = 16'h0000;
				seg_op_out_to_fifo = 16'h0000;
				seg_ID_out_to_fifo = 16'h0000;
				seg_req_push = 1'h0;
				seg_rd_rsp_fifo_pop = 1'h0;
				seg_pop_infifo = 1'h0;
				inc_req_made_seg = 1'h0;
				clr_req_made_seg = 1'h0;
				inc_req_rec_seg = 1'h0;
				clr_req_rec_seg = 1'h0;
				us_fifo_inject_data = 16'h0000;
				us_fifo_inject_eos = 1'h0;
				us_fifo_inject_push = 1'h1;
				seg_res_fifo_push_alloc = ~seg_res_fifo_full;
				seg_res_fifo_push_fill = ~seg_res_fifo_full;
				seg_res_fifo_fill_data_in = {16'h8180, readout_loop_sticky_sticky};
				seg_in_start_state = 1'h0;
				set_readout_loop_seg = 1'h0;
				set_pushed_done_seg = 1'h0;
				clr_pushed_done_seg = 1'h0;
				clr_readout_loop_seg = 1'h0;
				seg_in_done_state = 1'h0;
			end
			4'h5: begin : scan_seq_seg_LOOKUP_Output
				seg_addr_out_to_fifo = infifo_pos_in;
				seg_op_out_to_fifo = 16'h0001;
				seg_ID_out_to_fifo = 16'h0000;
				seg_req_push = (infifo_valid_in & ~infifo_eos_in) & ~crd_res_fifo_full;
				seg_rd_rsp_fifo_pop = 1'h1;
				seg_pop_infifo = (infifo_valid_in & ~crd_res_fifo_full) & (infifo_eos_in ? 1'h1 : seg_grant_push);
				inc_req_made_seg = 1'h0;
				clr_req_made_seg = 1'h1;
				inc_req_rec_seg = 1'h0;
				clr_req_rec_seg = 1'h1;
				us_fifo_inject_data = 16'h0000;
				us_fifo_inject_eos = 1'h0;
				us_fifo_inject_push = 1'h0;
				seg_res_fifo_push_alloc = ~crd_res_fifo_full & (seg_grant_push | (infifo_valid_in & infifo_eos_in));
				seg_res_fifo_push_fill = (infifo_valid_in & infifo_eos_in) & ~crd_res_fifo_full;
				seg_res_fifo_fill_data_in = (infifo_eos_in & (infifo_pos_in[9:8] == 2'h2) ? 17'h00000 : {infifo_eos_in, infifo_pos_in});
				set_pushed_done_seg = (done_in & ~crd_res_fifo_full) & spacc_mode;
				set_readout_loop_seg = (done_in & ~crd_res_fifo_full) & spacc_mode;
				seg_in_start_state = 1'h0;
				clr_pushed_done_seg = 1'h0;
				clr_readout_loop_seg = 1'h0;
				seg_in_done_state = 1'h0;
			end
			4'h6: begin : scan_seq_seg_PASS_DONE_SEG_Output
				seg_addr_out_to_fifo = 16'h0000;
				seg_op_out_to_fifo = 16'h0000;
				seg_ID_out_to_fifo = 16'h0000;
				seg_req_push = 1'h0;
				seg_rd_rsp_fifo_pop = 1'h1;
				seg_pop_infifo = (~readout_loop_sticky_sticky & done_in) & ~seg_res_fifo_full;
				inc_req_made_seg = 1'h0;
				clr_req_made_seg = 1'h0;
				inc_req_rec_seg = 1'h0;
				clr_req_rec_seg = 1'h0;
				us_fifo_inject_data = 16'h0000;
				us_fifo_inject_eos = 1'h0;
				us_fifo_inject_push = 1'h0;
				seg_res_fifo_push_alloc = ((readout_loop_sticky_sticky & pushed_done_sticky_sticky) | (~readout_loop_sticky_sticky & last_stop_done)) & ~seg_res_fifo_full;
				seg_res_fifo_push_fill = ((readout_loop_sticky_sticky & pushed_done_sticky_sticky) | (~readout_loop_sticky_sticky & last_stop_done)) & ~seg_res_fifo_full;
				seg_res_fifo_fill_data_in = 17'h10100;
				set_pushed_done_seg = (last_stop_done & ~seg_res_fifo_full) & spacc_mode;
				seg_in_start_state = 1'h0;
				set_readout_loop_seg = 1'h0;
				clr_pushed_done_seg = 1'h0;
				clr_readout_loop_seg = 1'h0;
				seg_in_done_state = 1'h0;
			end
			4'h7: begin : scan_seq_seg_PASS_STOP_SEG_Output
				seg_addr_out_to_fifo = 16'h0000;
				seg_op_out_to_fifo = 16'h0000;
				seg_ID_out_to_fifo = 16'h0000;
				seg_req_push = 1'h0;
				seg_rd_rsp_fifo_pop = 1'h1;
				seg_pop_infifo = (~seg_res_fifo_full & eos_in) & ~readout_loop_sticky_sticky;
				inc_req_made_seg = 1'h0;
				clr_req_made_seg = 1'h1;
				inc_req_rec_seg = 1'h0;
				clr_req_rec_seg = 1'h1;
				us_fifo_inject_data = 16'h0000;
				us_fifo_inject_eos = 1'h0;
				us_fifo_inject_push = 1'h0;
				seg_res_fifo_push_alloc = (infifo_valid_in | readout_loop_sticky_sticky) & ~seg_res_fifo_full;
				seg_res_fifo_push_fill = (infifo_valid_in | readout_loop_sticky_sticky) & ~seg_res_fifo_full;
				seg_res_fifo_fill_data_in = (readout_loop_sticky_sticky ? last_stop_token - 17'h00001 : (eos_in ? {1'h1, infifo_pos_in + 16'h0001} : 17'h10000));
				seg_in_start_state = 1'h0;
				set_readout_loop_seg = 1'h0;
				set_pushed_done_seg = 1'h0;
				clr_pushed_done_seg = 1'h0;
				clr_readout_loop_seg = 1'h0;
				seg_in_done_state = 1'h0;
			end
			4'h8: begin : scan_seq_seg_READ_Output
				seg_addr_out_to_fifo = (readout_loop_sticky_sticky ? 16'h0000 : infifo_pos_in);
				seg_op_out_to_fifo = 16'h0001;
				seg_ID_out_to_fifo = 16'h0000;
				seg_req_push = (((infifo_valid_in & ~infifo_eos_in) & ~dense) | readout_loop_sticky_sticky) & ~seg_res_fifo_full;
				seg_rd_rsp_fifo_pop = 1'h1;
				seg_pop_infifo = (((done_in | (dense & infifo_valid_in)) & ~seg_res_fifo_full) | maybe_in) & ~readout_loop_sticky_sticky;
				inc_req_made_seg = 1'h0;
				clr_req_made_seg = 1'h0;
				inc_req_rec_seg = 1'h0;
				clr_req_rec_seg = 1'h0;
				us_fifo_inject_data = 16'h0000;
				us_fifo_inject_eos = 1'h0;
				us_fifo_inject_push = 1'h0;
				seg_res_fifo_push_alloc = (done_in | dense ? ~seg_res_fifo_full & infifo_valid_in : (~seg_res_fifo_full & seg_grant_push) & ~maybe_in);
				seg_res_fifo_push_fill = (done_in | (dense & infifo_valid_in)) & ~seg_res_fifo_full;
				seg_res_fifo_fill_data_in = {infifo_eos_in, infifo_pos_in};
				seg_in_start_state = 1'h0;
				set_readout_loop_seg = 1'h0;
				set_pushed_done_seg = 1'h0;
				clr_pushed_done_seg = 1'h0;
				clr_readout_loop_seg = 1'h0;
				seg_in_done_state = 1'h0;
			end
			4'h9: begin : scan_seq_seg_READ_ALT_Output
				seg_addr_out_to_fifo = (readout_loop_sticky_sticky ? 16'h0001 : infifo_pos_in + 16'h0001);
				seg_op_out_to_fifo = 16'h0001;
				seg_ID_out_to_fifo = 16'h0000;
				seg_req_push = ~seg_res_fifo_full;
				seg_rd_rsp_fifo_pop = 1'h1;
				seg_pop_infifo = (seg_grant_push & ~seg_res_fifo_full) & ~readout_loop_sticky_sticky;
				inc_req_made_seg = 1'h0;
				clr_req_made_seg = 1'h0;
				inc_req_rec_seg = 1'h0;
				clr_req_rec_seg = 1'h0;
				us_fifo_inject_data = 16'h0000;
				us_fifo_inject_eos = 1'h0;
				us_fifo_inject_push = 1'h0;
				seg_res_fifo_push_alloc = 1'h0;
				seg_res_fifo_push_fill = 1'h0;
				seg_res_fifo_fill_data_in = 17'h00000;
				seg_in_start_state = 1'h0;
				set_readout_loop_seg = 1'h0;
				set_pushed_done_seg = 1'h0;
				clr_pushed_done_seg = 1'h0;
				clr_readout_loop_seg = 1'h0;
				seg_in_done_state = 1'h0;
			end
			4'ha: begin : scan_seq_seg_START_SEG_Output
				seg_addr_out_to_fifo = 16'h0000;
				seg_op_out_to_fifo = 16'h0000;
				seg_ID_out_to_fifo = 16'h0000;
				seg_req_push = 1'h0;
				seg_rd_rsp_fifo_pop = 1'h0;
				seg_pop_infifo = 1'h0;
				inc_req_made_seg = 1'h0;
				clr_req_made_seg = 1'h0;
				inc_req_rec_seg = 1'h0;
				clr_req_rec_seg = 1'h0;
				us_fifo_inject_data = 16'h0000;
				us_fifo_inject_eos = 1'h0;
				us_fifo_inject_push = 1'h0;
				seg_res_fifo_push_alloc = 1'h0;
				seg_res_fifo_push_fill = 1'h0;
				seg_res_fifo_fill_data_in = 17'h00000;
				set_readout_loop_seg = 1'h0;
				seg_in_start_state = 1'h1;
				set_pushed_done_seg = 1'h0;
				clr_pushed_done_seg = 1'h0;
				clr_readout_loop_seg = 1'h0;
				seg_in_done_state = 1'h0;
			end
			default: begin : scan_seq_seg_default_Output
				seg_addr_out_to_fifo = 16'h0000;
				seg_op_out_to_fifo = 16'h0000;
				seg_ID_out_to_fifo = 16'h0000;
				seg_req_push = 1'h0;
				seg_rd_rsp_fifo_pop = 1'h0;
				seg_pop_infifo = 1'h0;
				inc_req_made_seg = 1'h0;
				clr_req_made_seg = 1'h0;
				inc_req_rec_seg = 1'h0;
				clr_req_rec_seg = 1'h0;
				us_fifo_inject_data = 16'h0000;
				us_fifo_inject_eos = 1'h0;
				us_fifo_inject_push = 1'h0;
				seg_res_fifo_push_alloc = 1'h0;
				seg_res_fifo_push_fill = 1'h0;
				seg_res_fifo_fill_data_in = 17'h00000;
				set_readout_loop_seg = 1'h0;
				seg_in_start_state = 1'h1;
				set_pushed_done_seg = 1'h0;
				clr_pushed_done_seg = 1'h0;
				clr_readout_loop_seg = 1'h0;
				seg_in_done_state = 1'h0;
			end
		endcase
	reg_fifo_depth_2_w_17_afd_2 input_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(fifo_us_in_packed),
		.flush(flush),
		.pop(pop_infifo),
		.push(us_fifo_push),
		.rst_n(rst_n),
		.data_out(input_fifo_data_out),
		.empty(input_fifo_empty),
		.full(fifo_us_full)
	);
	reg_fifo_depth_2_w_17_afd_2 rd_rsp_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(rd_rsp_data_in[0+:17]),
		.flush(flush),
		.pop(1'h1),
		.push(rd_rsp_data_in_valid),
		.rst_n(rst_n),
		.data_out(rd_rsp_fifo_out_data),
		.empty(rd_rsp_fifo_empty),
		.full(rd_rsp_fifo_full)
	);
	arbiter_2_in_PRIO_algo rr_arbiter(
		.clk(gclk),
		.clk_en(clk_en),
		.flush(flush),
		.request_in(base_rr),
		.resource_ready(no_outfifo_full),
		.rst_n(rst_n),
		.grant_out(rr_arbiter_grant_out)
	);
	reg_fifo_depth_2_w_17_afd_2 addr_out_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(addr_out_fifo_data_in),
		.flush(flush),
		.pop(addr_out_ready),
		.push(addr_out_fifo_push),
		.rst_n(rst_n),
		.data_out(addr_out),
		.empty(addr_out_fifo_empty),
		.full(addr_out_fifo_full)
	);
	reg_fifo_depth_2_w_17_afd_2 op_out_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(op_out_fifo_data_in),
		.flush(flush),
		.pop(op_out_ready),
		.push(op_out_fifo_push),
		.rst_n(rst_n),
		.data_out(op_out),
		.empty(op_out_fifo_empty),
		.full(op_out_fifo_full)
	);
	reg_fifo_depth_2_w_17_afd_2 ID_out_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(ID_out_fifo_data_in),
		.flush(flush),
		.pop(ID_out_ready),
		.push(ID_out_fifo_push),
		.rst_n(rst_n),
		.data_out(ID_out),
		.empty(ID_out_fifo_empty),
		.full(ID_out_fifo_full)
	);
	reservation_fifo_depth_8_w_17_num_per_2 seg_res_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in_0(rd_rsp_fifo_out_data),
		.data_in_1(rd_rsp_fifo_out_data),
		.fill_data_in(seg_res_fifo_fill_data_in),
		.flush(flush),
		.pop(seg_res_fifo_pop_0),
		.push_alloc(seg_res_fifo_push_alloc_0),
		.push_fill(seg_res_fifo_push_fill_0),
		.push_reserve(seg_res_fifo_push_reserve_0),
		.rst_n(rst_n),
		.data_out_0(seg_res_fifo_data_out_0),
		.data_out_1(seg_res_fifo_data_out_1),
		.full(seg_res_fifo_full),
		.valid(seg_res_fifo_valid)
	);
	reservation_fifo_depth_8_w_17_num_per_1 crd_res_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in_0(crd_res_fifo_data_in_0),
		.fill_data_in(crd_res_fifo_fill_data_in),
		.flush(flush),
		.pop(crd_res_fifo_pop),
		.push_alloc(crd_res_fifo_push_alloc_0),
		.push_fill(crd_res_fifo_push_fill_0),
		.push_reserve(crd_res_fifo_push_reserve_0),
		.rst_n(rst_n),
		.data_out_0(crd_res_fifo_data_out),
		.full(crd_res_fifo_full),
		.valid(crd_res_fifo_valid)
	);
	reg_fifo_depth_0_w_17_afd_2 coordinate_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(coord_fifo_in_packed),
		.flush(flush),
		.pop(coord_out_ready),
		.push(coordinate_fifo_push),
		.rst_n(rst_n),
		.data_out(coord_fifo_out_packed),
		.empty(coordinate_fifo_empty),
		.full(coordinate_fifo_full)
	);
	reg_fifo_depth_0_w_17_afd_2 pos_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(pos_fifo_in_packed),
		.flush(flush),
		.pop(pos_out_ready),
		.push(pos_out_fifo_push),
		.rst_n(rst_n),
		.data_out(pos_fifo_out_packed),
		.empty(pos_fifo_empty),
		.full(pos_fifo_full)
	);
	reg_fifo_depth_0_w_17_afd_2 block_rd_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(crd_res_fifo_data_out),
		.flush(flush),
		.pop(block_rd_out_ready),
		.push(block_rd_fifo_push),
		.rst_n(rst_n),
		.data_out(block_rd_out),
		.empty(block_rd_fifo_empty),
		.full(block_rd_fifo_full)
	);
endmodule
module sched_gen_3_16 (
	clk,
	clk_en,
	cycle_count,
	enable,
	finished,
	flush,
	mux_sel,
	rst_n,
	sched_addr_gen_starting_addr,
	sched_addr_gen_strides_0,
	sched_addr_gen_strides_1,
	sched_addr_gen_strides_2,
	valid_output
);
	input wire clk;
	input wire clk_en;
	input wire [15:0] cycle_count;
	input wire enable;
	input wire finished;
	input wire flush;
	input wire [1:0] mux_sel;
	input wire rst_n;
	input wire [15:0] sched_addr_gen_starting_addr;
	input wire [15:0] sched_addr_gen_strides_0;
	input wire [15:0] sched_addr_gen_strides_1;
	input wire [15:0] sched_addr_gen_strides_2;
	output reg valid_output;
	wire [15:0] addr_out;
	wire [47:0] sched_addr_gen_strides;
	wire valid_gate;
	reg valid_gate_inv;
	reg valid_out;
	assign valid_gate = ~valid_gate_inv;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			valid_gate_inv <= 1'h0;
		else if (clk_en) begin
			if (flush)
				valid_gate_inv <= 1'h0;
			else if (finished)
				valid_gate_inv <= 1'h1;
		end
	always @(*) valid_out = ((cycle_count == addr_out) & valid_gate) & enable;
	always @(*) valid_output = valid_out;
	assign sched_addr_gen_strides[0+:16] = sched_addr_gen_strides_0;
	assign sched_addr_gen_strides[16+:16] = sched_addr_gen_strides_1;
	assign sched_addr_gen_strides[32+:16] = sched_addr_gen_strides_2;
	addr_gen_3_16 sched_addr_gen(
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.mux_sel(mux_sel),
		.restart(finished),
		.rst_n(rst_n),
		.starting_addr(sched_addr_gen_starting_addr),
		.step(valid_out),
		.strides(sched_addr_gen_strides),
		.addr_out(addr_out)
	);
endmodule
module sched_gen_6_16 (
	clk,
	clk_en,
	cycle_count,
	enable,
	finished,
	flush,
	mux_sel,
	rst_n,
	sched_addr_gen_starting_addr,
	sched_addr_gen_strides_0,
	sched_addr_gen_strides_1,
	sched_addr_gen_strides_2,
	sched_addr_gen_strides_3,
	sched_addr_gen_strides_4,
	sched_addr_gen_strides_5,
	valid_output
);
	input wire clk;
	input wire clk_en;
	input wire [15:0] cycle_count;
	input wire enable;
	input wire finished;
	input wire flush;
	input wire [2:0] mux_sel;
	input wire rst_n;
	input wire [15:0] sched_addr_gen_starting_addr;
	input wire [15:0] sched_addr_gen_strides_0;
	input wire [15:0] sched_addr_gen_strides_1;
	input wire [15:0] sched_addr_gen_strides_2;
	input wire [15:0] sched_addr_gen_strides_3;
	input wire [15:0] sched_addr_gen_strides_4;
	input wire [15:0] sched_addr_gen_strides_5;
	output reg valid_output;
	wire [15:0] addr_out;
	wire [95:0] sched_addr_gen_strides;
	wire valid_gate;
	reg valid_gate_inv;
	reg valid_out;
	assign valid_gate = ~valid_gate_inv;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			valid_gate_inv <= 1'h0;
		else if (clk_en) begin
			if (flush)
				valid_gate_inv <= 1'h0;
			else if (finished)
				valid_gate_inv <= 1'h1;
		end
	always @(*) valid_out = ((cycle_count == addr_out) & valid_gate) & enable;
	always @(*) valid_output = valid_out;
	assign sched_addr_gen_strides[0+:16] = sched_addr_gen_strides_0;
	assign sched_addr_gen_strides[16+:16] = sched_addr_gen_strides_1;
	assign sched_addr_gen_strides[32+:16] = sched_addr_gen_strides_2;
	assign sched_addr_gen_strides[48+:16] = sched_addr_gen_strides_3;
	assign sched_addr_gen_strides[64+:16] = sched_addr_gen_strides_4;
	assign sched_addr_gen_strides[80+:16] = sched_addr_gen_strides_5;
	addr_gen_6_16 sched_addr_gen(
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.mux_sel(mux_sel),
		.restart(finished),
		.rst_n(rst_n),
		.starting_addr(sched_addr_gen_starting_addr),
		.step(valid_out),
		.strides(sched_addr_gen_strides),
		.addr_out(addr_out)
	);
endmodule
module sched_gen_6_16_delay_addr_10_4 (
	clk,
	clk_en,
	cycle_count,
	enable,
	finished,
	flush,
	mux_sel,
	rst_n,
	sched_addr_gen_delay,
	sched_addr_gen_starting_addr,
	sched_addr_gen_strides_0,
	sched_addr_gen_strides_1,
	sched_addr_gen_strides_2,
	sched_addr_gen_strides_3,
	sched_addr_gen_strides_4,
	sched_addr_gen_strides_5,
	delay_en_out,
	valid_output,
	valid_output_d
);
	input wire clk;
	input wire clk_en;
	input wire [15:0] cycle_count;
	input wire enable;
	input wire finished;
	input wire flush;
	input wire [2:0] mux_sel;
	input wire rst_n;
	input wire [9:0] sched_addr_gen_delay;
	input wire [15:0] sched_addr_gen_starting_addr;
	input wire [15:0] sched_addr_gen_strides_0;
	input wire [15:0] sched_addr_gen_strides_1;
	input wire [15:0] sched_addr_gen_strides_2;
	input wire [15:0] sched_addr_gen_strides_3;
	input wire [15:0] sched_addr_gen_strides_4;
	input wire [15:0] sched_addr_gen_strides_5;
	output wire delay_en_out;
	output reg valid_output;
	output reg valid_output_d;
	reg [43:0] addr_fifo;
	reg addr_fifo_empty_n;
	wire [10:0] addr_fifo_in;
	wire [10:0] addr_fifo_out;
	wire addr_fifo_wr_en;
	wire [15:0] addr_out;
	wire [15:0] addr_out_d;
	wire delay_en;
	wire [1:0] next_rd_ptr;
	reg [1:0] rd_ptr;
	wire [9:0] sched_addr_gen_delay_out;
	wire [95:0] sched_addr_gen_strides;
	wire valid_gate;
	reg valid_gate_inv;
	reg valid_out;
	reg valid_out_d;
	reg [1:0] wr_ptr;
	assign valid_gate = ~valid_gate_inv;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			valid_gate_inv <= 1'h0;
		else if (clk_en) begin
			if (flush)
				valid_gate_inv <= 1'h0;
			else if (finished)
				valid_gate_inv <= 1'h1;
		end
	assign delay_en_out = delay_en;
	assign delay_en = sched_addr_gen_delay_out > 10'h000;
	assign next_rd_ptr = rd_ptr + 2'h1;
	assign addr_fifo_wr_en = valid_out;
	assign addr_fifo_in = addr_out_d[10:0];
	assign addr_fifo_out = addr_fifo[rd_ptr * 11+:11];
	always @(posedge clk or negedge rst_n)
		if (~rst_n) begin
			wr_ptr <= 2'h0;
			rd_ptr <= 2'h0;
			addr_fifo <= 44'h00000000000;
			addr_fifo_empty_n <= 1'h0;
		end
		else if (clk_en) begin
			if (flush) begin
				wr_ptr <= 2'h0;
				rd_ptr <= 2'h0;
				addr_fifo <= 44'h00000000000;
				addr_fifo_empty_n <= 1'h0;
			end
			else if (delay_en) begin
				if (addr_fifo_wr_en) begin
					wr_ptr <= wr_ptr + 2'h1;
					addr_fifo[wr_ptr * 11+:11] <= addr_fifo_in;
				end
				if (valid_out_d)
					rd_ptr <= next_rd_ptr;
				if (addr_fifo_wr_en)
					addr_fifo_empty_n <= 1'h1;
				else if (valid_out_d)
					addr_fifo_empty_n <= ~(next_rd_ptr == wr_ptr);
				else
					addr_fifo_empty_n <= addr_fifo_empty_n;
			end
		end
	always @(*) begin
		valid_out_d = ((cycle_count[10:0] == addr_fifo_out) & addr_fifo_empty_n) & enable;
		valid_output_d = valid_out_d;
	end
	always @(*) valid_out = ((cycle_count == addr_out) & valid_gate) & enable;
	always @(*) valid_output = valid_out;
	assign sched_addr_gen_strides[0+:16] = sched_addr_gen_strides_0;
	assign sched_addr_gen_strides[16+:16] = sched_addr_gen_strides_1;
	assign sched_addr_gen_strides[32+:16] = sched_addr_gen_strides_2;
	assign sched_addr_gen_strides[48+:16] = sched_addr_gen_strides_3;
	assign sched_addr_gen_strides[64+:16] = sched_addr_gen_strides_4;
	assign sched_addr_gen_strides[80+:16] = sched_addr_gen_strides_5;
	addr_gen_6_16_delay_addr_10 sched_addr_gen(
		.clk(clk),
		.clk_en(clk_en),
		.delay(sched_addr_gen_delay),
		.flush(flush),
		.mux_sel(mux_sel),
		.restart(finished),
		.rst_n(rst_n),
		.starting_addr(sched_addr_gen_starting_addr),
		.step(valid_out),
		.strides(sched_addr_gen_strides),
		.addr_out(addr_out),
		.delay_out(sched_addr_gen_delay_out),
		.delayed_addr_out(addr_out_d)
	);
endmodule
module sched_gen_6_16_delay_addr_10_8 (
	clk,
	clk_en,
	cycle_count,
	enable,
	finished,
	flush,
	mux_sel,
	rst_n,
	sched_addr_gen_delay,
	sched_addr_gen_starting_addr,
	sched_addr_gen_strides_0,
	sched_addr_gen_strides_1,
	sched_addr_gen_strides_2,
	sched_addr_gen_strides_3,
	sched_addr_gen_strides_4,
	sched_addr_gen_strides_5,
	delay_en_out,
	valid_output,
	valid_output_d
);
	input wire clk;
	input wire clk_en;
	input wire [15:0] cycle_count;
	input wire enable;
	input wire finished;
	input wire flush;
	input wire [2:0] mux_sel;
	input wire rst_n;
	input wire [9:0] sched_addr_gen_delay;
	input wire [15:0] sched_addr_gen_starting_addr;
	input wire [15:0] sched_addr_gen_strides_0;
	input wire [15:0] sched_addr_gen_strides_1;
	input wire [15:0] sched_addr_gen_strides_2;
	input wire [15:0] sched_addr_gen_strides_3;
	input wire [15:0] sched_addr_gen_strides_4;
	input wire [15:0] sched_addr_gen_strides_5;
	output wire delay_en_out;
	output reg valid_output;
	output reg valid_output_d;
	reg [87:0] addr_fifo;
	reg addr_fifo_empty_n;
	wire [10:0] addr_fifo_in;
	wire [10:0] addr_fifo_out;
	wire addr_fifo_wr_en;
	wire [15:0] addr_out;
	wire [15:0] addr_out_d;
	wire delay_en;
	wire [2:0] next_rd_ptr;
	reg [2:0] rd_ptr;
	wire [9:0] sched_addr_gen_delay_out;
	wire [95:0] sched_addr_gen_strides;
	wire valid_gate;
	reg valid_gate_inv;
	reg valid_out;
	reg valid_out_d;
	reg [2:0] wr_ptr;
	assign valid_gate = ~valid_gate_inv;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			valid_gate_inv <= 1'h0;
		else if (clk_en) begin
			if (flush)
				valid_gate_inv <= 1'h0;
			else if (finished)
				valid_gate_inv <= 1'h1;
		end
	assign delay_en_out = delay_en;
	assign delay_en = sched_addr_gen_delay_out > 10'h000;
	assign next_rd_ptr = rd_ptr + 3'h1;
	assign addr_fifo_wr_en = valid_out;
	assign addr_fifo_in = addr_out_d[10:0];
	assign addr_fifo_out = addr_fifo[rd_ptr * 11+:11];
	always @(posedge clk or negedge rst_n)
		if (~rst_n) begin
			wr_ptr <= 3'h0;
			rd_ptr <= 3'h0;
			addr_fifo <= 88'h0000000000000000000000;
			addr_fifo_empty_n <= 1'h0;
		end
		else if (clk_en) begin
			if (flush) begin
				wr_ptr <= 3'h0;
				rd_ptr <= 3'h0;
				addr_fifo <= 88'h0000000000000000000000;
				addr_fifo_empty_n <= 1'h0;
			end
			else if (delay_en) begin
				if (addr_fifo_wr_en) begin
					wr_ptr <= wr_ptr + 3'h1;
					addr_fifo[wr_ptr * 11+:11] <= addr_fifo_in;
				end
				if (valid_out_d)
					rd_ptr <= next_rd_ptr;
				if (addr_fifo_wr_en)
					addr_fifo_empty_n <= 1'h1;
				else if (valid_out_d)
					addr_fifo_empty_n <= ~(next_rd_ptr == wr_ptr);
				else
					addr_fifo_empty_n <= addr_fifo_empty_n;
			end
		end
	always @(*) begin
		valid_out_d = ((cycle_count[10:0] == addr_fifo_out) & addr_fifo_empty_n) & enable;
		valid_output_d = valid_out_d;
	end
	always @(*) valid_out = ((cycle_count == addr_out) & valid_gate) & enable;
	always @(*) valid_output = valid_out;
	assign sched_addr_gen_strides[0+:16] = sched_addr_gen_strides_0;
	assign sched_addr_gen_strides[16+:16] = sched_addr_gen_strides_1;
	assign sched_addr_gen_strides[32+:16] = sched_addr_gen_strides_2;
	assign sched_addr_gen_strides[48+:16] = sched_addr_gen_strides_3;
	assign sched_addr_gen_strides[64+:16] = sched_addr_gen_strides_4;
	assign sched_addr_gen_strides[80+:16] = sched_addr_gen_strides_5;
	addr_gen_6_16_delay_addr_10 sched_addr_gen(
		.clk(clk),
		.clk_en(clk_en),
		.delay(sched_addr_gen_delay),
		.flush(flush),
		.mux_sel(mux_sel),
		.restart(finished),
		.rst_n(rst_n),
		.starting_addr(sched_addr_gen_starting_addr),
		.step(valid_out),
		.strides(sched_addr_gen_strides),
		.addr_out(addr_out),
		.delay_out(sched_addr_gen_delay_out),
		.delayed_addr_out(addr_out_d)
	);
endmodule
module sram_sp__0 (
	clk,
	clk_en,
	data_in_p0,
	flush,
	read_addr_p0,
	read_enable_p0,
	write_addr_p0,
	write_enable_p0,
	data_out_p0
);
	input wire clk;
	input wire clk_en;
	input wire [63:0] data_in_p0;
	input wire flush;
	input wire [8:0] read_addr_p0;
	input wire read_enable_p0;
	input wire [8:0] write_addr_p0;
	input wire write_enable_p0;
	output reg [63:0] data_out_p0;
	reg [63:0] data_array [511:0];
	always @(posedge clk)
		if (clk_en) begin
			if (write_enable_p0 == 1'h1)
				data_array[write_addr_p0] <= data_in_p0;
			else if (read_enable_p0)
				data_out_p0 <= data_array[read_addr_p0];
		end
endmodule
module stencil_valid (
	clk,
	clk_en,
	flush,
	loops_stencil_valid_dimensionality,
	loops_stencil_valid_ranges_0,
	loops_stencil_valid_ranges_1,
	loops_stencil_valid_ranges_2,
	loops_stencil_valid_ranges_3,
	loops_stencil_valid_ranges_4,
	loops_stencil_valid_ranges_5,
	rst_n,
	stencil_valid_sched_gen_enable,
	stencil_valid_sched_gen_sched_addr_gen_starting_addr,
	stencil_valid_sched_gen_sched_addr_gen_strides_0,
	stencil_valid_sched_gen_sched_addr_gen_strides_1,
	stencil_valid_sched_gen_sched_addr_gen_strides_2,
	stencil_valid_sched_gen_sched_addr_gen_strides_3,
	stencil_valid_sched_gen_sched_addr_gen_strides_4,
	stencil_valid_sched_gen_sched_addr_gen_strides_5,
	stencil_valid
);
	input wire clk;
	input wire clk_en;
	input wire flush;
	input wire [3:0] loops_stencil_valid_dimensionality;
	input wire [10:0] loops_stencil_valid_ranges_0;
	input wire [10:0] loops_stencil_valid_ranges_1;
	input wire [10:0] loops_stencil_valid_ranges_2;
	input wire [10:0] loops_stencil_valid_ranges_3;
	input wire [10:0] loops_stencil_valid_ranges_4;
	input wire [10:0] loops_stencil_valid_ranges_5;
	input wire rst_n;
	input wire stencil_valid_sched_gen_enable;
	input wire [15:0] stencil_valid_sched_gen_sched_addr_gen_starting_addr;
	input wire [15:0] stencil_valid_sched_gen_sched_addr_gen_strides_0;
	input wire [15:0] stencil_valid_sched_gen_sched_addr_gen_strides_1;
	input wire [15:0] stencil_valid_sched_gen_sched_addr_gen_strides_2;
	input wire [15:0] stencil_valid_sched_gen_sched_addr_gen_strides_3;
	input wire [15:0] stencil_valid_sched_gen_sched_addr_gen_strides_4;
	input wire [15:0] stencil_valid_sched_gen_sched_addr_gen_strides_5;
	output wire stencil_valid;
	reg [15:0] cycle_count;
	reg flushed;
	wire [2:0] loops_stencil_valid_mux_sel_out;
	wire [65:0] loops_stencil_valid_ranges;
	wire loops_stencil_valid_restart;
	wire stencil_valid_internal;
	assign stencil_valid = stencil_valid_internal & flushed;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			cycle_count <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				cycle_count <= 16'h0000;
			else if (flushed)
				cycle_count <= cycle_count + 16'h0001;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			flushed <= 1'h0;
		else if (clk_en) begin
			if (flush)
				flushed <= 1'h1;
		end
	assign loops_stencil_valid_ranges[0+:11] = loops_stencil_valid_ranges_0;
	assign loops_stencil_valid_ranges[11+:11] = loops_stencil_valid_ranges_1;
	assign loops_stencil_valid_ranges[22+:11] = loops_stencil_valid_ranges_2;
	assign loops_stencil_valid_ranges[33+:11] = loops_stencil_valid_ranges_3;
	assign loops_stencil_valid_ranges[44+:11] = loops_stencil_valid_ranges_4;
	assign loops_stencil_valid_ranges[55+:11] = loops_stencil_valid_ranges_5;
	for_loop_6_11 loops_stencil_valid(
		.clk(clk),
		.clk_en(clk_en),
		.dimensionality(loops_stencil_valid_dimensionality),
		.flush(flush),
		.ranges(loops_stencil_valid_ranges),
		.rst_n(rst_n),
		.step(stencil_valid_internal),
		.mux_sel_out(loops_stencil_valid_mux_sel_out),
		.restart(loops_stencil_valid_restart)
	);
	sched_gen_6_16 stencil_valid_sched_gen(
		.clk(clk),
		.clk_en(clk_en),
		.cycle_count(cycle_count),
		.enable(stencil_valid_sched_gen_enable),
		.finished(loops_stencil_valid_restart),
		.flush(flush),
		.mux_sel(loops_stencil_valid_mux_sel_out),
		.rst_n(rst_n),
		.sched_addr_gen_starting_addr(stencil_valid_sched_gen_sched_addr_gen_starting_addr),
		.sched_addr_gen_strides_0(stencil_valid_sched_gen_sched_addr_gen_strides_0),
		.sched_addr_gen_strides_1(stencil_valid_sched_gen_sched_addr_gen_strides_1),
		.sched_addr_gen_strides_2(stencil_valid_sched_gen_sched_addr_gen_strides_2),
		.sched_addr_gen_strides_3(stencil_valid_sched_gen_sched_addr_gen_strides_3),
		.sched_addr_gen_strides_4(stencil_valid_sched_gen_sched_addr_gen_strides_4),
		.sched_addr_gen_strides_5(stencil_valid_sched_gen_sched_addr_gen_strides_5),
		.valid_output(stencil_valid_internal)
	);
endmodule
module stencil_valid_flat (
	clk,
	clk_en,
	flush,
	rst_n,
	stencil_valid_inst_loops_stencil_valid_dimensionality,
	stencil_valid_inst_loops_stencil_valid_ranges_0,
	stencil_valid_inst_loops_stencil_valid_ranges_1,
	stencil_valid_inst_loops_stencil_valid_ranges_2,
	stencil_valid_inst_loops_stencil_valid_ranges_3,
	stencil_valid_inst_loops_stencil_valid_ranges_4,
	stencil_valid_inst_loops_stencil_valid_ranges_5,
	stencil_valid_inst_stencil_valid_sched_gen_enable,
	stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr,
	stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0,
	stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1,
	stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2,
	stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3,
	stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4,
	stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5,
	stencil_valid_f_
);
	input wire clk;
	input wire clk_en;
	input wire flush;
	input wire rst_n;
	input wire [3:0] stencil_valid_inst_loops_stencil_valid_dimensionality;
	input wire [10:0] stencil_valid_inst_loops_stencil_valid_ranges_0;
	input wire [10:0] stencil_valid_inst_loops_stencil_valid_ranges_1;
	input wire [10:0] stencil_valid_inst_loops_stencil_valid_ranges_2;
	input wire [10:0] stencil_valid_inst_loops_stencil_valid_ranges_3;
	input wire [10:0] stencil_valid_inst_loops_stencil_valid_ranges_4;
	input wire [10:0] stencil_valid_inst_loops_stencil_valid_ranges_5;
	input wire stencil_valid_inst_stencil_valid_sched_gen_enable;
	input wire [15:0] stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr;
	input wire [15:0] stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0;
	input wire [15:0] stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1;
	input wire [15:0] stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2;
	input wire [15:0] stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3;
	input wire [15:0] stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4;
	input wire [15:0] stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5;
	output wire stencil_valid_f_;
	stencil_valid stencil_valid_inst(
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.loops_stencil_valid_dimensionality(stencil_valid_inst_loops_stencil_valid_dimensionality),
		.loops_stencil_valid_ranges_0(stencil_valid_inst_loops_stencil_valid_ranges_0),
		.loops_stencil_valid_ranges_1(stencil_valid_inst_loops_stencil_valid_ranges_1),
		.loops_stencil_valid_ranges_2(stencil_valid_inst_loops_stencil_valid_ranges_2),
		.loops_stencil_valid_ranges_3(stencil_valid_inst_loops_stencil_valid_ranges_3),
		.loops_stencil_valid_ranges_4(stencil_valid_inst_loops_stencil_valid_ranges_4),
		.loops_stencil_valid_ranges_5(stencil_valid_inst_loops_stencil_valid_ranges_5),
		.rst_n(rst_n),
		.stencil_valid_sched_gen_enable(stencil_valid_inst_stencil_valid_sched_gen_enable),
		.stencil_valid_sched_gen_sched_addr_gen_starting_addr(stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr),
		.stencil_valid_sched_gen_sched_addr_gen_strides_0(stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0),
		.stencil_valid_sched_gen_sched_addr_gen_strides_1(stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1),
		.stencil_valid_sched_gen_sched_addr_gen_strides_2(stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2),
		.stencil_valid_sched_gen_sched_addr_gen_strides_3(stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3),
		.stencil_valid_sched_gen_sched_addr_gen_strides_4(stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4),
		.stencil_valid_sched_gen_sched_addr_gen_strides_5(stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5),
		.stencil_valid(stencil_valid_f_)
	);
endmodule
module storage_config_seq_2_64_16 (
	clk,
	clk_en,
	config_addr_in,
	config_data_in,
	config_en,
	config_rd,
	config_wr,
	flush,
	rd_data_stg,
	rst_n,
	addr_out,
	rd_data_out,
	ren_out,
	wen_out,
	wr_data
);
	input wire clk;
	input wire clk_en;
	input wire [7:0] config_addr_in;
	input wire [15:0] config_data_in;
	input wire [1:0] config_en;
	input wire config_rd;
	input wire config_wr;
	input wire flush;
	input wire [63:0] rd_data_stg;
	input wire rst_n;
	output wire [8:0] addr_out;
	output wire [31:0] rd_data_out;
	output wire ren_out;
	output wire wen_out;
	output wire [63:0] wr_data;
	reg [1:0] cnt;
	reg [47:0] data_wr_reg;
	reg [1:0] rd_cnt;
	reg rd_valid;
	wire [1:0] reduce_en;
	reg set_to_addr;
	assign reduce_en[0] = |config_en[0];
	assign reduce_en[1] = |config_en[1];
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	always @(*) begin
		set_to_addr = 1'h0;
		begin : sv2v_autoblock_1
			reg [31:0] i;
			for (i = 0; i < 2; i = i + 1)
				if (reduce_en[sv2v_cast_1(i)])
					set_to_addr = sv2v_cast_1(i);
		end
	end
	assign addr_out = {set_to_addr, config_addr_in};
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			cnt <= 2'h0;
		else if (flush)
			cnt <= 2'h0;
		else if (config_wr & |config_en)
			cnt <= cnt + 2'h1;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			rd_valid <= 1'h0;
		else if (flush)
			rd_valid <= 1'h0;
		else
			rd_valid <= config_rd & |config_en;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			rd_cnt <= 2'h0;
		else if (flush)
			rd_cnt <= 2'h0;
		else if (rd_valid & ~(config_rd & |config_en))
			rd_cnt <= rd_cnt + 2'h1;
	assign rd_data_out[0+:16] = rd_data_stg[(0 + rd_cnt) * 16+:16];
	assign rd_data_out[16+:16] = rd_data_stg[(0 + rd_cnt) * 16+:16];
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			data_wr_reg <= 48'h000000000000;
		else if (flush)
			data_wr_reg <= 48'h000000000000;
		else if (config_wr & (cnt < 2'h3))
			data_wr_reg[cnt * 16+:16] <= config_data_in;
	assign wr_data[0+:16] = data_wr_reg[0+:16];
	assign wr_data[16+:16] = data_wr_reg[16+:16];
	assign wr_data[32+:16] = data_wr_reg[32+:16];
	assign wr_data[48+:16] = config_data_in;
	assign wen_out = config_wr & (cnt == 2'h3);
	assign ren_out = config_rd;
endmodule
module strg_ram_64_512_delay1 (
	clk,
	clk_en,
	data_from_strg,
	data_in,
	flush,
	rd_addr_in,
	ren,
	rst_n,
	wen,
	wr_addr_in,
	addr_out,
	data_out,
	data_to_strg,
	ready,
	ren_to_strg,
	valid_out,
	wen_to_strg
);
	input wire clk;
	input wire clk_en;
	input wire [63:0] data_from_strg;
	input wire [16:0] data_in;
	input wire flush;
	input wire [16:0] rd_addr_in;
	input wire ren;
	input wire rst_n;
	input wire wen;
	input wire [16:0] wr_addr_in;
	output reg [8:0] addr_out;
	output reg [16:0] data_out;
	output wire [63:0] data_to_strg;
	output reg ready;
	output wire ren_to_strg;
	output reg valid_out;
	output wire wen_to_strg;
	reg [15:0] addr_to_write;
	reg [63:0] data_combined;
	reg [15:0] data_to_write;
	reg [1:0] r_w_seq_current_state;
	reg [1:0] r_w_seq_next_state;
	wire [15:0] rd_addr;
	wire rd_bank;
	reg read_gate;
	wire [15:0] wr_addr;
	reg write_gate;
	assign wr_addr = wr_addr_in[15:0];
	assign rd_addr = wr_addr_in[15:0];
	assign rd_bank = 1'h0;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			data_to_write <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				data_to_write <= 16'h0000;
			else
				data_to_write <= data_in[15:0];
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			addr_to_write <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				addr_to_write <= 16'h0000;
			else
				addr_to_write <= wr_addr;
		end
	assign data_to_strg[0+:64] = data_combined;
	assign ren_to_strg = (wen | ren) & read_gate;
	assign wen_to_strg = write_gate;
	always @(*) begin
		addr_out[0+:9] = rd_addr[10:2];
		if (wen & ~write_gate)
			addr_out[0+:9] = wr_addr[10:2];
		else if (write_gate)
			addr_out[0+:9] = addr_to_write[10:2];
	end
	always @(*)
		if (addr_to_write[1:0] == 2'h0)
			data_combined[0+:16] = data_to_write;
		else
			data_combined[0+:16] = data_from_strg[(rd_bank * 4) * 16+:16];
	always @(*)
		if (addr_to_write[1:0] == 2'h1)
			data_combined[16+:16] = data_to_write;
		else
			data_combined[16+:16] = data_from_strg[((rd_bank * 4) + 1) * 16+:16];
	always @(*)
		if (addr_to_write[1:0] == 2'h2)
			data_combined[32+:16] = data_to_write;
		else
			data_combined[32+:16] = data_from_strg[((rd_bank * 4) + 2) * 16+:16];
	always @(*)
		if (addr_to_write[1:0] == 2'h3)
			data_combined[48+:16] = data_to_write;
		else
			data_combined[48+:16] = data_from_strg[((rd_bank * 4) + 3) * 16+:16];
	always @(posedge clk or negedge rst_n)
		if (!rst_n)
			r_w_seq_current_state <= 2'h0;
		else
			r_w_seq_current_state <= r_w_seq_next_state;
	always @(*) begin
		r_w_seq_next_state = r_w_seq_current_state;
		case (r_w_seq_current_state)
			2'h0:
				if (~wen & ~ren)
					r_w_seq_next_state = 2'h0;
				else if (ren & ~wen)
					r_w_seq_next_state = 2'h2;
				else if (wen)
					r_w_seq_next_state = 2'h1;
			2'h1: r_w_seq_next_state = 2'h0;
			2'h2:
				if (~wen & ~ren)
					r_w_seq_next_state = 2'h0;
				else if (ren & ~wen)
					r_w_seq_next_state = 2'h2;
				else if (wen)
					r_w_seq_next_state = 2'h1;
			2'h3: r_w_seq_next_state = 2'h3;
			default:
				;
		endcase
	end
	always @(*)
		case (r_w_seq_current_state)
			2'h0: begin : r_w_seq_IDLE_Output
				ready = 1'h1;
				valid_out = 1'h0;
				data_out[15:0] = 16'h0000;
				data_out[16] = 1'h0;
				write_gate = 1'h0;
				read_gate = 1'h1;
			end
			2'h1: begin : r_w_seq_MODIFY_Output
				ready = 1'h0;
				valid_out = 1'h0;
				data_out[15:0] = 16'h0000;
				data_out[16] = 1'h0;
				write_gate = 1'h1;
				read_gate = 1'h0;
			end
			2'h2: begin : r_w_seq_READ_Output
				ready = 1'h1;
				valid_out = 1'h1;
				data_out[15:0] = data_from_strg[((rd_bank * 4) + addr_to_write[1:0]) * 16+:16];
				data_out[16] = 1'h0;
				write_gate = 1'h0;
				read_gate = 1'h1;
			end
			2'h3: begin : r_w_seq__DEFAULT_Output
				ready = 1'h0;
				valid_out = 1'h0;
				data_out[15:0] = 16'h0000;
				data_out[16] = 1'h0;
				write_gate = 1'h0;
				read_gate = 1'h0;
			end
			default:
				;
		endcase
endmodule
module strg_ram_64_512_delay1_flat (
	clk,
	clk_en,
	data_in_f_,
	flush,
	rd_addr_in_f_,
	ren_f_,
	rst_n,
	strg_ram_64_512_delay1_inst_data_from_strg_lifted,
	wen_f_,
	wr_addr_in_f_,
	data_out_f_,
	ready_f_,
	strg_ram_64_512_delay1_inst_addr_out_lifted,
	strg_ram_64_512_delay1_inst_data_to_strg_lifted,
	strg_ram_64_512_delay1_inst_ren_to_strg_lifted,
	strg_ram_64_512_delay1_inst_wen_to_strg_lifted,
	valid_out_f_
);
	input wire clk;
	input wire clk_en;
	input wire [16:0] data_in_f_;
	input wire flush;
	input wire [16:0] rd_addr_in_f_;
	input wire ren_f_;
	input wire rst_n;
	input wire [63:0] strg_ram_64_512_delay1_inst_data_from_strg_lifted;
	input wire wen_f_;
	input wire [16:0] wr_addr_in_f_;
	output wire [16:0] data_out_f_;
	output wire ready_f_;
	output wire [8:0] strg_ram_64_512_delay1_inst_addr_out_lifted;
	output wire [63:0] strg_ram_64_512_delay1_inst_data_to_strg_lifted;
	output wire strg_ram_64_512_delay1_inst_ren_to_strg_lifted;
	output wire strg_ram_64_512_delay1_inst_wen_to_strg_lifted;
	output wire valid_out_f_;
	strg_ram_64_512_delay1 strg_ram_64_512_delay1_inst(
		.clk(clk),
		.clk_en(clk_en),
		.data_from_strg(strg_ram_64_512_delay1_inst_data_from_strg_lifted),
		.data_in(data_in_f_),
		.flush(flush),
		.rd_addr_in(rd_addr_in_f_),
		.ren(ren_f_),
		.rst_n(rst_n),
		.wen(wen_f_),
		.wr_addr_in(wr_addr_in_f_),
		.addr_out(strg_ram_64_512_delay1_inst_addr_out_lifted),
		.data_out(data_out_f_),
		.data_to_strg(strg_ram_64_512_delay1_inst_data_to_strg_lifted),
		.ready(ready_f_),
		.ren_to_strg(strg_ram_64_512_delay1_inst_ren_to_strg_lifted),
		.valid_out(valid_out_f_),
		.wen_to_strg(strg_ram_64_512_delay1_inst_wen_to_strg_lifted)
	);
endmodule
module strg_ub_agg_only (
	agg_read,
	agg_write_addr_gen_0_starting_addr,
	agg_write_addr_gen_0_strides_0,
	agg_write_addr_gen_0_strides_1,
	agg_write_addr_gen_0_strides_2,
	agg_write_addr_gen_1_starting_addr,
	agg_write_addr_gen_1_strides_0,
	agg_write_addr_gen_1_strides_1,
	agg_write_addr_gen_1_strides_2,
	agg_write_sched_gen_0_enable,
	agg_write_sched_gen_0_sched_addr_gen_starting_addr,
	agg_write_sched_gen_0_sched_addr_gen_strides_0,
	agg_write_sched_gen_0_sched_addr_gen_strides_1,
	agg_write_sched_gen_0_sched_addr_gen_strides_2,
	agg_write_sched_gen_1_enable,
	agg_write_sched_gen_1_sched_addr_gen_starting_addr,
	agg_write_sched_gen_1_sched_addr_gen_strides_0,
	agg_write_sched_gen_1_sched_addr_gen_strides_1,
	agg_write_sched_gen_1_sched_addr_gen_strides_2,
	clk,
	clk_en,
	cycle_count,
	data_in,
	flush,
	loops_in2buf_0_dimensionality,
	loops_in2buf_0_ranges_0,
	loops_in2buf_0_ranges_1,
	loops_in2buf_0_ranges_2,
	loops_in2buf_1_dimensionality,
	loops_in2buf_1_ranges_0,
	loops_in2buf_1_ranges_1,
	loops_in2buf_1_ranges_2,
	rst_n,
	sram_read_addr_in,
	tb_read_addr_d_in,
	tb_read_d_in,
	update_mode_in,
	agg_data_out,
	agg_write_addr_l2b_out,
	agg_write_mux_sel_out,
	agg_write_out,
	agg_write_restart_out
);
	input wire [1:0] agg_read;
	input wire [2:0] agg_write_addr_gen_0_starting_addr;
	input wire [2:0] agg_write_addr_gen_0_strides_0;
	input wire [2:0] agg_write_addr_gen_0_strides_1;
	input wire [2:0] agg_write_addr_gen_0_strides_2;
	input wire [2:0] agg_write_addr_gen_1_starting_addr;
	input wire [2:0] agg_write_addr_gen_1_strides_0;
	input wire [2:0] agg_write_addr_gen_1_strides_1;
	input wire [2:0] agg_write_addr_gen_1_strides_2;
	input wire agg_write_sched_gen_0_enable;
	input wire [15:0] agg_write_sched_gen_0_sched_addr_gen_starting_addr;
	input wire [15:0] agg_write_sched_gen_0_sched_addr_gen_strides_0;
	input wire [15:0] agg_write_sched_gen_0_sched_addr_gen_strides_1;
	input wire [15:0] agg_write_sched_gen_0_sched_addr_gen_strides_2;
	input wire agg_write_sched_gen_1_enable;
	input wire [15:0] agg_write_sched_gen_1_sched_addr_gen_starting_addr;
	input wire [15:0] agg_write_sched_gen_1_sched_addr_gen_strides_0;
	input wire [15:0] agg_write_sched_gen_1_sched_addr_gen_strides_1;
	input wire [15:0] agg_write_sched_gen_1_sched_addr_gen_strides_2;
	input wire clk;
	input wire clk_en;
	input wire [15:0] cycle_count;
	input wire [31:0] data_in;
	input wire flush;
	input wire [2:0] loops_in2buf_0_dimensionality;
	input wire [10:0] loops_in2buf_0_ranges_0;
	input wire [10:0] loops_in2buf_0_ranges_1;
	input wire [10:0] loops_in2buf_0_ranges_2;
	input wire [2:0] loops_in2buf_1_dimensionality;
	input wire [10:0] loops_in2buf_1_ranges_0;
	input wire [10:0] loops_in2buf_1_ranges_1;
	input wire [10:0] loops_in2buf_1_ranges_2;
	input wire rst_n;
	input wire [17:0] sram_read_addr_in;
	input wire [5:0] tb_read_addr_d_in;
	input wire [1:0] tb_read_d_in;
	input wire [3:0] update_mode_in;
	output reg [127:0] agg_data_out;
	output wire [3:0] agg_write_addr_l2b_out;
	output wire [5:0] agg_write_mux_sel_out;
	output wire [1:0] agg_write_out;
	output wire [1:0] agg_write_restart_out;
	reg [255:0] agg;
	wire [1:0] agg_read_addr;
	wire [15:0] agg_read_addr_gen_out;
	wire [1:0] agg_read_addr_in;
	wire [1:0] agg_write;
	wire [5:0] agg_write_addr;
	wire [2:0] agg_write_addr_gen_0_addr_out;
	wire [8:0] agg_write_addr_gen_0_strides;
	wire [2:0] agg_write_addr_gen_1_addr_out;
	wire [8:0] agg_write_addr_gen_1_strides;
	wire agg_write_sched_gen_0_valid_output;
	wire agg_write_sched_gen_1_valid_output;
	wire [2:0] fl_mux_sel_0;
	wire [2:0] fl_mux_sel_1;
	wire [1:0] loops_in2buf_0_mux_sel_out;
	wire [32:0] loops_in2buf_0_ranges;
	wire loops_in2buf_0_restart;
	wire [1:0] loops_in2buf_1_mux_sel_out;
	wire [32:0] loops_in2buf_1_ranges;
	wire loops_in2buf_1_restart;
	wire [1:0] mode_0;
	wire [1:0] mode_1;
	wire [2:0] tb_addr_0;
	wire [2:0] tb_addr_1;
	wire tb_read_0;
	wire tb_read_1;
	assign agg_write_out = agg_write;
	assign mode_0 = update_mode_in[0+:2];
	assign agg_write_addr_l2b_out[0+:2] = agg_write_addr[1-:2];
	assign tb_read_0 = (mode_0[0] ? tb_read_d_in[1] : tb_read_d_in[0]);
	assign tb_addr_0 = (mode_0[0] ? tb_read_addr_d_in[3+:3] : tb_read_addr_d_in[0+:3]);
	assign fl_mux_sel_0[1:0] = loops_in2buf_0_mux_sel_out;
	assign fl_mux_sel_0[2] = 1'h0;
	assign agg_write_mux_sel_out[0+:3] = fl_mux_sel_0;
	assign agg_write_restart_out[0] = loops_in2buf_0_restart;
	assign agg_write_addr[0+:3] = (mode_0[1] ? tb_addr_0 : agg_write_addr_gen_0_addr_out);
	assign agg_write[0] = (mode_0[1] ? tb_read_0 : agg_write_sched_gen_0_valid_output);
	always @(posedge clk)
		if (clk_en) begin
			if (agg_write[0])
				agg[(((0 + agg_write_addr[2]) * 4) + agg_write_addr[1-:2]) * 16+:16] <= data_in[0+:16];
		end
	assign agg_read_addr_in[0] = sram_read_addr_in[0];
	assign agg_read_addr_gen_out[0] = agg_read_addr_in[0];
	assign agg_read_addr_gen_out[7-:7] = 7'h00;
	assign agg_read_addr[0] = agg_read_addr_gen_out[0];
	always @(*) agg_data_out[0+:64] = agg[16 * ((0 + agg_read_addr[0]) * 4)+:64];
	assign mode_1 = update_mode_in[2+:2];
	assign agg_write_addr_l2b_out[2+:2] = agg_write_addr[4-:2];
	assign tb_read_1 = (mode_1[0] ? tb_read_d_in[1] : tb_read_d_in[0]);
	assign tb_addr_1 = (mode_1[0] ? tb_read_addr_d_in[3+:3] : tb_read_addr_d_in[0+:3]);
	assign fl_mux_sel_1[1:0] = loops_in2buf_1_mux_sel_out;
	assign fl_mux_sel_1[2] = 1'h0;
	assign agg_write_mux_sel_out[3+:3] = fl_mux_sel_1;
	assign agg_write_restart_out[1] = loops_in2buf_1_restart;
	assign agg_write_addr[3+:3] = (mode_1[1] ? tb_addr_1 : agg_write_addr_gen_1_addr_out);
	assign agg_write[1] = (mode_1[1] ? tb_read_1 : agg_write_sched_gen_1_valid_output);
	always @(posedge clk)
		if (clk_en) begin
			if (agg_write[1])
				agg[(((2 + agg_write_addr[5]) * 4) + agg_write_addr[4-:2]) * 16+:16] <= data_in[16+:16];
		end
	assign agg_read_addr_in[1] = sram_read_addr_in[9];
	assign agg_read_addr_gen_out[8] = agg_read_addr_in[1];
	assign agg_read_addr_gen_out[15-:7] = 7'h00;
	assign agg_read_addr[1] = agg_read_addr_gen_out[8];
	always @(*) agg_data_out[64+:64] = agg[16 * ((2 + agg_read_addr[1]) * 4)+:64];
	assign loops_in2buf_0_ranges[0+:11] = loops_in2buf_0_ranges_0;
	assign loops_in2buf_0_ranges[11+:11] = loops_in2buf_0_ranges_1;
	assign loops_in2buf_0_ranges[22+:11] = loops_in2buf_0_ranges_2;
	assign agg_write_addr_gen_0_strides[0+:3] = agg_write_addr_gen_0_strides_0;
	assign agg_write_addr_gen_0_strides[3+:3] = agg_write_addr_gen_0_strides_1;
	assign agg_write_addr_gen_0_strides[6+:3] = agg_write_addr_gen_0_strides_2;
	assign loops_in2buf_1_ranges[0+:11] = loops_in2buf_1_ranges_0;
	assign loops_in2buf_1_ranges[11+:11] = loops_in2buf_1_ranges_1;
	assign loops_in2buf_1_ranges[22+:11] = loops_in2buf_1_ranges_2;
	assign agg_write_addr_gen_1_strides[0+:3] = agg_write_addr_gen_1_strides_0;
	assign agg_write_addr_gen_1_strides[3+:3] = agg_write_addr_gen_1_strides_1;
	assign agg_write_addr_gen_1_strides[6+:3] = agg_write_addr_gen_1_strides_2;
	for_loop_3_11 loops_in2buf_0(
		.clk(clk),
		.clk_en(clk_en),
		.dimensionality(loops_in2buf_0_dimensionality),
		.flush(flush),
		.ranges(loops_in2buf_0_ranges),
		.rst_n(rst_n),
		.step(agg_write[0]),
		.mux_sel_out(loops_in2buf_0_mux_sel_out),
		.restart(loops_in2buf_0_restart)
	);
	addr_gen_3_3 agg_write_addr_gen_0(
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.mux_sel(loops_in2buf_0_mux_sel_out),
		.restart(loops_in2buf_0_restart),
		.rst_n(rst_n),
		.starting_addr(agg_write_addr_gen_0_starting_addr),
		.step(agg_write[0]),
		.strides(agg_write_addr_gen_0_strides),
		.addr_out(agg_write_addr_gen_0_addr_out)
	);
	sched_gen_3_16 agg_write_sched_gen_0(
		.clk(clk),
		.clk_en(clk_en),
		.cycle_count(cycle_count),
		.enable(agg_write_sched_gen_0_enable),
		.finished(loops_in2buf_0_restart),
		.flush(flush),
		.mux_sel(loops_in2buf_0_mux_sel_out),
		.rst_n(rst_n),
		.sched_addr_gen_starting_addr(agg_write_sched_gen_0_sched_addr_gen_starting_addr),
		.sched_addr_gen_strides_0(agg_write_sched_gen_0_sched_addr_gen_strides_0),
		.sched_addr_gen_strides_1(agg_write_sched_gen_0_sched_addr_gen_strides_1),
		.sched_addr_gen_strides_2(agg_write_sched_gen_0_sched_addr_gen_strides_2),
		.valid_output(agg_write_sched_gen_0_valid_output)
	);
	for_loop_3_11 loops_in2buf_1(
		.clk(clk),
		.clk_en(clk_en),
		.dimensionality(loops_in2buf_1_dimensionality),
		.flush(flush),
		.ranges(loops_in2buf_1_ranges),
		.rst_n(rst_n),
		.step(agg_write[1]),
		.mux_sel_out(loops_in2buf_1_mux_sel_out),
		.restart(loops_in2buf_1_restart)
	);
	addr_gen_3_3 agg_write_addr_gen_1(
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.mux_sel(loops_in2buf_1_mux_sel_out),
		.restart(loops_in2buf_1_restart),
		.rst_n(rst_n),
		.starting_addr(agg_write_addr_gen_1_starting_addr),
		.step(agg_write[1]),
		.strides(agg_write_addr_gen_1_strides),
		.addr_out(agg_write_addr_gen_1_addr_out)
	);
	sched_gen_3_16 agg_write_sched_gen_1(
		.clk(clk),
		.clk_en(clk_en),
		.cycle_count(cycle_count),
		.enable(agg_write_sched_gen_1_enable),
		.finished(loops_in2buf_1_restart),
		.flush(flush),
		.mux_sel(loops_in2buf_1_mux_sel_out),
		.rst_n(rst_n),
		.sched_addr_gen_starting_addr(agg_write_sched_gen_1_sched_addr_gen_starting_addr),
		.sched_addr_gen_strides_0(agg_write_sched_gen_1_sched_addr_gen_strides_0),
		.sched_addr_gen_strides_1(agg_write_sched_gen_1_sched_addr_gen_strides_1),
		.sched_addr_gen_strides_2(agg_write_sched_gen_1_sched_addr_gen_strides_2),
		.valid_output(agg_write_sched_gen_1_valid_output)
	);
endmodule
module strg_ub_agg_sram_shared (
	agg_read_sched_gen_0_agg_read_padding,
	agg_read_sched_gen_1_agg_read_padding,
	agg_sram_shared_addr_gen_0_starting_addr,
	agg_sram_shared_addr_gen_1_starting_addr,
	agg_write_addr_l2b_in,
	agg_write_in,
	agg_write_mux_sel_in,
	agg_write_restart_in,
	clk,
	clk_en,
	flush,
	mode_0,
	mode_1,
	rst_n,
	sram_read_addr_in,
	sram_read_d_in,
	sram_read_in,
	agg_read_out,
	agg_sram_shared_addr_out,
	update_mode_out
);
	input wire [7:0] agg_read_sched_gen_0_agg_read_padding;
	input wire [7:0] agg_read_sched_gen_1_agg_read_padding;
	input wire [8:0] agg_sram_shared_addr_gen_0_starting_addr;
	input wire [8:0] agg_sram_shared_addr_gen_1_starting_addr;
	input wire [3:0] agg_write_addr_l2b_in;
	input wire [1:0] agg_write_in;
	input wire [5:0] agg_write_mux_sel_in;
	input wire [1:0] agg_write_restart_in;
	input wire clk;
	input wire clk_en;
	input wire flush;
	input wire [1:0] mode_0;
	input wire [1:0] mode_1;
	input wire rst_n;
	input wire [17:0] sram_read_addr_in;
	input wire [1:0] sram_read_d_in;
	input wire [1:0] sram_read_in;
	output wire [1:0] agg_read_out;
	output wire [17:0] agg_sram_shared_addr_out;
	output wire [3:0] update_mode_out;
	wire [1:0] agg_read;
	wire agg_read_sched_gen_0_valid_output;
	wire agg_read_sched_gen_1_valid_output;
	wire [8:0] agg_sram_shared_addr_gen_0_addr_out;
	wire [8:0] agg_sram_shared_addr_gen_1_addr_out;
	assign agg_read_out = agg_read;
	assign update_mode_out[0+:2] = mode_0;
	assign agg_read[0] = agg_read_sched_gen_0_valid_output;
	assign agg_sram_shared_addr_out[0+:9] = agg_sram_shared_addr_gen_0_addr_out;
	assign update_mode_out[2+:2] = mode_1;
	assign agg_read[1] = agg_read_sched_gen_1_valid_output;
	assign agg_sram_shared_addr_out[9+:9] = agg_sram_shared_addr_gen_1_addr_out;
	agg_sram_shared_sched_gen agg_read_sched_gen_0(
		.agg_read_padding(agg_read_sched_gen_0_agg_read_padding),
		.agg_write(agg_write_in[0]),
		.agg_write_addr_l2b(agg_write_addr_l2b_in[0+:2]),
		.agg_write_mux_sel(agg_write_mux_sel_in[0+:3]),
		.agg_write_restart(agg_write_restart_in[0]),
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.mode(mode_0),
		.rst_n(rst_n),
		.sram_read_d(sram_read_d_in),
		.valid_output(agg_read_sched_gen_0_valid_output)
	);
	agg_sram_shared_addr_gen agg_sram_shared_addr_gen_0(
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.mode(mode_0),
		.rst_n(rst_n),
		.sram_read(sram_read_in),
		.sram_read_addr(sram_read_addr_in),
		.starting_addr(agg_sram_shared_addr_gen_0_starting_addr),
		.step(agg_read[0]),
		.addr_out(agg_sram_shared_addr_gen_0_addr_out)
	);
	agg_sram_shared_sched_gen agg_read_sched_gen_1(
		.agg_read_padding(agg_read_sched_gen_1_agg_read_padding),
		.agg_write(agg_write_in[1]),
		.agg_write_addr_l2b(agg_write_addr_l2b_in[2+:2]),
		.agg_write_mux_sel(agg_write_mux_sel_in[3+:3]),
		.agg_write_restart(agg_write_restart_in[1]),
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.mode(mode_1),
		.rst_n(rst_n),
		.sram_read_d(sram_read_d_in),
		.valid_output(agg_read_sched_gen_1_valid_output)
	);
	agg_sram_shared_addr_gen agg_sram_shared_addr_gen_1(
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.mode(mode_1),
		.rst_n(rst_n),
		.sram_read(sram_read_in),
		.sram_read_addr(sram_read_addr_in),
		.starting_addr(agg_sram_shared_addr_gen_1_starting_addr),
		.step(agg_read[1]),
		.addr_out(agg_sram_shared_addr_gen_1_addr_out)
	);
endmodule
module strg_ub_sram_only (
	agg_data_out,
	agg_read,
	clk,
	clk_en,
	cycle_count,
	flush,
	loops_sram2tb_mux_sel,
	loops_sram2tb_restart,
	output_addr_gen_0_starting_addr,
	output_addr_gen_0_strides_0,
	output_addr_gen_0_strides_1,
	output_addr_gen_0_strides_2,
	output_addr_gen_0_strides_3,
	output_addr_gen_0_strides_4,
	output_addr_gen_0_strides_5,
	output_addr_gen_1_starting_addr,
	output_addr_gen_1_strides_0,
	output_addr_gen_1_strides_1,
	output_addr_gen_1_strides_2,
	output_addr_gen_1_strides_3,
	output_addr_gen_1_strides_4,
	output_addr_gen_1_strides_5,
	rst_n,
	sram_read_addr_in,
	t_read,
	addr_to_sram,
	cen_to_sram,
	data_to_sram,
	sram_read_addr_out,
	wen_to_sram
);
	input wire [127:0] agg_data_out;
	input wire [1:0] agg_read;
	input wire clk;
	input wire clk_en;
	input wire [15:0] cycle_count;
	input wire flush;
	input wire [5:0] loops_sram2tb_mux_sel;
	input wire [1:0] loops_sram2tb_restart;
	input wire [8:0] output_addr_gen_0_starting_addr;
	input wire [8:0] output_addr_gen_0_strides_0;
	input wire [8:0] output_addr_gen_0_strides_1;
	input wire [8:0] output_addr_gen_0_strides_2;
	input wire [8:0] output_addr_gen_0_strides_3;
	input wire [8:0] output_addr_gen_0_strides_4;
	input wire [8:0] output_addr_gen_0_strides_5;
	input wire [8:0] output_addr_gen_1_starting_addr;
	input wire [8:0] output_addr_gen_1_strides_0;
	input wire [8:0] output_addr_gen_1_strides_1;
	input wire [8:0] output_addr_gen_1_strides_2;
	input wire [8:0] output_addr_gen_1_strides_3;
	input wire [8:0] output_addr_gen_1_strides_4;
	input wire [8:0] output_addr_gen_1_strides_5;
	input wire rst_n;
	input wire [17:0] sram_read_addr_in;
	input wire [1:0] t_read;
	output wire [8:0] addr_to_sram;
	output wire cen_to_sram;
	output wire [63:0] data_to_sram;
	output wire [17:0] sram_read_addr_out;
	output wire wen_to_sram;
	reg [8:0] addr;
	reg [63:0] decode_ret_agg_read_agg_data_out;
	reg [15:0] decode_ret_agg_read_s_write_addr;
	reg [15:0] decode_ret_t_read_s_read_addr;
	reg decode_sel_done_agg_read_agg_data_out;
	reg decode_sel_done_agg_read_s_write_addr;
	reg decode_sel_done_t_read_s_read_addr;
	wire [8:0] output_addr_gen_0_addr_out;
	wire [53:0] output_addr_gen_0_strides;
	wire [8:0] output_addr_gen_1_addr_out;
	wire [53:0] output_addr_gen_1_strides;
	wire read;
	wire [31:0] s_read_addr;
	wire [31:0] s_write_addr;
	wire [63:0] sram_write_data;
	wire write;
	assign s_write_addr[8-:9] = sram_read_addr_in[0+:9];
	assign s_write_addr[15-:7] = 7'h00;
	assign s_write_addr[24-:9] = sram_read_addr_in[9+:9];
	assign s_write_addr[31-:7] = 7'h00;
	assign s_read_addr[8-:9] = output_addr_gen_0_addr_out;
	assign s_read_addr[15-:7] = 7'h00;
	assign sram_read_addr_out[0+:9] = output_addr_gen_0_addr_out;
	assign s_read_addr[24-:9] = output_addr_gen_1_addr_out;
	assign s_read_addr[31-:7] = 7'h00;
	assign sram_read_addr_out[9+:9] = output_addr_gen_1_addr_out;
	assign data_to_sram = sram_write_data;
	assign wen_to_sram = write;
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	always @(*) begin
		decode_sel_done_agg_read_s_write_addr = 1'h0;
		decode_ret_agg_read_s_write_addr = 16'h0000;
		begin : sv2v_autoblock_1
			reg [31:0] i;
			for (i = 0; i < 2; i = i + 1)
				if (~decode_sel_done_agg_read_s_write_addr & agg_read[sv2v_cast_1(i)]) begin
					decode_ret_agg_read_s_write_addr = s_write_addr[sv2v_cast_1(i) * 16+:16];
					decode_sel_done_agg_read_s_write_addr = 1'h1;
				end
		end
	end
	always @(*) begin
		decode_sel_done_t_read_s_read_addr = 1'h0;
		decode_ret_t_read_s_read_addr = 16'h0000;
		begin : sv2v_autoblock_2
			reg [31:0] i;
			for (i = 0; i < 2; i = i + 1)
				if (~decode_sel_done_t_read_s_read_addr & t_read[sv2v_cast_1(i)]) begin
					decode_ret_t_read_s_read_addr = s_read_addr[sv2v_cast_1(i) * 16+:16];
					decode_sel_done_t_read_s_read_addr = 1'h1;
				end
		end
	end
	assign cen_to_sram = write | read;
	assign addr_to_sram = addr;
	always @(*)
		if (write)
			addr = decode_ret_agg_read_s_write_addr[8:0];
		else
			addr = decode_ret_t_read_s_read_addr[8:0];
	assign write = |agg_read;
	assign read = |t_read;
	always @(*) begin
		decode_sel_done_agg_read_agg_data_out = 1'h0;
		decode_ret_agg_read_agg_data_out = 64'h0000000000000000;
		begin : sv2v_autoblock_3
			reg [31:0] i;
			for (i = 0; i < 2; i = i + 1)
				if (~decode_sel_done_agg_read_agg_data_out & agg_read[sv2v_cast_1(i)]) begin
					decode_ret_agg_read_agg_data_out = agg_data_out[16 * (sv2v_cast_1(i) * 4)+:64];
					decode_sel_done_agg_read_agg_data_out = 1'h1;
				end
		end
	end
	assign sram_write_data = decode_ret_agg_read_agg_data_out;
	assign output_addr_gen_0_strides[0+:9] = output_addr_gen_0_strides_0;
	assign output_addr_gen_0_strides[9+:9] = output_addr_gen_0_strides_1;
	assign output_addr_gen_0_strides[18+:9] = output_addr_gen_0_strides_2;
	assign output_addr_gen_0_strides[27+:9] = output_addr_gen_0_strides_3;
	assign output_addr_gen_0_strides[36+:9] = output_addr_gen_0_strides_4;
	assign output_addr_gen_0_strides[45+:9] = output_addr_gen_0_strides_5;
	assign output_addr_gen_1_strides[0+:9] = output_addr_gen_1_strides_0;
	assign output_addr_gen_1_strides[9+:9] = output_addr_gen_1_strides_1;
	assign output_addr_gen_1_strides[18+:9] = output_addr_gen_1_strides_2;
	assign output_addr_gen_1_strides[27+:9] = output_addr_gen_1_strides_3;
	assign output_addr_gen_1_strides[36+:9] = output_addr_gen_1_strides_4;
	assign output_addr_gen_1_strides[45+:9] = output_addr_gen_1_strides_5;
	addr_gen_6_9 output_addr_gen_0(
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.mux_sel(loops_sram2tb_mux_sel[0+:3]),
		.restart(loops_sram2tb_restart[0]),
		.rst_n(rst_n),
		.starting_addr(output_addr_gen_0_starting_addr),
		.step(t_read[0]),
		.strides(output_addr_gen_0_strides),
		.addr_out(output_addr_gen_0_addr_out)
	);
	addr_gen_6_9 output_addr_gen_1(
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.mux_sel(loops_sram2tb_mux_sel[3+:3]),
		.restart(loops_sram2tb_restart[1]),
		.rst_n(rst_n),
		.starting_addr(output_addr_gen_1_starting_addr),
		.step(t_read[1]),
		.strides(output_addr_gen_1_strides),
		.addr_out(output_addr_gen_1_addr_out)
	);
endmodule
module strg_ub_sram_tb_shared (
	clk,
	clk_en,
	cycle_count,
	flush,
	loops_buf2out_autovec_read_0_dimensionality,
	loops_buf2out_autovec_read_0_ranges_0,
	loops_buf2out_autovec_read_0_ranges_1,
	loops_buf2out_autovec_read_0_ranges_2,
	loops_buf2out_autovec_read_0_ranges_3,
	loops_buf2out_autovec_read_0_ranges_4,
	loops_buf2out_autovec_read_0_ranges_5,
	loops_buf2out_autovec_read_1_dimensionality,
	loops_buf2out_autovec_read_1_ranges_0,
	loops_buf2out_autovec_read_1_ranges_1,
	loops_buf2out_autovec_read_1_ranges_2,
	loops_buf2out_autovec_read_1_ranges_3,
	loops_buf2out_autovec_read_1_ranges_4,
	loops_buf2out_autovec_read_1_ranges_5,
	output_sched_gen_0_enable,
	output_sched_gen_0_sched_addr_gen_delay,
	output_sched_gen_0_sched_addr_gen_starting_addr,
	output_sched_gen_0_sched_addr_gen_strides_0,
	output_sched_gen_0_sched_addr_gen_strides_1,
	output_sched_gen_0_sched_addr_gen_strides_2,
	output_sched_gen_0_sched_addr_gen_strides_3,
	output_sched_gen_0_sched_addr_gen_strides_4,
	output_sched_gen_0_sched_addr_gen_strides_5,
	output_sched_gen_1_enable,
	output_sched_gen_1_sched_addr_gen_delay,
	output_sched_gen_1_sched_addr_gen_starting_addr,
	output_sched_gen_1_sched_addr_gen_strides_0,
	output_sched_gen_1_sched_addr_gen_strides_1,
	output_sched_gen_1_sched_addr_gen_strides_2,
	output_sched_gen_1_sched_addr_gen_strides_3,
	output_sched_gen_1_sched_addr_gen_strides_4,
	output_sched_gen_1_sched_addr_gen_strides_5,
	rst_n,
	loops_sram2tb_mux_sel,
	loops_sram2tb_restart,
	sram_read_d,
	t_read_out
);
	input wire clk;
	input wire clk_en;
	input wire [15:0] cycle_count;
	input wire flush;
	input wire [3:0] loops_buf2out_autovec_read_0_dimensionality;
	input wire [10:0] loops_buf2out_autovec_read_0_ranges_0;
	input wire [10:0] loops_buf2out_autovec_read_0_ranges_1;
	input wire [10:0] loops_buf2out_autovec_read_0_ranges_2;
	input wire [10:0] loops_buf2out_autovec_read_0_ranges_3;
	input wire [10:0] loops_buf2out_autovec_read_0_ranges_4;
	input wire [10:0] loops_buf2out_autovec_read_0_ranges_5;
	input wire [3:0] loops_buf2out_autovec_read_1_dimensionality;
	input wire [10:0] loops_buf2out_autovec_read_1_ranges_0;
	input wire [10:0] loops_buf2out_autovec_read_1_ranges_1;
	input wire [10:0] loops_buf2out_autovec_read_1_ranges_2;
	input wire [10:0] loops_buf2out_autovec_read_1_ranges_3;
	input wire [10:0] loops_buf2out_autovec_read_1_ranges_4;
	input wire [10:0] loops_buf2out_autovec_read_1_ranges_5;
	input wire output_sched_gen_0_enable;
	input wire [9:0] output_sched_gen_0_sched_addr_gen_delay;
	input wire [15:0] output_sched_gen_0_sched_addr_gen_starting_addr;
	input wire [15:0] output_sched_gen_0_sched_addr_gen_strides_0;
	input wire [15:0] output_sched_gen_0_sched_addr_gen_strides_1;
	input wire [15:0] output_sched_gen_0_sched_addr_gen_strides_2;
	input wire [15:0] output_sched_gen_0_sched_addr_gen_strides_3;
	input wire [15:0] output_sched_gen_0_sched_addr_gen_strides_4;
	input wire [15:0] output_sched_gen_0_sched_addr_gen_strides_5;
	input wire output_sched_gen_1_enable;
	input wire [9:0] output_sched_gen_1_sched_addr_gen_delay;
	input wire [15:0] output_sched_gen_1_sched_addr_gen_starting_addr;
	input wire [15:0] output_sched_gen_1_sched_addr_gen_strides_0;
	input wire [15:0] output_sched_gen_1_sched_addr_gen_strides_1;
	input wire [15:0] output_sched_gen_1_sched_addr_gen_strides_2;
	input wire [15:0] output_sched_gen_1_sched_addr_gen_strides_3;
	input wire [15:0] output_sched_gen_1_sched_addr_gen_strides_4;
	input wire [15:0] output_sched_gen_1_sched_addr_gen_strides_5;
	input wire rst_n;
	output wire [5:0] loops_sram2tb_mux_sel;
	output wire [1:0] loops_sram2tb_restart;
	output wire [1:0] sram_read_d;
	output wire [1:0] t_read_out;
	wire [2:0] loops_buf2out_autovec_read_0_mux_sel_out;
	wire [65:0] loops_buf2out_autovec_read_0_ranges;
	wire loops_buf2out_autovec_read_0_restart;
	wire [2:0] loops_buf2out_autovec_read_1_mux_sel_out;
	wire [65:0] loops_buf2out_autovec_read_1_ranges;
	wire loops_buf2out_autovec_read_1_restart;
	wire output_sched_gen_0_valid_output;
	wire output_sched_gen_0_valid_output_d;
	wire output_sched_gen_1_valid_output;
	wire output_sched_gen_1_valid_output_d;
	wire [1:0] t_read;
	assign t_read_out = t_read;
	assign loops_sram2tb_mux_sel[0+:3] = loops_buf2out_autovec_read_0_mux_sel_out;
	assign loops_sram2tb_restart[0] = loops_buf2out_autovec_read_0_restart;
	assign t_read[0] = output_sched_gen_0_valid_output;
	assign sram_read_d[0] = output_sched_gen_0_valid_output_d;
	assign loops_sram2tb_mux_sel[3+:3] = loops_buf2out_autovec_read_1_mux_sel_out;
	assign loops_sram2tb_restart[1] = loops_buf2out_autovec_read_1_restart;
	assign t_read[1] = output_sched_gen_1_valid_output;
	assign sram_read_d[1] = output_sched_gen_1_valid_output_d;
	assign loops_buf2out_autovec_read_0_ranges[0+:11] = loops_buf2out_autovec_read_0_ranges_0;
	assign loops_buf2out_autovec_read_0_ranges[11+:11] = loops_buf2out_autovec_read_0_ranges_1;
	assign loops_buf2out_autovec_read_0_ranges[22+:11] = loops_buf2out_autovec_read_0_ranges_2;
	assign loops_buf2out_autovec_read_0_ranges[33+:11] = loops_buf2out_autovec_read_0_ranges_3;
	assign loops_buf2out_autovec_read_0_ranges[44+:11] = loops_buf2out_autovec_read_0_ranges_4;
	assign loops_buf2out_autovec_read_0_ranges[55+:11] = loops_buf2out_autovec_read_0_ranges_5;
	assign loops_buf2out_autovec_read_1_ranges[0+:11] = loops_buf2out_autovec_read_1_ranges_0;
	assign loops_buf2out_autovec_read_1_ranges[11+:11] = loops_buf2out_autovec_read_1_ranges_1;
	assign loops_buf2out_autovec_read_1_ranges[22+:11] = loops_buf2out_autovec_read_1_ranges_2;
	assign loops_buf2out_autovec_read_1_ranges[33+:11] = loops_buf2out_autovec_read_1_ranges_3;
	assign loops_buf2out_autovec_read_1_ranges[44+:11] = loops_buf2out_autovec_read_1_ranges_4;
	assign loops_buf2out_autovec_read_1_ranges[55+:11] = loops_buf2out_autovec_read_1_ranges_5;
	for_loop_6_11 loops_buf2out_autovec_read_0(
		.clk(clk),
		.clk_en(clk_en),
		.dimensionality(loops_buf2out_autovec_read_0_dimensionality),
		.flush(flush),
		.ranges(loops_buf2out_autovec_read_0_ranges),
		.rst_n(rst_n),
		.step(t_read[0]),
		.mux_sel_out(loops_buf2out_autovec_read_0_mux_sel_out),
		.restart(loops_buf2out_autovec_read_0_restart)
	);
	sched_gen_6_16_delay_addr_10_4 output_sched_gen_0(
		.clk(clk),
		.clk_en(clk_en),
		.cycle_count(cycle_count),
		.enable(output_sched_gen_0_enable),
		.finished(loops_buf2out_autovec_read_0_restart),
		.flush(flush),
		.mux_sel(loops_buf2out_autovec_read_0_mux_sel_out),
		.rst_n(rst_n),
		.sched_addr_gen_delay(output_sched_gen_0_sched_addr_gen_delay),
		.sched_addr_gen_starting_addr(output_sched_gen_0_sched_addr_gen_starting_addr),
		.sched_addr_gen_strides_0(output_sched_gen_0_sched_addr_gen_strides_0),
		.sched_addr_gen_strides_1(output_sched_gen_0_sched_addr_gen_strides_1),
		.sched_addr_gen_strides_2(output_sched_gen_0_sched_addr_gen_strides_2),
		.sched_addr_gen_strides_3(output_sched_gen_0_sched_addr_gen_strides_3),
		.sched_addr_gen_strides_4(output_sched_gen_0_sched_addr_gen_strides_4),
		.sched_addr_gen_strides_5(output_sched_gen_0_sched_addr_gen_strides_5),
		.valid_output(output_sched_gen_0_valid_output),
		.valid_output_d(output_sched_gen_0_valid_output_d)
	);
	for_loop_6_11 loops_buf2out_autovec_read_1(
		.clk(clk),
		.clk_en(clk_en),
		.dimensionality(loops_buf2out_autovec_read_1_dimensionality),
		.flush(flush),
		.ranges(loops_buf2out_autovec_read_1_ranges),
		.rst_n(rst_n),
		.step(t_read[1]),
		.mux_sel_out(loops_buf2out_autovec_read_1_mux_sel_out),
		.restart(loops_buf2out_autovec_read_1_restart)
	);
	sched_gen_6_16_delay_addr_10_4 output_sched_gen_1(
		.clk(clk),
		.clk_en(clk_en),
		.cycle_count(cycle_count),
		.enable(output_sched_gen_1_enable),
		.finished(loops_buf2out_autovec_read_1_restart),
		.flush(flush),
		.mux_sel(loops_buf2out_autovec_read_1_mux_sel_out),
		.rst_n(rst_n),
		.sched_addr_gen_delay(output_sched_gen_1_sched_addr_gen_delay),
		.sched_addr_gen_starting_addr(output_sched_gen_1_sched_addr_gen_starting_addr),
		.sched_addr_gen_strides_0(output_sched_gen_1_sched_addr_gen_strides_0),
		.sched_addr_gen_strides_1(output_sched_gen_1_sched_addr_gen_strides_1),
		.sched_addr_gen_strides_2(output_sched_gen_1_sched_addr_gen_strides_2),
		.sched_addr_gen_strides_3(output_sched_gen_1_sched_addr_gen_strides_3),
		.sched_addr_gen_strides_4(output_sched_gen_1_sched_addr_gen_strides_4),
		.sched_addr_gen_strides_5(output_sched_gen_1_sched_addr_gen_strides_5),
		.valid_output(output_sched_gen_1_valid_output),
		.valid_output_d(output_sched_gen_1_valid_output_d)
	);
endmodule
module strg_ub_tb_only (
	clk,
	clk_en,
	cycle_count,
	flush,
	loops_buf2out_read_0_dimensionality,
	loops_buf2out_read_0_ranges_0,
	loops_buf2out_read_0_ranges_1,
	loops_buf2out_read_0_ranges_2,
	loops_buf2out_read_0_ranges_3,
	loops_buf2out_read_0_ranges_4,
	loops_buf2out_read_0_ranges_5,
	loops_buf2out_read_1_dimensionality,
	loops_buf2out_read_1_ranges_0,
	loops_buf2out_read_1_ranges_1,
	loops_buf2out_read_1_ranges_2,
	loops_buf2out_read_1_ranges_3,
	loops_buf2out_read_1_ranges_4,
	loops_buf2out_read_1_ranges_5,
	loops_sram2tb_mux_sel,
	loops_sram2tb_restart,
	rst_n,
	shared_tb_0,
	sram_read_data,
	t_read,
	tb_read_addr_gen_0_starting_addr,
	tb_read_addr_gen_0_strides_0,
	tb_read_addr_gen_0_strides_1,
	tb_read_addr_gen_0_strides_2,
	tb_read_addr_gen_0_strides_3,
	tb_read_addr_gen_0_strides_4,
	tb_read_addr_gen_0_strides_5,
	tb_read_addr_gen_1_starting_addr,
	tb_read_addr_gen_1_strides_0,
	tb_read_addr_gen_1_strides_1,
	tb_read_addr_gen_1_strides_2,
	tb_read_addr_gen_1_strides_3,
	tb_read_addr_gen_1_strides_4,
	tb_read_addr_gen_1_strides_5,
	tb_read_sched_gen_0_enable,
	tb_read_sched_gen_0_sched_addr_gen_delay,
	tb_read_sched_gen_0_sched_addr_gen_starting_addr,
	tb_read_sched_gen_0_sched_addr_gen_strides_0,
	tb_read_sched_gen_0_sched_addr_gen_strides_1,
	tb_read_sched_gen_0_sched_addr_gen_strides_2,
	tb_read_sched_gen_0_sched_addr_gen_strides_3,
	tb_read_sched_gen_0_sched_addr_gen_strides_4,
	tb_read_sched_gen_0_sched_addr_gen_strides_5,
	tb_read_sched_gen_1_enable,
	tb_read_sched_gen_1_sched_addr_gen_delay,
	tb_read_sched_gen_1_sched_addr_gen_starting_addr,
	tb_read_sched_gen_1_sched_addr_gen_strides_0,
	tb_read_sched_gen_1_sched_addr_gen_strides_1,
	tb_read_sched_gen_1_sched_addr_gen_strides_2,
	tb_read_sched_gen_1_sched_addr_gen_strides_3,
	tb_read_sched_gen_1_sched_addr_gen_strides_4,
	tb_read_sched_gen_1_sched_addr_gen_strides_5,
	tb_write_addr_gen_0_starting_addr,
	tb_write_addr_gen_0_strides_0,
	tb_write_addr_gen_0_strides_1,
	tb_write_addr_gen_0_strides_2,
	tb_write_addr_gen_0_strides_3,
	tb_write_addr_gen_0_strides_4,
	tb_write_addr_gen_0_strides_5,
	tb_write_addr_gen_1_starting_addr,
	tb_write_addr_gen_1_strides_0,
	tb_write_addr_gen_1_strides_1,
	tb_write_addr_gen_1_strides_2,
	tb_write_addr_gen_1_strides_3,
	tb_write_addr_gen_1_strides_4,
	tb_write_addr_gen_1_strides_5,
	accessor_output,
	data_out,
	tb_read_addr_d_out,
	tb_read_d_out
);
	input wire clk;
	input wire clk_en;
	input wire [15:0] cycle_count;
	input wire flush;
	input wire [3:0] loops_buf2out_read_0_dimensionality;
	input wire [10:0] loops_buf2out_read_0_ranges_0;
	input wire [10:0] loops_buf2out_read_0_ranges_1;
	input wire [10:0] loops_buf2out_read_0_ranges_2;
	input wire [10:0] loops_buf2out_read_0_ranges_3;
	input wire [10:0] loops_buf2out_read_0_ranges_4;
	input wire [10:0] loops_buf2out_read_0_ranges_5;
	input wire [3:0] loops_buf2out_read_1_dimensionality;
	input wire [10:0] loops_buf2out_read_1_ranges_0;
	input wire [10:0] loops_buf2out_read_1_ranges_1;
	input wire [10:0] loops_buf2out_read_1_ranges_2;
	input wire [10:0] loops_buf2out_read_1_ranges_3;
	input wire [10:0] loops_buf2out_read_1_ranges_4;
	input wire [10:0] loops_buf2out_read_1_ranges_5;
	input wire [5:0] loops_sram2tb_mux_sel;
	input wire [1:0] loops_sram2tb_restart;
	input wire rst_n;
	input wire shared_tb_0;
	input wire [63:0] sram_read_data;
	input wire [1:0] t_read;
	input wire [3:0] tb_read_addr_gen_0_starting_addr;
	input wire [3:0] tb_read_addr_gen_0_strides_0;
	input wire [3:0] tb_read_addr_gen_0_strides_1;
	input wire [3:0] tb_read_addr_gen_0_strides_2;
	input wire [3:0] tb_read_addr_gen_0_strides_3;
	input wire [3:0] tb_read_addr_gen_0_strides_4;
	input wire [3:0] tb_read_addr_gen_0_strides_5;
	input wire [3:0] tb_read_addr_gen_1_starting_addr;
	input wire [3:0] tb_read_addr_gen_1_strides_0;
	input wire [3:0] tb_read_addr_gen_1_strides_1;
	input wire [3:0] tb_read_addr_gen_1_strides_2;
	input wire [3:0] tb_read_addr_gen_1_strides_3;
	input wire [3:0] tb_read_addr_gen_1_strides_4;
	input wire [3:0] tb_read_addr_gen_1_strides_5;
	input wire tb_read_sched_gen_0_enable;
	input wire [9:0] tb_read_sched_gen_0_sched_addr_gen_delay;
	input wire [15:0] tb_read_sched_gen_0_sched_addr_gen_starting_addr;
	input wire [15:0] tb_read_sched_gen_0_sched_addr_gen_strides_0;
	input wire [15:0] tb_read_sched_gen_0_sched_addr_gen_strides_1;
	input wire [15:0] tb_read_sched_gen_0_sched_addr_gen_strides_2;
	input wire [15:0] tb_read_sched_gen_0_sched_addr_gen_strides_3;
	input wire [15:0] tb_read_sched_gen_0_sched_addr_gen_strides_4;
	input wire [15:0] tb_read_sched_gen_0_sched_addr_gen_strides_5;
	input wire tb_read_sched_gen_1_enable;
	input wire [9:0] tb_read_sched_gen_1_sched_addr_gen_delay;
	input wire [15:0] tb_read_sched_gen_1_sched_addr_gen_starting_addr;
	input wire [15:0] tb_read_sched_gen_1_sched_addr_gen_strides_0;
	input wire [15:0] tb_read_sched_gen_1_sched_addr_gen_strides_1;
	input wire [15:0] tb_read_sched_gen_1_sched_addr_gen_strides_2;
	input wire [15:0] tb_read_sched_gen_1_sched_addr_gen_strides_3;
	input wire [15:0] tb_read_sched_gen_1_sched_addr_gen_strides_4;
	input wire [15:0] tb_read_sched_gen_1_sched_addr_gen_strides_5;
	input wire [3:0] tb_write_addr_gen_0_starting_addr;
	input wire [3:0] tb_write_addr_gen_0_strides_0;
	input wire [3:0] tb_write_addr_gen_0_strides_1;
	input wire [3:0] tb_write_addr_gen_0_strides_2;
	input wire [3:0] tb_write_addr_gen_0_strides_3;
	input wire [3:0] tb_write_addr_gen_0_strides_4;
	input wire [3:0] tb_write_addr_gen_0_strides_5;
	input wire [3:0] tb_write_addr_gen_1_starting_addr;
	input wire [3:0] tb_write_addr_gen_1_strides_0;
	input wire [3:0] tb_write_addr_gen_1_strides_1;
	input wire [3:0] tb_write_addr_gen_1_strides_2;
	input wire [3:0] tb_write_addr_gen_1_strides_3;
	input wire [3:0] tb_write_addr_gen_1_strides_4;
	input wire [3:0] tb_write_addr_gen_1_strides_5;
	output wire [1:0] accessor_output;
	output reg [31:0] data_out;
	output wire [5:0] tb_read_addr_d_out;
	output wire [1:0] tb_read_d_out;
	wire [2:0] addr_fifo_in_0;
	wire [2:0] addr_fifo_in_1;
	wire delay_en_0;
	wire delay_en_1;
	wire [2:0] loops_buf2out_read_0_mux_sel_out;
	wire [65:0] loops_buf2out_read_0_ranges;
	wire loops_buf2out_read_0_restart;
	wire [2:0] loops_buf2out_read_1_mux_sel_out;
	wire [65:0] loops_buf2out_read_1_ranges;
	wire loops_buf2out_read_1_restart;
	reg [5:0] mux_sel_d1;
	reg [2:0] rd_ptr_0;
	reg [2:0] rd_ptr_1;
	reg [1:0] restart_d1;
	reg [1:0] t_read_d1;
	reg [255:0] tb;
	reg [23:0] tb_addr_fifo_0;
	reg [23:0] tb_addr_fifo_1;
	wire [1:0] tb_read;
	wire [7:0] tb_read_addr;
	wire [3:0] tb_read_addr_gen_0_addr_out;
	wire [23:0] tb_read_addr_gen_0_strides;
	wire [3:0] tb_read_addr_gen_1_addr_out;
	wire [23:0] tb_read_addr_gen_1_strides;
	wire tb_read_d_0;
	wire tb_read_d_1;
	wire tb_read_sched_gen_0_valid_output;
	wire tb_read_sched_gen_1_valid_output;
	wire tb_read_sel_0;
	wire [5:0] tb_write_addr;
	wire [3:0] tb_write_addr_gen_0_addr_out;
	wire [23:0] tb_write_addr_gen_0_strides;
	wire [3:0] tb_write_addr_gen_1_addr_out;
	wire [23:0] tb_write_addr_gen_1_strides;
	wire tb_write_sel_0;
	reg [2:0] wr_ptr_0;
	reg [2:0] wr_ptr_1;
	assign accessor_output = tb_read;
	always @(posedge clk or negedge rst_n)
		if (~rst_n) begin
			t_read_d1[0] <= 1'h0;
			mux_sel_d1[0+:3] <= 3'h0;
			restart_d1[0] <= 1'h0;
		end
		else if (clk_en) begin
			if (flush) begin
				t_read_d1[0] <= 1'h0;
				mux_sel_d1[0+:3] <= 3'h0;
				restart_d1[0] <= 1'h0;
			end
			else begin
				t_read_d1[0] <= t_read[0];
				mux_sel_d1[0+:3] <= loops_sram2tb_mux_sel[0+:3];
				restart_d1[0] <= loops_sram2tb_restart[0];
			end
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n) begin
			t_read_d1[1] <= 1'h0;
			mux_sel_d1[3+:3] <= 3'h0;
			restart_d1[1] <= 1'h0;
		end
		else if (clk_en) begin
			if (flush) begin
				t_read_d1[1] <= 1'h0;
				mux_sel_d1[3+:3] <= 3'h0;
				restart_d1[1] <= 1'h0;
			end
			else begin
				t_read_d1[1] <= t_read[1];
				mux_sel_d1[3+:3] <= loops_sram2tb_mux_sel[3+:3];
				restart_d1[1] <= loops_sram2tb_restart[1];
			end
		end
	assign tb_write_sel_0 = (shared_tb_0 ? tb_write_addr[1] : 1'h0);
	assign tb_read_sel_0 = (shared_tb_0 ? tb_read_addr[3] : 1'h0);
	assign tb_write_addr[0+:3] = tb_write_addr_gen_0_addr_out[2:0];
	assign tb_read_addr[0+:4] = tb_read_addr_gen_0_addr_out;
	assign tb_read[0] = tb_read_sched_gen_0_valid_output;
	assign addr_fifo_in_0 = tb_read_addr_gen_0_addr_out[2:0];
	always @(posedge clk or negedge rst_n)
		if (~rst_n) begin
			wr_ptr_0 <= 3'h0;
			rd_ptr_0 <= 3'h0;
			tb_addr_fifo_0 <= 24'h000000;
		end
		else if (clk_en) begin
			if (flush) begin
				wr_ptr_0 <= 3'h0;
				rd_ptr_0 <= 3'h0;
				tb_addr_fifo_0 <= 24'h000000;
			end
			else if (delay_en_0) begin
				if (tb_read[0]) begin
					tb_addr_fifo_0[wr_ptr_0 * 3+:3] <= addr_fifo_in_0;
					wr_ptr_0 <= wr_ptr_0 + 3'h1;
				end
				if (tb_read_d_0)
					rd_ptr_0 <= rd_ptr_0 + 3'h1;
			end
		end
	assign tb_read_d_out[0] = (delay_en_0 ? tb_read_d_0 : tb_read[0]);
	assign tb_read_addr_d_out[0+:3] = (delay_en_0 ? tb_addr_fifo_0[rd_ptr_0 * 3+:3] : addr_fifo_in_0);
	always @(*) data_out[0+:16] = tb[((((tb_read_sel_0 * 2) + tb_read_addr[2]) * 4) + tb_read_addr[1-:2]) * 16+:16];
	assign tb_write_addr[3+:3] = tb_write_addr_gen_1_addr_out[2:0];
	assign tb_read_addr[4+:4] = tb_read_addr_gen_1_addr_out;
	assign tb_read[1] = tb_read_sched_gen_1_valid_output;
	assign addr_fifo_in_1 = tb_read_addr_gen_1_addr_out[2:0];
	always @(posedge clk or negedge rst_n)
		if (~rst_n) begin
			wr_ptr_1 <= 3'h0;
			rd_ptr_1 <= 3'h0;
			tb_addr_fifo_1 <= 24'h000000;
		end
		else if (clk_en) begin
			if (flush) begin
				wr_ptr_1 <= 3'h0;
				rd_ptr_1 <= 3'h0;
				tb_addr_fifo_1 <= 24'h000000;
			end
			else if (delay_en_1) begin
				if (tb_read[1]) begin
					tb_addr_fifo_1[wr_ptr_1 * 3+:3] <= addr_fifo_in_1;
					wr_ptr_1 <= wr_ptr_1 + 3'h1;
				end
				if (tb_read_d_1)
					rd_ptr_1 <= rd_ptr_1 + 3'h1;
			end
		end
	assign tb_read_d_out[1] = (delay_en_1 ? tb_read_d_1 : tb_read[1]);
	assign tb_read_addr_d_out[3+:3] = (delay_en_1 ? tb_addr_fifo_1[rd_ptr_1 * 3+:3] : addr_fifo_in_1);
	always @(*) data_out[16+:16] = tb[(((2 + tb_read_addr[6]) * 4) + tb_read_addr[5-:2]) * 16+:16];
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	always @(posedge clk)
		if (clk_en) begin : sv2v_autoblock_1
			reg [31:0] i;
			for (i = 0; i < 2; i = i + 1)
				if (t_read_d1[sv2v_cast_1(i)]) begin
					if (i == 32'h00000000)
						tb[16 * (((tb_write_sel_0 * 2) + tb_write_addr[sv2v_cast_1(i) * 3]) * 4)+:64] <= sram_read_data;
					else
						tb[16 * (((sv2v_cast_1(i) * 2) + tb_write_addr[sv2v_cast_1(i) * 3]) * 4)+:64] <= sram_read_data;
				end
		end
	assign tb_write_addr_gen_0_strides[0+:4] = tb_write_addr_gen_0_strides_0;
	assign tb_write_addr_gen_0_strides[4+:4] = tb_write_addr_gen_0_strides_1;
	assign tb_write_addr_gen_0_strides[8+:4] = tb_write_addr_gen_0_strides_2;
	assign tb_write_addr_gen_0_strides[12+:4] = tb_write_addr_gen_0_strides_3;
	assign tb_write_addr_gen_0_strides[16+:4] = tb_write_addr_gen_0_strides_4;
	assign tb_write_addr_gen_0_strides[20+:4] = tb_write_addr_gen_0_strides_5;
	assign loops_buf2out_read_0_ranges[0+:11] = loops_buf2out_read_0_ranges_0;
	assign loops_buf2out_read_0_ranges[11+:11] = loops_buf2out_read_0_ranges_1;
	assign loops_buf2out_read_0_ranges[22+:11] = loops_buf2out_read_0_ranges_2;
	assign loops_buf2out_read_0_ranges[33+:11] = loops_buf2out_read_0_ranges_3;
	assign loops_buf2out_read_0_ranges[44+:11] = loops_buf2out_read_0_ranges_4;
	assign loops_buf2out_read_0_ranges[55+:11] = loops_buf2out_read_0_ranges_5;
	assign tb_read_addr_gen_0_strides[0+:4] = tb_read_addr_gen_0_strides_0;
	assign tb_read_addr_gen_0_strides[4+:4] = tb_read_addr_gen_0_strides_1;
	assign tb_read_addr_gen_0_strides[8+:4] = tb_read_addr_gen_0_strides_2;
	assign tb_read_addr_gen_0_strides[12+:4] = tb_read_addr_gen_0_strides_3;
	assign tb_read_addr_gen_0_strides[16+:4] = tb_read_addr_gen_0_strides_4;
	assign tb_read_addr_gen_0_strides[20+:4] = tb_read_addr_gen_0_strides_5;
	assign tb_write_addr_gen_1_strides[0+:4] = tb_write_addr_gen_1_strides_0;
	assign tb_write_addr_gen_1_strides[4+:4] = tb_write_addr_gen_1_strides_1;
	assign tb_write_addr_gen_1_strides[8+:4] = tb_write_addr_gen_1_strides_2;
	assign tb_write_addr_gen_1_strides[12+:4] = tb_write_addr_gen_1_strides_3;
	assign tb_write_addr_gen_1_strides[16+:4] = tb_write_addr_gen_1_strides_4;
	assign tb_write_addr_gen_1_strides[20+:4] = tb_write_addr_gen_1_strides_5;
	assign loops_buf2out_read_1_ranges[0+:11] = loops_buf2out_read_1_ranges_0;
	assign loops_buf2out_read_1_ranges[11+:11] = loops_buf2out_read_1_ranges_1;
	assign loops_buf2out_read_1_ranges[22+:11] = loops_buf2out_read_1_ranges_2;
	assign loops_buf2out_read_1_ranges[33+:11] = loops_buf2out_read_1_ranges_3;
	assign loops_buf2out_read_1_ranges[44+:11] = loops_buf2out_read_1_ranges_4;
	assign loops_buf2out_read_1_ranges[55+:11] = loops_buf2out_read_1_ranges_5;
	assign tb_read_addr_gen_1_strides[0+:4] = tb_read_addr_gen_1_strides_0;
	assign tb_read_addr_gen_1_strides[4+:4] = tb_read_addr_gen_1_strides_1;
	assign tb_read_addr_gen_1_strides[8+:4] = tb_read_addr_gen_1_strides_2;
	assign tb_read_addr_gen_1_strides[12+:4] = tb_read_addr_gen_1_strides_3;
	assign tb_read_addr_gen_1_strides[16+:4] = tb_read_addr_gen_1_strides_4;
	assign tb_read_addr_gen_1_strides[20+:4] = tb_read_addr_gen_1_strides_5;
	addr_gen_6_4 tb_write_addr_gen_0(
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.mux_sel(mux_sel_d1[0+:3]),
		.restart(restart_d1[0]),
		.rst_n(rst_n),
		.starting_addr(tb_write_addr_gen_0_starting_addr),
		.step(t_read_d1[0]),
		.strides(tb_write_addr_gen_0_strides),
		.addr_out(tb_write_addr_gen_0_addr_out)
	);
	for_loop_6_11 loops_buf2out_read_0(
		.clk(clk),
		.clk_en(clk_en),
		.dimensionality(loops_buf2out_read_0_dimensionality),
		.flush(flush),
		.ranges(loops_buf2out_read_0_ranges),
		.rst_n(rst_n),
		.step(tb_read[0]),
		.mux_sel_out(loops_buf2out_read_0_mux_sel_out),
		.restart(loops_buf2out_read_0_restart)
	);
	addr_gen_6_4 tb_read_addr_gen_0(
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.mux_sel(loops_buf2out_read_0_mux_sel_out),
		.restart(loops_buf2out_read_0_restart),
		.rst_n(rst_n),
		.starting_addr(tb_read_addr_gen_0_starting_addr),
		.step(tb_read[0]),
		.strides(tb_read_addr_gen_0_strides),
		.addr_out(tb_read_addr_gen_0_addr_out)
	);
	sched_gen_6_16_delay_addr_10_8 tb_read_sched_gen_0(
		.clk(clk),
		.clk_en(clk_en),
		.cycle_count(cycle_count),
		.enable(tb_read_sched_gen_0_enable),
		.finished(loops_buf2out_read_0_restart),
		.flush(flush),
		.mux_sel(loops_buf2out_read_0_mux_sel_out),
		.rst_n(rst_n),
		.sched_addr_gen_delay(tb_read_sched_gen_0_sched_addr_gen_delay),
		.sched_addr_gen_starting_addr(tb_read_sched_gen_0_sched_addr_gen_starting_addr),
		.sched_addr_gen_strides_0(tb_read_sched_gen_0_sched_addr_gen_strides_0),
		.sched_addr_gen_strides_1(tb_read_sched_gen_0_sched_addr_gen_strides_1),
		.sched_addr_gen_strides_2(tb_read_sched_gen_0_sched_addr_gen_strides_2),
		.sched_addr_gen_strides_3(tb_read_sched_gen_0_sched_addr_gen_strides_3),
		.sched_addr_gen_strides_4(tb_read_sched_gen_0_sched_addr_gen_strides_4),
		.sched_addr_gen_strides_5(tb_read_sched_gen_0_sched_addr_gen_strides_5),
		.delay_en_out(delay_en_0),
		.valid_output(tb_read_sched_gen_0_valid_output),
		.valid_output_d(tb_read_d_0)
	);
	addr_gen_6_4 tb_write_addr_gen_1(
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.mux_sel(mux_sel_d1[3+:3]),
		.restart(restart_d1[1]),
		.rst_n(rst_n),
		.starting_addr(tb_write_addr_gen_1_starting_addr),
		.step(t_read_d1[1]),
		.strides(tb_write_addr_gen_1_strides),
		.addr_out(tb_write_addr_gen_1_addr_out)
	);
	for_loop_6_11 loops_buf2out_read_1(
		.clk(clk),
		.clk_en(clk_en),
		.dimensionality(loops_buf2out_read_1_dimensionality),
		.flush(flush),
		.ranges(loops_buf2out_read_1_ranges),
		.rst_n(rst_n),
		.step(tb_read[1]),
		.mux_sel_out(loops_buf2out_read_1_mux_sel_out),
		.restart(loops_buf2out_read_1_restart)
	);
	addr_gen_6_4 tb_read_addr_gen_1(
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.mux_sel(loops_buf2out_read_1_mux_sel_out),
		.restart(loops_buf2out_read_1_restart),
		.rst_n(rst_n),
		.starting_addr(tb_read_addr_gen_1_starting_addr),
		.step(tb_read[1]),
		.strides(tb_read_addr_gen_1_strides),
		.addr_out(tb_read_addr_gen_1_addr_out)
	);
	sched_gen_6_16_delay_addr_10_8 tb_read_sched_gen_1(
		.clk(clk),
		.clk_en(clk_en),
		.cycle_count(cycle_count),
		.enable(tb_read_sched_gen_1_enable),
		.finished(loops_buf2out_read_1_restart),
		.flush(flush),
		.mux_sel(loops_buf2out_read_1_mux_sel_out),
		.rst_n(rst_n),
		.sched_addr_gen_delay(tb_read_sched_gen_1_sched_addr_gen_delay),
		.sched_addr_gen_starting_addr(tb_read_sched_gen_1_sched_addr_gen_starting_addr),
		.sched_addr_gen_strides_0(tb_read_sched_gen_1_sched_addr_gen_strides_0),
		.sched_addr_gen_strides_1(tb_read_sched_gen_1_sched_addr_gen_strides_1),
		.sched_addr_gen_strides_2(tb_read_sched_gen_1_sched_addr_gen_strides_2),
		.sched_addr_gen_strides_3(tb_read_sched_gen_1_sched_addr_gen_strides_3),
		.sched_addr_gen_strides_4(tb_read_sched_gen_1_sched_addr_gen_strides_4),
		.sched_addr_gen_strides_5(tb_read_sched_gen_1_sched_addr_gen_strides_5),
		.delay_en_out(delay_en_1),
		.valid_output(tb_read_sched_gen_1_valid_output),
		.valid_output_d(tb_read_d_1)
	);
endmodule
module strg_ub_vec (
	agg_only_agg_write_addr_gen_0_starting_addr,
	agg_only_agg_write_addr_gen_0_strides_0,
	agg_only_agg_write_addr_gen_0_strides_1,
	agg_only_agg_write_addr_gen_0_strides_2,
	agg_only_agg_write_addr_gen_1_starting_addr,
	agg_only_agg_write_addr_gen_1_strides_0,
	agg_only_agg_write_addr_gen_1_strides_1,
	agg_only_agg_write_addr_gen_1_strides_2,
	agg_only_agg_write_sched_gen_0_enable,
	agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr,
	agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0,
	agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1,
	agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2,
	agg_only_agg_write_sched_gen_1_enable,
	agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr,
	agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0,
	agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1,
	agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2,
	agg_only_loops_in2buf_0_dimensionality,
	agg_only_loops_in2buf_0_ranges_0,
	agg_only_loops_in2buf_0_ranges_1,
	agg_only_loops_in2buf_0_ranges_2,
	agg_only_loops_in2buf_1_dimensionality,
	agg_only_loops_in2buf_1_ranges_0,
	agg_only_loops_in2buf_1_ranges_1,
	agg_only_loops_in2buf_1_ranges_2,
	agg_sram_shared_agg_read_sched_gen_0_agg_read_padding,
	agg_sram_shared_agg_read_sched_gen_1_agg_read_padding,
	agg_sram_shared_agg_sram_shared_addr_gen_0_starting_addr,
	agg_sram_shared_agg_sram_shared_addr_gen_1_starting_addr,
	agg_sram_shared_mode_0,
	agg_sram_shared_mode_1,
	chain_chain_en,
	chain_data_in,
	clk,
	clk_en,
	data_from_strg,
	data_in,
	flush,
	rst_n,
	sram_only_output_addr_gen_0_starting_addr,
	sram_only_output_addr_gen_0_strides_0,
	sram_only_output_addr_gen_0_strides_1,
	sram_only_output_addr_gen_0_strides_2,
	sram_only_output_addr_gen_0_strides_3,
	sram_only_output_addr_gen_0_strides_4,
	sram_only_output_addr_gen_0_strides_5,
	sram_only_output_addr_gen_1_starting_addr,
	sram_only_output_addr_gen_1_strides_0,
	sram_only_output_addr_gen_1_strides_1,
	sram_only_output_addr_gen_1_strides_2,
	sram_only_output_addr_gen_1_strides_3,
	sram_only_output_addr_gen_1_strides_4,
	sram_only_output_addr_gen_1_strides_5,
	sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality,
	sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0,
	sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1,
	sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2,
	sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3,
	sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4,
	sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5,
	sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality,
	sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0,
	sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1,
	sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2,
	sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3,
	sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4,
	sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5,
	sram_tb_shared_output_sched_gen_0_enable,
	sram_tb_shared_output_sched_gen_0_sched_addr_gen_delay,
	sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr,
	sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0,
	sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1,
	sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2,
	sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3,
	sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4,
	sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5,
	sram_tb_shared_output_sched_gen_1_enable,
	sram_tb_shared_output_sched_gen_1_sched_addr_gen_delay,
	sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr,
	sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0,
	sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1,
	sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2,
	sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3,
	sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4,
	sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5,
	tb_only_loops_buf2out_read_0_dimensionality,
	tb_only_loops_buf2out_read_0_ranges_0,
	tb_only_loops_buf2out_read_0_ranges_1,
	tb_only_loops_buf2out_read_0_ranges_2,
	tb_only_loops_buf2out_read_0_ranges_3,
	tb_only_loops_buf2out_read_0_ranges_4,
	tb_only_loops_buf2out_read_0_ranges_5,
	tb_only_loops_buf2out_read_1_dimensionality,
	tb_only_loops_buf2out_read_1_ranges_0,
	tb_only_loops_buf2out_read_1_ranges_1,
	tb_only_loops_buf2out_read_1_ranges_2,
	tb_only_loops_buf2out_read_1_ranges_3,
	tb_only_loops_buf2out_read_1_ranges_4,
	tb_only_loops_buf2out_read_1_ranges_5,
	tb_only_shared_tb_0,
	tb_only_tb_read_addr_gen_0_starting_addr,
	tb_only_tb_read_addr_gen_0_strides_0,
	tb_only_tb_read_addr_gen_0_strides_1,
	tb_only_tb_read_addr_gen_0_strides_2,
	tb_only_tb_read_addr_gen_0_strides_3,
	tb_only_tb_read_addr_gen_0_strides_4,
	tb_only_tb_read_addr_gen_0_strides_5,
	tb_only_tb_read_addr_gen_1_starting_addr,
	tb_only_tb_read_addr_gen_1_strides_0,
	tb_only_tb_read_addr_gen_1_strides_1,
	tb_only_tb_read_addr_gen_1_strides_2,
	tb_only_tb_read_addr_gen_1_strides_3,
	tb_only_tb_read_addr_gen_1_strides_4,
	tb_only_tb_read_addr_gen_1_strides_5,
	tb_only_tb_read_sched_gen_0_enable,
	tb_only_tb_read_sched_gen_0_sched_addr_gen_delay,
	tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr,
	tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0,
	tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1,
	tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2,
	tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3,
	tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4,
	tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5,
	tb_only_tb_read_sched_gen_1_enable,
	tb_only_tb_read_sched_gen_1_sched_addr_gen_delay,
	tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr,
	tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0,
	tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1,
	tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2,
	tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3,
	tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4,
	tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5,
	tb_only_tb_write_addr_gen_0_starting_addr,
	tb_only_tb_write_addr_gen_0_strides_0,
	tb_only_tb_write_addr_gen_0_strides_1,
	tb_only_tb_write_addr_gen_0_strides_2,
	tb_only_tb_write_addr_gen_0_strides_3,
	tb_only_tb_write_addr_gen_0_strides_4,
	tb_only_tb_write_addr_gen_0_strides_5,
	tb_only_tb_write_addr_gen_1_starting_addr,
	tb_only_tb_write_addr_gen_1_strides_0,
	tb_only_tb_write_addr_gen_1_strides_1,
	tb_only_tb_write_addr_gen_1_strides_2,
	tb_only_tb_write_addr_gen_1_strides_3,
	tb_only_tb_write_addr_gen_1_strides_4,
	tb_only_tb_write_addr_gen_1_strides_5,
	accessor_output,
	addr_out,
	data_out,
	data_to_strg,
	ren_to_strg,
	wen_to_strg
);
	input wire [2:0] agg_only_agg_write_addr_gen_0_starting_addr;
	input wire [2:0] agg_only_agg_write_addr_gen_0_strides_0;
	input wire [2:0] agg_only_agg_write_addr_gen_0_strides_1;
	input wire [2:0] agg_only_agg_write_addr_gen_0_strides_2;
	input wire [2:0] agg_only_agg_write_addr_gen_1_starting_addr;
	input wire [2:0] agg_only_agg_write_addr_gen_1_strides_0;
	input wire [2:0] agg_only_agg_write_addr_gen_1_strides_1;
	input wire [2:0] agg_only_agg_write_addr_gen_1_strides_2;
	input wire agg_only_agg_write_sched_gen_0_enable;
	input wire [15:0] agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr;
	input wire [15:0] agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0;
	input wire [15:0] agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1;
	input wire [15:0] agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2;
	input wire agg_only_agg_write_sched_gen_1_enable;
	input wire [15:0] agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr;
	input wire [15:0] agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0;
	input wire [15:0] agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1;
	input wire [15:0] agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2;
	input wire [2:0] agg_only_loops_in2buf_0_dimensionality;
	input wire [10:0] agg_only_loops_in2buf_0_ranges_0;
	input wire [10:0] agg_only_loops_in2buf_0_ranges_1;
	input wire [10:0] agg_only_loops_in2buf_0_ranges_2;
	input wire [2:0] agg_only_loops_in2buf_1_dimensionality;
	input wire [10:0] agg_only_loops_in2buf_1_ranges_0;
	input wire [10:0] agg_only_loops_in2buf_1_ranges_1;
	input wire [10:0] agg_only_loops_in2buf_1_ranges_2;
	input wire [7:0] agg_sram_shared_agg_read_sched_gen_0_agg_read_padding;
	input wire [7:0] agg_sram_shared_agg_read_sched_gen_1_agg_read_padding;
	input wire [8:0] agg_sram_shared_agg_sram_shared_addr_gen_0_starting_addr;
	input wire [8:0] agg_sram_shared_agg_sram_shared_addr_gen_1_starting_addr;
	input wire [1:0] agg_sram_shared_mode_0;
	input wire [1:0] agg_sram_shared_mode_1;
	input wire chain_chain_en;
	input wire [33:0] chain_data_in;
	input wire clk;
	input wire clk_en;
	input wire [63:0] data_from_strg;
	input wire [33:0] data_in;
	input wire flush;
	input wire rst_n;
	input wire [8:0] sram_only_output_addr_gen_0_starting_addr;
	input wire [8:0] sram_only_output_addr_gen_0_strides_0;
	input wire [8:0] sram_only_output_addr_gen_0_strides_1;
	input wire [8:0] sram_only_output_addr_gen_0_strides_2;
	input wire [8:0] sram_only_output_addr_gen_0_strides_3;
	input wire [8:0] sram_only_output_addr_gen_0_strides_4;
	input wire [8:0] sram_only_output_addr_gen_0_strides_5;
	input wire [8:0] sram_only_output_addr_gen_1_starting_addr;
	input wire [8:0] sram_only_output_addr_gen_1_strides_0;
	input wire [8:0] sram_only_output_addr_gen_1_strides_1;
	input wire [8:0] sram_only_output_addr_gen_1_strides_2;
	input wire [8:0] sram_only_output_addr_gen_1_strides_3;
	input wire [8:0] sram_only_output_addr_gen_1_strides_4;
	input wire [8:0] sram_only_output_addr_gen_1_strides_5;
	input wire [3:0] sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality;
	input wire [10:0] sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0;
	input wire [10:0] sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1;
	input wire [10:0] sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2;
	input wire [10:0] sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3;
	input wire [10:0] sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4;
	input wire [10:0] sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5;
	input wire [3:0] sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality;
	input wire [10:0] sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0;
	input wire [10:0] sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1;
	input wire [10:0] sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2;
	input wire [10:0] sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3;
	input wire [10:0] sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4;
	input wire [10:0] sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5;
	input wire sram_tb_shared_output_sched_gen_0_enable;
	input wire [9:0] sram_tb_shared_output_sched_gen_0_sched_addr_gen_delay;
	input wire [15:0] sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr;
	input wire [15:0] sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0;
	input wire [15:0] sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1;
	input wire [15:0] sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2;
	input wire [15:0] sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3;
	input wire [15:0] sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4;
	input wire [15:0] sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5;
	input wire sram_tb_shared_output_sched_gen_1_enable;
	input wire [9:0] sram_tb_shared_output_sched_gen_1_sched_addr_gen_delay;
	input wire [15:0] sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr;
	input wire [15:0] sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0;
	input wire [15:0] sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1;
	input wire [15:0] sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2;
	input wire [15:0] sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3;
	input wire [15:0] sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4;
	input wire [15:0] sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5;
	input wire [3:0] tb_only_loops_buf2out_read_0_dimensionality;
	input wire [10:0] tb_only_loops_buf2out_read_0_ranges_0;
	input wire [10:0] tb_only_loops_buf2out_read_0_ranges_1;
	input wire [10:0] tb_only_loops_buf2out_read_0_ranges_2;
	input wire [10:0] tb_only_loops_buf2out_read_0_ranges_3;
	input wire [10:0] tb_only_loops_buf2out_read_0_ranges_4;
	input wire [10:0] tb_only_loops_buf2out_read_0_ranges_5;
	input wire [3:0] tb_only_loops_buf2out_read_1_dimensionality;
	input wire [10:0] tb_only_loops_buf2out_read_1_ranges_0;
	input wire [10:0] tb_only_loops_buf2out_read_1_ranges_1;
	input wire [10:0] tb_only_loops_buf2out_read_1_ranges_2;
	input wire [10:0] tb_only_loops_buf2out_read_1_ranges_3;
	input wire [10:0] tb_only_loops_buf2out_read_1_ranges_4;
	input wire [10:0] tb_only_loops_buf2out_read_1_ranges_5;
	input wire tb_only_shared_tb_0;
	input wire [3:0] tb_only_tb_read_addr_gen_0_starting_addr;
	input wire [3:0] tb_only_tb_read_addr_gen_0_strides_0;
	input wire [3:0] tb_only_tb_read_addr_gen_0_strides_1;
	input wire [3:0] tb_only_tb_read_addr_gen_0_strides_2;
	input wire [3:0] tb_only_tb_read_addr_gen_0_strides_3;
	input wire [3:0] tb_only_tb_read_addr_gen_0_strides_4;
	input wire [3:0] tb_only_tb_read_addr_gen_0_strides_5;
	input wire [3:0] tb_only_tb_read_addr_gen_1_starting_addr;
	input wire [3:0] tb_only_tb_read_addr_gen_1_strides_0;
	input wire [3:0] tb_only_tb_read_addr_gen_1_strides_1;
	input wire [3:0] tb_only_tb_read_addr_gen_1_strides_2;
	input wire [3:0] tb_only_tb_read_addr_gen_1_strides_3;
	input wire [3:0] tb_only_tb_read_addr_gen_1_strides_4;
	input wire [3:0] tb_only_tb_read_addr_gen_1_strides_5;
	input wire tb_only_tb_read_sched_gen_0_enable;
	input wire [9:0] tb_only_tb_read_sched_gen_0_sched_addr_gen_delay;
	input wire [15:0] tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr;
	input wire [15:0] tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0;
	input wire [15:0] tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1;
	input wire [15:0] tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2;
	input wire [15:0] tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3;
	input wire [15:0] tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4;
	input wire [15:0] tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5;
	input wire tb_only_tb_read_sched_gen_1_enable;
	input wire [9:0] tb_only_tb_read_sched_gen_1_sched_addr_gen_delay;
	input wire [15:0] tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr;
	input wire [15:0] tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0;
	input wire [15:0] tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1;
	input wire [15:0] tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2;
	input wire [15:0] tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3;
	input wire [15:0] tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4;
	input wire [15:0] tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5;
	input wire [3:0] tb_only_tb_write_addr_gen_0_starting_addr;
	input wire [3:0] tb_only_tb_write_addr_gen_0_strides_0;
	input wire [3:0] tb_only_tb_write_addr_gen_0_strides_1;
	input wire [3:0] tb_only_tb_write_addr_gen_0_strides_2;
	input wire [3:0] tb_only_tb_write_addr_gen_0_strides_3;
	input wire [3:0] tb_only_tb_write_addr_gen_0_strides_4;
	input wire [3:0] tb_only_tb_write_addr_gen_0_strides_5;
	input wire [3:0] tb_only_tb_write_addr_gen_1_starting_addr;
	input wire [3:0] tb_only_tb_write_addr_gen_1_strides_0;
	input wire [3:0] tb_only_tb_write_addr_gen_1_strides_1;
	input wire [3:0] tb_only_tb_write_addr_gen_1_strides_2;
	input wire [3:0] tb_only_tb_write_addr_gen_1_strides_3;
	input wire [3:0] tb_only_tb_write_addr_gen_1_strides_4;
	input wire [3:0] tb_only_tb_write_addr_gen_1_strides_5;
	output wire [1:0] accessor_output;
	output wire [8:0] addr_out;
	output wire [33:0] data_out;
	output wire [63:0] data_to_strg;
	output wire ren_to_strg;
	output wire wen_to_strg;
	wire [1:0] accessor_output_int;
	wire [127:0] agg_only_agg_data_out;
	wire [1:0] agg_only_agg_read;
	wire [3:0] agg_only_agg_write_addr_l2b_out;
	wire [5:0] agg_only_agg_write_mux_sel_out;
	wire [1:0] agg_only_agg_write_out;
	wire [1:0] agg_only_agg_write_restart_out;
	wire [17:0] agg_only_sram_read_addr_in;
	wire [5:0] agg_only_tb_read_addr_d_in;
	wire [1:0] agg_only_tb_read_d_in;
	wire [3:0] agg_only_update_mode_in;
	wire [1:0] agg_sram_shared_agg_read_out;
	wire [17:0] agg_sram_shared_agg_sram_shared_addr_out;
	wire [17:0] agg_sram_shared_sram_read_addr_in;
	wire [1:0] agg_sram_shared_sram_read_d_in;
	wire [1:0] agg_sram_shared_sram_read_in;
	wire [31:0] chain_data_in_thin;
	reg [15:0] cycle_count;
	wire [31:0] data_in_thin;
	wire [31:0] data_out_int;
	wire [31:0] data_out_int_thin;
	wire [5:0] sram_only_loops_sram2tb_mux_sel;
	wire [1:0] sram_only_loops_sram2tb_restart;
	wire [1:0] sram_only_t_read;
	wire [5:0] sram_tb_shared_loops_sram2tb_mux_sel;
	wire [1:0] sram_tb_shared_loops_sram2tb_restart;
	wire [1:0] sram_tb_shared_t_read_out;
	assign data_in_thin[0+:16] = data_in[15-:16];
	assign data_in_thin[16+:16] = data_in[32-:16];
	assign data_out[15-:16] = data_out_int_thin[0+:16];
	assign data_out[16] = 1'h0;
	assign data_out[32-:16] = data_out_int_thin[16+:16];
	assign data_out[33] = 1'h0;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			cycle_count <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				cycle_count <= 16'h0000;
			else
				cycle_count <= cycle_count + 16'h0001;
		end
	assign agg_only_sram_read_addr_in = agg_sram_shared_agg_sram_shared_addr_out;
	assign agg_sram_shared_sram_read_in = sram_tb_shared_t_read_out;
	assign agg_only_agg_read = agg_sram_shared_agg_read_out;
	assign sram_only_loops_sram2tb_mux_sel = sram_tb_shared_loops_sram2tb_mux_sel;
	assign sram_only_loops_sram2tb_restart = sram_tb_shared_loops_sram2tb_restart;
	assign sram_only_t_read = sram_tb_shared_t_read_out;
	assign ren_to_strg = |sram_tb_shared_t_read_out;
	assign chain_data_in_thin[0+:16] = chain_data_in[15-:16];
	assign chain_data_in_thin[16+:16] = chain_data_in[32-:16];
	assign accessor_output = accessor_output_int;
	strg_ub_agg_only agg_only(
		.agg_read(agg_only_agg_read),
		.agg_write_addr_gen_0_starting_addr(agg_only_agg_write_addr_gen_0_starting_addr),
		.agg_write_addr_gen_0_strides_0(agg_only_agg_write_addr_gen_0_strides_0),
		.agg_write_addr_gen_0_strides_1(agg_only_agg_write_addr_gen_0_strides_1),
		.agg_write_addr_gen_0_strides_2(agg_only_agg_write_addr_gen_0_strides_2),
		.agg_write_addr_gen_1_starting_addr(agg_only_agg_write_addr_gen_1_starting_addr),
		.agg_write_addr_gen_1_strides_0(agg_only_agg_write_addr_gen_1_strides_0),
		.agg_write_addr_gen_1_strides_1(agg_only_agg_write_addr_gen_1_strides_1),
		.agg_write_addr_gen_1_strides_2(agg_only_agg_write_addr_gen_1_strides_2),
		.agg_write_sched_gen_0_enable(agg_only_agg_write_sched_gen_0_enable),
		.agg_write_sched_gen_0_sched_addr_gen_starting_addr(agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr),
		.agg_write_sched_gen_0_sched_addr_gen_strides_0(agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0),
		.agg_write_sched_gen_0_sched_addr_gen_strides_1(agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1),
		.agg_write_sched_gen_0_sched_addr_gen_strides_2(agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2),
		.agg_write_sched_gen_1_enable(agg_only_agg_write_sched_gen_1_enable),
		.agg_write_sched_gen_1_sched_addr_gen_starting_addr(agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr),
		.agg_write_sched_gen_1_sched_addr_gen_strides_0(agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0),
		.agg_write_sched_gen_1_sched_addr_gen_strides_1(agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1),
		.agg_write_sched_gen_1_sched_addr_gen_strides_2(agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2),
		.clk(clk),
		.clk_en(clk_en),
		.cycle_count(cycle_count),
		.data_in(data_in_thin),
		.flush(flush),
		.loops_in2buf_0_dimensionality(agg_only_loops_in2buf_0_dimensionality),
		.loops_in2buf_0_ranges_0(agg_only_loops_in2buf_0_ranges_0),
		.loops_in2buf_0_ranges_1(agg_only_loops_in2buf_0_ranges_1),
		.loops_in2buf_0_ranges_2(agg_only_loops_in2buf_0_ranges_2),
		.loops_in2buf_1_dimensionality(agg_only_loops_in2buf_1_dimensionality),
		.loops_in2buf_1_ranges_0(agg_only_loops_in2buf_1_ranges_0),
		.loops_in2buf_1_ranges_1(agg_only_loops_in2buf_1_ranges_1),
		.loops_in2buf_1_ranges_2(agg_only_loops_in2buf_1_ranges_2),
		.rst_n(rst_n),
		.sram_read_addr_in(agg_only_sram_read_addr_in),
		.tb_read_addr_d_in(agg_only_tb_read_addr_d_in),
		.tb_read_d_in(agg_only_tb_read_d_in),
		.update_mode_in(agg_only_update_mode_in),
		.agg_data_out(agg_only_agg_data_out),
		.agg_write_addr_l2b_out(agg_only_agg_write_addr_l2b_out),
		.agg_write_mux_sel_out(agg_only_agg_write_mux_sel_out),
		.agg_write_out(agg_only_agg_write_out),
		.agg_write_restart_out(agg_only_agg_write_restart_out)
	);
	strg_ub_agg_sram_shared agg_sram_shared(
		.agg_read_sched_gen_0_agg_read_padding(agg_sram_shared_agg_read_sched_gen_0_agg_read_padding),
		.agg_read_sched_gen_1_agg_read_padding(agg_sram_shared_agg_read_sched_gen_1_agg_read_padding),
		.agg_sram_shared_addr_gen_0_starting_addr(agg_sram_shared_agg_sram_shared_addr_gen_0_starting_addr),
		.agg_sram_shared_addr_gen_1_starting_addr(agg_sram_shared_agg_sram_shared_addr_gen_1_starting_addr),
		.agg_write_addr_l2b_in(agg_only_agg_write_addr_l2b_out),
		.agg_write_in(agg_only_agg_write_out),
		.agg_write_mux_sel_in(agg_only_agg_write_mux_sel_out),
		.agg_write_restart_in(agg_only_agg_write_restart_out),
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.mode_0(agg_sram_shared_mode_0),
		.mode_1(agg_sram_shared_mode_1),
		.rst_n(rst_n),
		.sram_read_addr_in(agg_sram_shared_sram_read_addr_in),
		.sram_read_d_in(agg_sram_shared_sram_read_d_in),
		.sram_read_in(agg_sram_shared_sram_read_in),
		.agg_read_out(agg_sram_shared_agg_read_out),
		.agg_sram_shared_addr_out(agg_sram_shared_agg_sram_shared_addr_out),
		.update_mode_out(agg_only_update_mode_in)
	);
	strg_ub_sram_only sram_only(
		.agg_data_out(agg_only_agg_data_out),
		.agg_read(agg_sram_shared_agg_read_out),
		.clk(clk),
		.clk_en(clk_en),
		.cycle_count(cycle_count),
		.flush(flush),
		.loops_sram2tb_mux_sel(sram_only_loops_sram2tb_mux_sel),
		.loops_sram2tb_restart(sram_only_loops_sram2tb_restart),
		.output_addr_gen_0_starting_addr(sram_only_output_addr_gen_0_starting_addr),
		.output_addr_gen_0_strides_0(sram_only_output_addr_gen_0_strides_0),
		.output_addr_gen_0_strides_1(sram_only_output_addr_gen_0_strides_1),
		.output_addr_gen_0_strides_2(sram_only_output_addr_gen_0_strides_2),
		.output_addr_gen_0_strides_3(sram_only_output_addr_gen_0_strides_3),
		.output_addr_gen_0_strides_4(sram_only_output_addr_gen_0_strides_4),
		.output_addr_gen_0_strides_5(sram_only_output_addr_gen_0_strides_5),
		.output_addr_gen_1_starting_addr(sram_only_output_addr_gen_1_starting_addr),
		.output_addr_gen_1_strides_0(sram_only_output_addr_gen_1_strides_0),
		.output_addr_gen_1_strides_1(sram_only_output_addr_gen_1_strides_1),
		.output_addr_gen_1_strides_2(sram_only_output_addr_gen_1_strides_2),
		.output_addr_gen_1_strides_3(sram_only_output_addr_gen_1_strides_3),
		.output_addr_gen_1_strides_4(sram_only_output_addr_gen_1_strides_4),
		.output_addr_gen_1_strides_5(sram_only_output_addr_gen_1_strides_5),
		.rst_n(rst_n),
		.sram_read_addr_in(agg_sram_shared_agg_sram_shared_addr_out),
		.t_read(sram_only_t_read),
		.addr_to_sram(addr_out),
		.data_to_sram(data_to_strg),
		.sram_read_addr_out(agg_sram_shared_sram_read_addr_in),
		.wen_to_sram(wen_to_strg)
	);
	strg_ub_sram_tb_shared sram_tb_shared(
		.clk(clk),
		.clk_en(clk_en),
		.cycle_count(cycle_count),
		.flush(flush),
		.loops_buf2out_autovec_read_0_dimensionality(sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality),
		.loops_buf2out_autovec_read_0_ranges_0(sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0),
		.loops_buf2out_autovec_read_0_ranges_1(sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1),
		.loops_buf2out_autovec_read_0_ranges_2(sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2),
		.loops_buf2out_autovec_read_0_ranges_3(sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3),
		.loops_buf2out_autovec_read_0_ranges_4(sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4),
		.loops_buf2out_autovec_read_0_ranges_5(sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5),
		.loops_buf2out_autovec_read_1_dimensionality(sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality),
		.loops_buf2out_autovec_read_1_ranges_0(sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0),
		.loops_buf2out_autovec_read_1_ranges_1(sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1),
		.loops_buf2out_autovec_read_1_ranges_2(sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2),
		.loops_buf2out_autovec_read_1_ranges_3(sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3),
		.loops_buf2out_autovec_read_1_ranges_4(sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4),
		.loops_buf2out_autovec_read_1_ranges_5(sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5),
		.output_sched_gen_0_enable(sram_tb_shared_output_sched_gen_0_enable),
		.output_sched_gen_0_sched_addr_gen_delay(sram_tb_shared_output_sched_gen_0_sched_addr_gen_delay),
		.output_sched_gen_0_sched_addr_gen_starting_addr(sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr),
		.output_sched_gen_0_sched_addr_gen_strides_0(sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0),
		.output_sched_gen_0_sched_addr_gen_strides_1(sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1),
		.output_sched_gen_0_sched_addr_gen_strides_2(sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2),
		.output_sched_gen_0_sched_addr_gen_strides_3(sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3),
		.output_sched_gen_0_sched_addr_gen_strides_4(sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4),
		.output_sched_gen_0_sched_addr_gen_strides_5(sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5),
		.output_sched_gen_1_enable(sram_tb_shared_output_sched_gen_1_enable),
		.output_sched_gen_1_sched_addr_gen_delay(sram_tb_shared_output_sched_gen_1_sched_addr_gen_delay),
		.output_sched_gen_1_sched_addr_gen_starting_addr(sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr),
		.output_sched_gen_1_sched_addr_gen_strides_0(sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0),
		.output_sched_gen_1_sched_addr_gen_strides_1(sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1),
		.output_sched_gen_1_sched_addr_gen_strides_2(sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2),
		.output_sched_gen_1_sched_addr_gen_strides_3(sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3),
		.output_sched_gen_1_sched_addr_gen_strides_4(sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4),
		.output_sched_gen_1_sched_addr_gen_strides_5(sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5),
		.rst_n(rst_n),
		.loops_sram2tb_mux_sel(sram_tb_shared_loops_sram2tb_mux_sel),
		.loops_sram2tb_restart(sram_tb_shared_loops_sram2tb_restart),
		.sram_read_d(agg_sram_shared_sram_read_d_in),
		.t_read_out(sram_tb_shared_t_read_out)
	);
	strg_ub_tb_only tb_only(
		.clk(clk),
		.clk_en(clk_en),
		.cycle_count(cycle_count),
		.flush(flush),
		.loops_buf2out_read_0_dimensionality(tb_only_loops_buf2out_read_0_dimensionality),
		.loops_buf2out_read_0_ranges_0(tb_only_loops_buf2out_read_0_ranges_0),
		.loops_buf2out_read_0_ranges_1(tb_only_loops_buf2out_read_0_ranges_1),
		.loops_buf2out_read_0_ranges_2(tb_only_loops_buf2out_read_0_ranges_2),
		.loops_buf2out_read_0_ranges_3(tb_only_loops_buf2out_read_0_ranges_3),
		.loops_buf2out_read_0_ranges_4(tb_only_loops_buf2out_read_0_ranges_4),
		.loops_buf2out_read_0_ranges_5(tb_only_loops_buf2out_read_0_ranges_5),
		.loops_buf2out_read_1_dimensionality(tb_only_loops_buf2out_read_1_dimensionality),
		.loops_buf2out_read_1_ranges_0(tb_only_loops_buf2out_read_1_ranges_0),
		.loops_buf2out_read_1_ranges_1(tb_only_loops_buf2out_read_1_ranges_1),
		.loops_buf2out_read_1_ranges_2(tb_only_loops_buf2out_read_1_ranges_2),
		.loops_buf2out_read_1_ranges_3(tb_only_loops_buf2out_read_1_ranges_3),
		.loops_buf2out_read_1_ranges_4(tb_only_loops_buf2out_read_1_ranges_4),
		.loops_buf2out_read_1_ranges_5(tb_only_loops_buf2out_read_1_ranges_5),
		.loops_sram2tb_mux_sel(sram_tb_shared_loops_sram2tb_mux_sel),
		.loops_sram2tb_restart(sram_tb_shared_loops_sram2tb_restart),
		.rst_n(rst_n),
		.shared_tb_0(tb_only_shared_tb_0),
		.sram_read_data(data_from_strg),
		.t_read(sram_tb_shared_t_read_out),
		.tb_read_addr_gen_0_starting_addr(tb_only_tb_read_addr_gen_0_starting_addr),
		.tb_read_addr_gen_0_strides_0(tb_only_tb_read_addr_gen_0_strides_0),
		.tb_read_addr_gen_0_strides_1(tb_only_tb_read_addr_gen_0_strides_1),
		.tb_read_addr_gen_0_strides_2(tb_only_tb_read_addr_gen_0_strides_2),
		.tb_read_addr_gen_0_strides_3(tb_only_tb_read_addr_gen_0_strides_3),
		.tb_read_addr_gen_0_strides_4(tb_only_tb_read_addr_gen_0_strides_4),
		.tb_read_addr_gen_0_strides_5(tb_only_tb_read_addr_gen_0_strides_5),
		.tb_read_addr_gen_1_starting_addr(tb_only_tb_read_addr_gen_1_starting_addr),
		.tb_read_addr_gen_1_strides_0(tb_only_tb_read_addr_gen_1_strides_0),
		.tb_read_addr_gen_1_strides_1(tb_only_tb_read_addr_gen_1_strides_1),
		.tb_read_addr_gen_1_strides_2(tb_only_tb_read_addr_gen_1_strides_2),
		.tb_read_addr_gen_1_strides_3(tb_only_tb_read_addr_gen_1_strides_3),
		.tb_read_addr_gen_1_strides_4(tb_only_tb_read_addr_gen_1_strides_4),
		.tb_read_addr_gen_1_strides_5(tb_only_tb_read_addr_gen_1_strides_5),
		.tb_read_sched_gen_0_enable(tb_only_tb_read_sched_gen_0_enable),
		.tb_read_sched_gen_0_sched_addr_gen_delay(tb_only_tb_read_sched_gen_0_sched_addr_gen_delay),
		.tb_read_sched_gen_0_sched_addr_gen_starting_addr(tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr),
		.tb_read_sched_gen_0_sched_addr_gen_strides_0(tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0),
		.tb_read_sched_gen_0_sched_addr_gen_strides_1(tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1),
		.tb_read_sched_gen_0_sched_addr_gen_strides_2(tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2),
		.tb_read_sched_gen_0_sched_addr_gen_strides_3(tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3),
		.tb_read_sched_gen_0_sched_addr_gen_strides_4(tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4),
		.tb_read_sched_gen_0_sched_addr_gen_strides_5(tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5),
		.tb_read_sched_gen_1_enable(tb_only_tb_read_sched_gen_1_enable),
		.tb_read_sched_gen_1_sched_addr_gen_delay(tb_only_tb_read_sched_gen_1_sched_addr_gen_delay),
		.tb_read_sched_gen_1_sched_addr_gen_starting_addr(tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr),
		.tb_read_sched_gen_1_sched_addr_gen_strides_0(tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0),
		.tb_read_sched_gen_1_sched_addr_gen_strides_1(tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1),
		.tb_read_sched_gen_1_sched_addr_gen_strides_2(tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2),
		.tb_read_sched_gen_1_sched_addr_gen_strides_3(tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3),
		.tb_read_sched_gen_1_sched_addr_gen_strides_4(tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4),
		.tb_read_sched_gen_1_sched_addr_gen_strides_5(tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5),
		.tb_write_addr_gen_0_starting_addr(tb_only_tb_write_addr_gen_0_starting_addr),
		.tb_write_addr_gen_0_strides_0(tb_only_tb_write_addr_gen_0_strides_0),
		.tb_write_addr_gen_0_strides_1(tb_only_tb_write_addr_gen_0_strides_1),
		.tb_write_addr_gen_0_strides_2(tb_only_tb_write_addr_gen_0_strides_2),
		.tb_write_addr_gen_0_strides_3(tb_only_tb_write_addr_gen_0_strides_3),
		.tb_write_addr_gen_0_strides_4(tb_only_tb_write_addr_gen_0_strides_4),
		.tb_write_addr_gen_0_strides_5(tb_only_tb_write_addr_gen_0_strides_5),
		.tb_write_addr_gen_1_starting_addr(tb_only_tb_write_addr_gen_1_starting_addr),
		.tb_write_addr_gen_1_strides_0(tb_only_tb_write_addr_gen_1_strides_0),
		.tb_write_addr_gen_1_strides_1(tb_only_tb_write_addr_gen_1_strides_1),
		.tb_write_addr_gen_1_strides_2(tb_only_tb_write_addr_gen_1_strides_2),
		.tb_write_addr_gen_1_strides_3(tb_only_tb_write_addr_gen_1_strides_3),
		.tb_write_addr_gen_1_strides_4(tb_only_tb_write_addr_gen_1_strides_4),
		.tb_write_addr_gen_1_strides_5(tb_only_tb_write_addr_gen_1_strides_5),
		.accessor_output(accessor_output_int),
		.data_out(data_out_int),
		.tb_read_addr_d_out(agg_only_tb_read_addr_d_in),
		.tb_read_d_out(agg_only_tb_read_d_in)
	);
	Chain_2_16 chain(
		.accessor_output(accessor_output_int),
		.chain_data_in(chain_data_in_thin),
		.chain_en(chain_chain_en),
		.clk_en(clk_en),
		.curr_tile_data_out(data_out_int),
		.flush(flush),
		.data_out_tile(data_out_int_thin)
	);
endmodule
module strg_ub_vec_flat (
	chain_data_in_f_0,
	chain_data_in_f_1,
	clk,
	clk_en,
	data_in_f_0,
	data_in_f_1,
	flush,
	rst_n,
	strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr,
	strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0,
	strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1,
	strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2,
	strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr,
	strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0,
	strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1,
	strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2,
	strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable,
	strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr,
	strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0,
	strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1,
	strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2,
	strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable,
	strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr,
	strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0,
	strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1,
	strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2,
	strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality,
	strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0,
	strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1,
	strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2,
	strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality,
	strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0,
	strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1,
	strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2,
	strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_agg_read_padding,
	strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_agg_read_padding,
	strg_ub_vec_inst_agg_sram_shared_agg_sram_shared_addr_gen_0_starting_addr,
	strg_ub_vec_inst_agg_sram_shared_agg_sram_shared_addr_gen_1_starting_addr,
	strg_ub_vec_inst_agg_sram_shared_mode_0,
	strg_ub_vec_inst_agg_sram_shared_mode_1,
	strg_ub_vec_inst_chain_chain_en,
	strg_ub_vec_inst_data_from_strg_lifted,
	strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr,
	strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0,
	strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1,
	strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2,
	strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3,
	strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4,
	strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5,
	strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr,
	strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0,
	strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1,
	strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2,
	strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3,
	strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4,
	strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5,
	strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality,
	strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0,
	strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1,
	strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2,
	strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3,
	strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4,
	strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5,
	strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality,
	strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0,
	strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1,
	strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2,
	strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3,
	strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4,
	strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5,
	strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable,
	strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_delay,
	strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr,
	strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0,
	strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1,
	strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2,
	strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3,
	strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4,
	strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5,
	strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable,
	strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_delay,
	strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr,
	strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0,
	strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1,
	strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2,
	strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3,
	strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4,
	strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5,
	strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality,
	strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0,
	strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1,
	strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2,
	strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3,
	strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4,
	strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5,
	strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality,
	strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0,
	strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1,
	strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2,
	strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3,
	strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4,
	strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5,
	strg_ub_vec_inst_tb_only_shared_tb_0,
	strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr,
	strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0,
	strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1,
	strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2,
	strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3,
	strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4,
	strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5,
	strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr,
	strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0,
	strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1,
	strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2,
	strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3,
	strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4,
	strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5,
	strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable,
	strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_delay,
	strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr,
	strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0,
	strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1,
	strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2,
	strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3,
	strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4,
	strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5,
	strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable,
	strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_delay,
	strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr,
	strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0,
	strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1,
	strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2,
	strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3,
	strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4,
	strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5,
	strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr,
	strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0,
	strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1,
	strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2,
	strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3,
	strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4,
	strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5,
	strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr,
	strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0,
	strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1,
	strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2,
	strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3,
	strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4,
	strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5,
	accessor_output_f_b_0,
	accessor_output_f_b_1,
	data_out_f_0,
	data_out_f_1,
	strg_ub_vec_inst_addr_out_lifted,
	strg_ub_vec_inst_data_to_strg_lifted,
	strg_ub_vec_inst_ren_to_strg_lifted,
	strg_ub_vec_inst_wen_to_strg_lifted
);
	input wire [16:0] chain_data_in_f_0;
	input wire [16:0] chain_data_in_f_1;
	input wire clk;
	input wire clk_en;
	input wire [16:0] data_in_f_0;
	input wire [16:0] data_in_f_1;
	input wire flush;
	input wire rst_n;
	input wire [2:0] strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr;
	input wire [2:0] strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0;
	input wire [2:0] strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1;
	input wire [2:0] strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2;
	input wire [2:0] strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr;
	input wire [2:0] strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0;
	input wire [2:0] strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1;
	input wire [2:0] strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2;
	input wire strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable;
	input wire [15:0] strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr;
	input wire [15:0] strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0;
	input wire [15:0] strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1;
	input wire [15:0] strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2;
	input wire strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable;
	input wire [15:0] strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr;
	input wire [15:0] strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0;
	input wire [15:0] strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1;
	input wire [15:0] strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2;
	input wire [2:0] strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality;
	input wire [10:0] strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0;
	input wire [10:0] strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1;
	input wire [10:0] strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2;
	input wire [2:0] strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality;
	input wire [10:0] strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0;
	input wire [10:0] strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1;
	input wire [10:0] strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2;
	input wire [7:0] strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_agg_read_padding;
	input wire [7:0] strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_agg_read_padding;
	input wire [8:0] strg_ub_vec_inst_agg_sram_shared_agg_sram_shared_addr_gen_0_starting_addr;
	input wire [8:0] strg_ub_vec_inst_agg_sram_shared_agg_sram_shared_addr_gen_1_starting_addr;
	input wire [1:0] strg_ub_vec_inst_agg_sram_shared_mode_0;
	input wire [1:0] strg_ub_vec_inst_agg_sram_shared_mode_1;
	input wire strg_ub_vec_inst_chain_chain_en;
	input wire [63:0] strg_ub_vec_inst_data_from_strg_lifted;
	input wire [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr;
	input wire [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0;
	input wire [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1;
	input wire [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2;
	input wire [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3;
	input wire [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4;
	input wire [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5;
	input wire [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr;
	input wire [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0;
	input wire [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1;
	input wire [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2;
	input wire [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3;
	input wire [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4;
	input wire [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5;
	input wire [3:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality;
	input wire [10:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0;
	input wire [10:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1;
	input wire [10:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2;
	input wire [10:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3;
	input wire [10:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4;
	input wire [10:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5;
	input wire [3:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality;
	input wire [10:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0;
	input wire [10:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1;
	input wire [10:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2;
	input wire [10:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3;
	input wire [10:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4;
	input wire [10:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5;
	input wire strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable;
	input wire [9:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_delay;
	input wire [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr;
	input wire [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0;
	input wire [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1;
	input wire [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2;
	input wire [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3;
	input wire [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4;
	input wire [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5;
	input wire strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable;
	input wire [9:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_delay;
	input wire [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr;
	input wire [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0;
	input wire [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1;
	input wire [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2;
	input wire [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3;
	input wire [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4;
	input wire [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5;
	input wire [3:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality;
	input wire [10:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0;
	input wire [10:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1;
	input wire [10:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2;
	input wire [10:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3;
	input wire [10:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4;
	input wire [10:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5;
	input wire [3:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality;
	input wire [10:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0;
	input wire [10:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1;
	input wire [10:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2;
	input wire [10:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3;
	input wire [10:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4;
	input wire [10:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5;
	input wire strg_ub_vec_inst_tb_only_shared_tb_0;
	input wire [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr;
	input wire [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0;
	input wire [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1;
	input wire [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2;
	input wire [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3;
	input wire [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4;
	input wire [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5;
	input wire [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr;
	input wire [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0;
	input wire [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1;
	input wire [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2;
	input wire [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3;
	input wire [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4;
	input wire [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5;
	input wire strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable;
	input wire [9:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_delay;
	input wire [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr;
	input wire [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0;
	input wire [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1;
	input wire [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2;
	input wire [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3;
	input wire [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4;
	input wire [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5;
	input wire strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable;
	input wire [9:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_delay;
	input wire [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr;
	input wire [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0;
	input wire [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1;
	input wire [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2;
	input wire [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3;
	input wire [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4;
	input wire [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5;
	input wire [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr;
	input wire [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0;
	input wire [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1;
	input wire [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2;
	input wire [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3;
	input wire [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4;
	input wire [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5;
	input wire [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr;
	input wire [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0;
	input wire [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1;
	input wire [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2;
	input wire [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3;
	input wire [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4;
	input wire [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5;
	output wire accessor_output_f_b_0;
	output wire accessor_output_f_b_1;
	output wire [16:0] data_out_f_0;
	output wire [16:0] data_out_f_1;
	output wire [8:0] strg_ub_vec_inst_addr_out_lifted;
	output wire [63:0] strg_ub_vec_inst_data_to_strg_lifted;
	output wire strg_ub_vec_inst_ren_to_strg_lifted;
	output wire strg_ub_vec_inst_wen_to_strg_lifted;
	wire [1:0] strg_ub_vec_inst_accessor_output;
	wire [33:0] strg_ub_vec_inst_chain_data_in;
	wire [33:0] strg_ub_vec_inst_data_in;
	wire [33:0] strg_ub_vec_inst_data_out;
	assign strg_ub_vec_inst_data_in[0+:17] = data_in_f_0;
	assign strg_ub_vec_inst_data_in[17+:17] = data_in_f_1;
	assign strg_ub_vec_inst_chain_data_in[0+:17] = chain_data_in_f_0;
	assign strg_ub_vec_inst_chain_data_in[17+:17] = chain_data_in_f_1;
	assign data_out_f_0 = strg_ub_vec_inst_data_out[0+:17];
	assign data_out_f_1 = strg_ub_vec_inst_data_out[17+:17];
	assign accessor_output_f_b_0 = strg_ub_vec_inst_accessor_output[0];
	assign accessor_output_f_b_1 = strg_ub_vec_inst_accessor_output[1];
	strg_ub_vec strg_ub_vec_inst(
		.agg_only_agg_write_addr_gen_0_starting_addr(strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr),
		.agg_only_agg_write_addr_gen_0_strides_0(strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0),
		.agg_only_agg_write_addr_gen_0_strides_1(strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1),
		.agg_only_agg_write_addr_gen_0_strides_2(strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2),
		.agg_only_agg_write_addr_gen_1_starting_addr(strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr),
		.agg_only_agg_write_addr_gen_1_strides_0(strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0),
		.agg_only_agg_write_addr_gen_1_strides_1(strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1),
		.agg_only_agg_write_addr_gen_1_strides_2(strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2),
		.agg_only_agg_write_sched_gen_0_enable(strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable),
		.agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr(strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr),
		.agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0(strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0),
		.agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1(strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1),
		.agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2(strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2),
		.agg_only_agg_write_sched_gen_1_enable(strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable),
		.agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr(strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr),
		.agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0(strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0),
		.agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1(strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1),
		.agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2(strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2),
		.agg_only_loops_in2buf_0_dimensionality(strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality),
		.agg_only_loops_in2buf_0_ranges_0(strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0),
		.agg_only_loops_in2buf_0_ranges_1(strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1),
		.agg_only_loops_in2buf_0_ranges_2(strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2),
		.agg_only_loops_in2buf_1_dimensionality(strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality),
		.agg_only_loops_in2buf_1_ranges_0(strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0),
		.agg_only_loops_in2buf_1_ranges_1(strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1),
		.agg_only_loops_in2buf_1_ranges_2(strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2),
		.agg_sram_shared_agg_read_sched_gen_0_agg_read_padding(strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_agg_read_padding),
		.agg_sram_shared_agg_read_sched_gen_1_agg_read_padding(strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_agg_read_padding),
		.agg_sram_shared_agg_sram_shared_addr_gen_0_starting_addr(strg_ub_vec_inst_agg_sram_shared_agg_sram_shared_addr_gen_0_starting_addr),
		.agg_sram_shared_agg_sram_shared_addr_gen_1_starting_addr(strg_ub_vec_inst_agg_sram_shared_agg_sram_shared_addr_gen_1_starting_addr),
		.agg_sram_shared_mode_0(strg_ub_vec_inst_agg_sram_shared_mode_0),
		.agg_sram_shared_mode_1(strg_ub_vec_inst_agg_sram_shared_mode_1),
		.chain_chain_en(strg_ub_vec_inst_chain_chain_en),
		.chain_data_in(strg_ub_vec_inst_chain_data_in),
		.clk(clk),
		.clk_en(clk_en),
		.data_from_strg(strg_ub_vec_inst_data_from_strg_lifted),
		.data_in(strg_ub_vec_inst_data_in),
		.flush(flush),
		.rst_n(rst_n),
		.sram_only_output_addr_gen_0_starting_addr(strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr),
		.sram_only_output_addr_gen_0_strides_0(strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0),
		.sram_only_output_addr_gen_0_strides_1(strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1),
		.sram_only_output_addr_gen_0_strides_2(strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2),
		.sram_only_output_addr_gen_0_strides_3(strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3),
		.sram_only_output_addr_gen_0_strides_4(strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4),
		.sram_only_output_addr_gen_0_strides_5(strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5),
		.sram_only_output_addr_gen_1_starting_addr(strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr),
		.sram_only_output_addr_gen_1_strides_0(strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0),
		.sram_only_output_addr_gen_1_strides_1(strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1),
		.sram_only_output_addr_gen_1_strides_2(strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2),
		.sram_only_output_addr_gen_1_strides_3(strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3),
		.sram_only_output_addr_gen_1_strides_4(strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4),
		.sram_only_output_addr_gen_1_strides_5(strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5),
		.sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality),
		.sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0),
		.sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1),
		.sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2),
		.sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3),
		.sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4),
		.sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5),
		.sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality),
		.sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0),
		.sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1),
		.sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2),
		.sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3),
		.sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4),
		.sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5),
		.sram_tb_shared_output_sched_gen_0_enable(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable),
		.sram_tb_shared_output_sched_gen_0_sched_addr_gen_delay(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_delay),
		.sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr),
		.sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0),
		.sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1),
		.sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2),
		.sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3),
		.sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4),
		.sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5),
		.sram_tb_shared_output_sched_gen_1_enable(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable),
		.sram_tb_shared_output_sched_gen_1_sched_addr_gen_delay(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_delay),
		.sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr),
		.sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0),
		.sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1),
		.sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2),
		.sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3),
		.sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4),
		.sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5),
		.tb_only_loops_buf2out_read_0_dimensionality(strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality),
		.tb_only_loops_buf2out_read_0_ranges_0(strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0),
		.tb_only_loops_buf2out_read_0_ranges_1(strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1),
		.tb_only_loops_buf2out_read_0_ranges_2(strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2),
		.tb_only_loops_buf2out_read_0_ranges_3(strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3),
		.tb_only_loops_buf2out_read_0_ranges_4(strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4),
		.tb_only_loops_buf2out_read_0_ranges_5(strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5),
		.tb_only_loops_buf2out_read_1_dimensionality(strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality),
		.tb_only_loops_buf2out_read_1_ranges_0(strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0),
		.tb_only_loops_buf2out_read_1_ranges_1(strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1),
		.tb_only_loops_buf2out_read_1_ranges_2(strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2),
		.tb_only_loops_buf2out_read_1_ranges_3(strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3),
		.tb_only_loops_buf2out_read_1_ranges_4(strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4),
		.tb_only_loops_buf2out_read_1_ranges_5(strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5),
		.tb_only_shared_tb_0(strg_ub_vec_inst_tb_only_shared_tb_0),
		.tb_only_tb_read_addr_gen_0_starting_addr(strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr),
		.tb_only_tb_read_addr_gen_0_strides_0(strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0),
		.tb_only_tb_read_addr_gen_0_strides_1(strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1),
		.tb_only_tb_read_addr_gen_0_strides_2(strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2),
		.tb_only_tb_read_addr_gen_0_strides_3(strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3),
		.tb_only_tb_read_addr_gen_0_strides_4(strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4),
		.tb_only_tb_read_addr_gen_0_strides_5(strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5),
		.tb_only_tb_read_addr_gen_1_starting_addr(strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr),
		.tb_only_tb_read_addr_gen_1_strides_0(strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0),
		.tb_only_tb_read_addr_gen_1_strides_1(strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1),
		.tb_only_tb_read_addr_gen_1_strides_2(strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2),
		.tb_only_tb_read_addr_gen_1_strides_3(strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3),
		.tb_only_tb_read_addr_gen_1_strides_4(strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4),
		.tb_only_tb_read_addr_gen_1_strides_5(strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5),
		.tb_only_tb_read_sched_gen_0_enable(strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable),
		.tb_only_tb_read_sched_gen_0_sched_addr_gen_delay(strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_delay),
		.tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr(strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr),
		.tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0(strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0),
		.tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1(strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1),
		.tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2(strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2),
		.tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3(strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3),
		.tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4(strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4),
		.tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5(strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5),
		.tb_only_tb_read_sched_gen_1_enable(strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable),
		.tb_only_tb_read_sched_gen_1_sched_addr_gen_delay(strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_delay),
		.tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr(strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr),
		.tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0(strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0),
		.tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1(strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1),
		.tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2(strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2),
		.tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3(strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3),
		.tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4(strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4),
		.tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5(strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5),
		.tb_only_tb_write_addr_gen_0_starting_addr(strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr),
		.tb_only_tb_write_addr_gen_0_strides_0(strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0),
		.tb_only_tb_write_addr_gen_0_strides_1(strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1),
		.tb_only_tb_write_addr_gen_0_strides_2(strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2),
		.tb_only_tb_write_addr_gen_0_strides_3(strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3),
		.tb_only_tb_write_addr_gen_0_strides_4(strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4),
		.tb_only_tb_write_addr_gen_0_strides_5(strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5),
		.tb_only_tb_write_addr_gen_1_starting_addr(strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr),
		.tb_only_tb_write_addr_gen_1_strides_0(strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0),
		.tb_only_tb_write_addr_gen_1_strides_1(strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1),
		.tb_only_tb_write_addr_gen_1_strides_2(strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2),
		.tb_only_tb_write_addr_gen_1_strides_3(strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3),
		.tb_only_tb_write_addr_gen_1_strides_4(strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4),
		.tb_only_tb_write_addr_gen_1_strides_5(strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5),
		.accessor_output(strg_ub_vec_inst_accessor_output),
		.addr_out(strg_ub_vec_inst_addr_out_lifted),
		.data_out(strg_ub_vec_inst_data_out),
		.data_to_strg(strg_ub_vec_inst_data_to_strg_lifted),
		.ren_to_strg(strg_ub_vec_inst_ren_to_strg_lifted),
		.wen_to_strg(strg_ub_vec_inst_wen_to_strg_lifted)
	);
endmodule
module write_scanner (
	ID_out_ready,
	addr_in,
	addr_in_valid,
	addr_out_ready,
	block_mode,
	block_wr_in,
	block_wr_in_valid,
	clk,
	clk_en,
	compressed,
	data_in,
	data_in_valid,
	data_out_ready,
	flush,
	init_blank,
	lowest_level,
	rst_n,
	spacc_mode,
	stop_lvl,
	tile_en,
	ID_out,
	ID_out_valid,
	addr_in_ready,
	addr_out,
	addr_out_valid,
	block_wr_in_ready,
	data_in_ready,
	data_out,
	data_out_valid
);
	input wire ID_out_ready;
	input wire [16:0] addr_in;
	input wire addr_in_valid;
	input wire addr_out_ready;
	input wire block_mode;
	input wire [16:0] block_wr_in;
	input wire block_wr_in_valid;
	input wire clk;
	input wire clk_en;
	input wire compressed;
	input wire [16:0] data_in;
	input wire data_in_valid;
	input wire data_out_ready;
	input wire flush;
	input wire init_blank;
	input wire lowest_level;
	input wire rst_n;
	input wire spacc_mode;
	input wire [15:0] stop_lvl;
	input wire tile_en;
	output wire [16:0] ID_out;
	output wire ID_out_valid;
	output wire addr_in_ready;
	output wire [16:0] addr_out;
	output wire addr_out_valid;
	output wire block_wr_in_ready;
	output wire data_in_ready;
	output wire [16:0] data_out;
	output wire data_out_valid;
	wire [16:0] ID_out_fifo_data_in;
	wire ID_out_fifo_empty;
	wire ID_out_fifo_full;
	wire ID_out_fifo_push;
	reg [15:0] ID_to_fifo;
	reg IN_DONE;
	wire addr_done_in;
	wire [15:0] addr_infifo_data_in;
	wire addr_infifo_eos_in;
	wire [16:0] addr_infifo_in_packed;
	wire [16:0] addr_infifo_out_packed;
	wire addr_infifo_valid_in;
	wire addr_input_fifo_empty;
	wire addr_input_fifo_full;
	wire [16:0] addr_out_fifo_data_in;
	wire addr_out_fifo_empty;
	wire addr_out_fifo_full;
	wire addr_out_fifo_push;
	reg [15:0] addr_to_fifo;
	wire blank_done_stick_sticky;
	reg blank_done_stick_was_high;
	reg [15:0] block_size;
	wire block_wr_fifo_valid;
	wire [15:0] block_wr_input_fifo_data_out;
	wire block_wr_input_fifo_empty;
	wire block_wr_input_fifo_full;
	reg [15:0] block_write_count;
	reg clr_blank_done;
	reg clr_block_write;
	reg clr_coord_addr;
	reg clr_curr_coord;
	reg clr_seg_addr;
	reg clr_seg_ctr;
	reg clr_wen_made;
	reg [15:0] coord_addr;
	wire data_done_in;
	wire [15:0] data_infifo_data_in;
	reg [15:0] data_infifo_data_in_d1;
	wire data_infifo_eos_in;
	wire [16:0] data_infifo_in_packed;
	wire [16:0] data_infifo_out_packed;
	wire data_infifo_valid_in;
	wire data_input_fifo_empty;
	wire data_input_fifo_full;
	wire [16:0] data_out_fifo_data_in;
	wire data_out_fifo_empty;
	wire data_out_fifo_full;
	wire data_out_fifo_push;
	reg [15:0] data_to_fifo;
	wire gclk;
	reg inc_block_write;
	reg inc_coord_addr;
	reg inc_seg_addr;
	reg inc_seg_ctr;
	reg [1:0] infifo_pop;
	wire matching_stop;
	wire new_coord;
	reg op_to_fifo;
	reg pop_block_wr;
	reg push_to_outs;
	reg [4:0] scan_seq_current_state;
	reg [4:0] scan_seq_next_state;
	reg [15:0] segment_addr;
	reg [15:0] segment_counter;
	reg set_blank_done;
	reg set_block_size;
	reg set_curr_coord;
	wire stop_in;
	wire stop_lvl_geq;
	wire stop_lvl_geq_p1;
	wire stop_lvl_new_blank_sticky_sticky;
	reg stop_lvl_new_blank_sticky_was_high;
	wire valid_coord_sticky_sticky;
	reg valid_coord_sticky_was_high;
	wire wen_made_sticky;
	reg wen_made_was_high;
	assign gclk = clk & tile_en;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			blank_done_stick_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				blank_done_stick_was_high <= 1'h0;
			else if (clr_blank_done)
				blank_done_stick_was_high <= 1'h0;
			else if (set_blank_done)
				blank_done_stick_was_high <= 1'h1;
		end
	assign blank_done_stick_sticky = blank_done_stick_was_high;
	assign data_infifo_in_packed[16] = data_in[16];
	assign data_infifo_in_packed[15:0] = data_in[15:0];
	assign data_infifo_eos_in = data_infifo_out_packed[16];
	assign data_infifo_data_in = data_infifo_out_packed[15:0];
	assign data_in_ready = ~data_input_fifo_full;
	assign data_infifo_valid_in = ~data_input_fifo_empty;
	assign addr_infifo_in_packed[16] = addr_in[16];
	assign addr_infifo_in_packed[15:0] = addr_in[15:0];
	assign addr_infifo_eos_in = addr_infifo_out_packed[16];
	assign addr_infifo_data_in = addr_infifo_out_packed[15:0];
	assign addr_in_ready = ~addr_input_fifo_full;
	assign addr_infifo_valid_in = ~addr_input_fifo_empty;
	assign block_wr_in_ready = ~block_wr_input_fifo_full;
	assign block_wr_fifo_valid = ~block_wr_input_fifo_empty;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			block_size <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				block_size <= 16'h0000;
			else if (set_block_size)
				block_size <= block_wr_input_fifo_data_out;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			block_write_count <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				block_write_count <= 16'h0000;
			else if (clr_block_write)
				block_write_count <= 16'h0000;
			else if (inc_block_write)
				block_write_count <= block_write_count + 16'h0001;
		end
	assign data_out_fifo_data_in = {op_to_fifo, data_to_fifo};
	assign data_out_valid = ~data_out_fifo_empty;
	assign addr_out_fifo_data_in = {1'h0, addr_to_fifo};
	assign addr_out_valid = ~addr_out_fifo_empty;
	assign ID_out_fifo_data_in = {1'h0, ID_to_fifo};
	assign ID_out_valid = ~ID_out_fifo_empty;
	assign {data_out_fifo_push, addr_out_fifo_push, ID_out_fifo_push} = {push_to_outs, push_to_outs, push_to_outs};
	assign stop_lvl_geq = ((data_infifo_eos_in & data_infifo_valid_in) & (data_infifo_data_in[9:8] == 2'h0)) & (data_infifo_data_in[7:0] >= stop_lvl[7:0]);
	assign stop_lvl_geq_p1 = ((data_infifo_eos_in & data_infifo_valid_in) & (data_infifo_data_in[9:8] == 2'h0)) & (data_infifo_data_in[7:0] >= (stop_lvl[7:0] + 8'h01));
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			stop_lvl_new_blank_sticky_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				stop_lvl_new_blank_sticky_was_high <= 1'h0;
			else if (clr_blank_done)
				stop_lvl_new_blank_sticky_was_high <= 1'h0;
			else if (stop_lvl_geq_p1)
				stop_lvl_new_blank_sticky_was_high <= 1'h1;
		end
	assign stop_lvl_new_blank_sticky_sticky = stop_lvl_new_blank_sticky_was_high;
	assign data_done_in = (data_infifo_valid_in & data_infifo_eos_in) & (data_infifo_data_in[9:8] == 2'h1);
	assign addr_done_in = (addr_infifo_valid_in & addr_infifo_eos_in) & (addr_infifo_data_in[9:8] == 2'h1);
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			segment_addr <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				segment_addr <= 16'h0000;
			else if (clr_seg_addr)
				segment_addr <= 16'h0000;
			else if (inc_seg_addr)
				segment_addr <= segment_addr + 16'h0001;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			coord_addr <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				coord_addr <= 16'h0000;
			else if (clr_coord_addr)
				coord_addr <= 16'h0000;
			else if (inc_coord_addr)
				coord_addr <= coord_addr + 16'h0001;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			segment_counter <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				segment_counter <= 16'h0000;
			else if (clr_seg_ctr)
				segment_counter <= 16'h0000;
			else if (inc_seg_ctr)
				segment_counter <= segment_counter + 16'h0001;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			data_infifo_data_in_d1 <= 16'h0000;
		else if (clk_en) begin
			if (flush)
				data_infifo_data_in_d1 <= 16'h0000;
			else if (set_curr_coord)
				data_infifo_data_in_d1 <= data_infifo_data_in;
		end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			valid_coord_sticky_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				valid_coord_sticky_was_high <= 1'h0;
			else if (clr_curr_coord)
				valid_coord_sticky_was_high <= 1'h0;
			else if (set_curr_coord)
				valid_coord_sticky_was_high <= 1'h1;
		end
	assign valid_coord_sticky_sticky = valid_coord_sticky_was_high;
	assign new_coord = (data_infifo_valid_in & ~data_infifo_eos_in) & (~valid_coord_sticky_sticky | (data_infifo_data_in != data_infifo_data_in_d1));
	assign stop_in = data_infifo_valid_in & data_infifo_eos_in;
	assign matching_stop = data_infifo_valid_in & data_infifo_eos_in;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			wen_made_was_high <= 1'h0;
		else if (clk_en) begin
			if (flush)
				wen_made_was_high <= 1'h0;
			else if (clr_wen_made)
				wen_made_was_high <= 1'h0;
			else if (push_to_outs)
				wen_made_was_high <= 1'h1;
		end
	assign wen_made_sticky = wen_made_was_high;
	always @(posedge clk or negedge rst_n)
		if (!rst_n)
			scan_seq_current_state <= 5'h0b;
		else if (clk_en) begin
			if (flush)
				scan_seq_current_state <= 5'h0b;
			else
				scan_seq_current_state <= scan_seq_next_state;
		end
	always @(*) begin
		scan_seq_next_state = scan_seq_current_state;
		case (scan_seq_current_state)
			5'h00:
				if (~(&(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full})))
					scan_seq_next_state = 5'h00;
				else if (~lowest_level & &(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full}))
					scan_seq_next_state = 5'h01;
				else if ((lowest_level & block_mode) & &(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full}))
					scan_seq_next_state = 5'h02;
				else if ((lowest_level & ~block_mode) & &(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full}))
					scan_seq_next_state = 5'h0a;
			5'h01:
				if (~(&(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full})))
					scan_seq_next_state = 5'h01;
				else if (block_mode & &(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full}))
					scan_seq_next_state = 5'h02;
				else if (~block_mode & &(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full}))
					scan_seq_next_state = 5'h0f;
			5'h02:
				if (block_wr_fifo_valid)
					scan_seq_next_state = 5'h03;
				else
					scan_seq_next_state = 5'h02;
			5'h03:
				if ((block_write_count == block_size) & ~lowest_level)
					scan_seq_next_state = 5'h04;
				else if ((block_write_count == block_size) & lowest_level)
					scan_seq_next_state = 5'h09;
				else
					scan_seq_next_state = 5'h03;
			5'h04:
				if (block_wr_fifo_valid)
					scan_seq_next_state = 5'h05;
				else
					scan_seq_next_state = 5'h04;
			5'h05:
				if (block_write_count == block_size)
					scan_seq_next_state = 5'h08;
				else
					scan_seq_next_state = 5'h05;
			5'h06:
				if (data_done_in | (spacc_mode & stop_lvl_geq))
					scan_seq_next_state = 5'h09;
				else
					scan_seq_next_state = 5'h06;
			5'h07: scan_seq_next_state = 5'h0b;
			5'h08:
				if (&(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full}))
					scan_seq_next_state = 5'h09;
				else
					scan_seq_next_state = 5'h08;
			5'h09:
				if (&(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full}))
					scan_seq_next_state = 5'h07;
				else
					scan_seq_next_state = 5'h09;
			5'h0a:
				if (init_blank & ~blank_done_stick_sticky)
					scan_seq_next_state = 5'h09;
				else if (compressed & (~init_blank | blank_done_stick_sticky))
					scan_seq_next_state = 5'h06;
				else if (~compressed & (~init_blank | blank_done_stick_sticky))
					scan_seq_next_state = 5'h10;
			5'h0b:
				if (tile_en)
					scan_seq_next_state = 5'h00;
				else
					scan_seq_next_state = 5'h0b;
			5'h0c:
				if (new_coord)
					scan_seq_next_state = 5'h0d;
				else if (matching_stop | (init_blank & ~blank_done_stick_sticky))
					scan_seq_next_state = 5'h0e;
				else
					scan_seq_next_state = 5'h0c;
			5'h0d:
				if (new_coord | stop_in)
					scan_seq_next_state = 5'h0c;
				else
					scan_seq_next_state = 5'h0d;
			5'h0e:
				if ((init_blank ? (data_infifo_valid_in & ~data_infifo_eos_in) & blank_done_stick_sticky : data_infifo_valid_in & ~data_infifo_eos_in))
					scan_seq_next_state = 5'h0c;
				else if ((spacc_mode ? (data_done_in | (init_blank & ~blank_done_stick_sticky)) | stop_lvl_geq : data_done_in))
					scan_seq_next_state = 5'h08;
				else
					scan_seq_next_state = 5'h0e;
			5'h0f:
				if (&(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full}))
					scan_seq_next_state = 5'h0c;
				else if (~(&(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full})))
					scan_seq_next_state = 5'h0f;
			5'h10:
				if ((data_done_in & addr_done_in) | (spacc_mode & stop_lvl_geq))
					scan_seq_next_state = 5'h09;
				else
					scan_seq_next_state = 5'h10;
			default: scan_seq_next_state = scan_seq_current_state;
		endcase
	end
	always @(*)
		case (scan_seq_current_state)
			5'h00: begin : scan_seq_ALLOCATE1_Output
				data_to_fifo = 16'h0000;
				op_to_fifo = 1'h0;
				addr_to_fifo = 16'h0000;
				ID_to_fifo = 16'h0000;
				push_to_outs = 1'h1;
				inc_seg_addr = 1'h0;
				clr_seg_addr = 1'h0;
				inc_coord_addr = 1'h0;
				clr_coord_addr = 1'h0;
				inc_seg_ctr = 1'h0;
				clr_seg_ctr = 1'h0;
				set_curr_coord = 1'h0;
				clr_curr_coord = 1'h0;
				infifo_pop[0] = 1'h0;
				infifo_pop[1] = 1'h0;
				clr_wen_made = 1'h0;
				set_block_size = 1'h0;
				inc_block_write = 1'h0;
				clr_block_write = 1'h0;
				IN_DONE = 1'h0;
				clr_blank_done = 1'h0;
				set_blank_done = 1'h0;
				pop_block_wr = 1'h0;
			end
			5'h01: begin : scan_seq_ALLOCATE2_Output
				data_to_fifo = 16'h0000;
				op_to_fifo = 1'h0;
				addr_to_fifo = 16'h0000;
				ID_to_fifo = 16'h0001;
				push_to_outs = 1'h1;
				inc_seg_addr = 1'h0;
				clr_seg_addr = 1'h0;
				inc_coord_addr = 1'h0;
				clr_coord_addr = 1'h0;
				inc_seg_ctr = 1'h0;
				clr_seg_ctr = 1'h0;
				set_curr_coord = 1'h0;
				clr_curr_coord = 1'h0;
				infifo_pop[0] = 1'h0;
				infifo_pop[1] = 1'h0;
				clr_wen_made = 1'h0;
				set_block_size = 1'h0;
				inc_block_write = 1'h0;
				clr_block_write = 1'h0;
				IN_DONE = 1'h0;
				clr_blank_done = 1'h0;
				set_blank_done = 1'h0;
				pop_block_wr = 1'h0;
			end
			5'h02: begin : scan_seq_BLOCK_1_SZ_Output
				data_to_fifo = 16'h0000;
				op_to_fifo = 1'h0;
				addr_to_fifo = 16'h0000;
				ID_to_fifo = 16'h0001;
				push_to_outs = 1'h0;
				inc_seg_addr = 1'h0;
				clr_seg_addr = 1'h0;
				inc_coord_addr = 1'h0;
				clr_coord_addr = 1'h0;
				inc_seg_ctr = 1'h0;
				clr_seg_ctr = 1'h0;
				set_curr_coord = 1'h0;
				clr_curr_coord = 1'h0;
				infifo_pop[0] = 1'h0;
				infifo_pop[1] = 1'h0;
				clr_wen_made = 1'h0;
				set_block_size = block_wr_fifo_valid;
				inc_block_write = 1'h0;
				clr_block_write = 1'h1;
				pop_block_wr = block_wr_fifo_valid;
				IN_DONE = 1'h0;
				clr_blank_done = 1'h0;
				set_blank_done = 1'h0;
			end
			5'h03: begin : scan_seq_BLOCK_1_WR_Output
				data_to_fifo = block_wr_input_fifo_data_out;
				op_to_fifo = 1'h1;
				addr_to_fifo = block_write_count;
				ID_to_fifo = 16'h0000;
				push_to_outs = block_wr_fifo_valid & (block_write_count < block_size);
				inc_seg_addr = 1'h0;
				clr_seg_addr = 1'h0;
				inc_coord_addr = 1'h0;
				clr_coord_addr = 1'h0;
				inc_seg_ctr = 1'h0;
				clr_seg_ctr = 1'h0;
				set_curr_coord = 1'h0;
				clr_curr_coord = 1'h0;
				infifo_pop[0] = 1'h0;
				infifo_pop[1] = 1'h0;
				clr_wen_made = 1'h0;
				set_block_size = 1'h0;
				inc_block_write = (block_wr_fifo_valid & (block_write_count < block_size)) & &(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full});
				clr_block_write = 1'h0;
				pop_block_wr = (block_wr_fifo_valid & (block_write_count < block_size)) & &(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full});
				IN_DONE = 1'h0;
				clr_blank_done = 1'h0;
				set_blank_done = 1'h0;
			end
			5'h04: begin : scan_seq_BLOCK_2_SZ_Output
				data_to_fifo = 16'h0000;
				op_to_fifo = 1'h0;
				addr_to_fifo = 16'h0000;
				ID_to_fifo = 16'h0000;
				push_to_outs = 1'h0;
				inc_seg_addr = 1'h0;
				clr_seg_addr = 1'h0;
				inc_coord_addr = 1'h0;
				clr_coord_addr = 1'h0;
				inc_seg_ctr = 1'h0;
				clr_seg_ctr = 1'h0;
				set_curr_coord = 1'h0;
				clr_curr_coord = 1'h0;
				infifo_pop[0] = 1'h0;
				infifo_pop[1] = 1'h0;
				clr_wen_made = 1'h0;
				set_block_size = block_wr_fifo_valid;
				inc_block_write = 1'h0;
				clr_block_write = 1'h1;
				pop_block_wr = block_wr_fifo_valid;
				IN_DONE = 1'h0;
				clr_blank_done = 1'h0;
				set_blank_done = 1'h0;
			end
			5'h05: begin : scan_seq_BLOCK_2_WR_Output
				data_to_fifo = block_wr_input_fifo_data_out;
				op_to_fifo = 1'h1;
				addr_to_fifo = block_write_count;
				ID_to_fifo = 16'h0001;
				push_to_outs = block_wr_fifo_valid & (block_write_count < block_size);
				inc_seg_addr = 1'h0;
				clr_seg_addr = 1'h0;
				inc_coord_addr = 1'h0;
				clr_coord_addr = 1'h0;
				inc_seg_ctr = 1'h0;
				clr_seg_ctr = 1'h0;
				set_curr_coord = 1'h0;
				clr_curr_coord = 1'h0;
				infifo_pop[0] = 1'h0;
				infifo_pop[1] = 1'h0;
				clr_wen_made = 1'h0;
				set_block_size = 1'h0;
				inc_block_write = (block_wr_fifo_valid & (block_write_count < block_size)) & &(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full});
				clr_block_write = 1'h0;
				pop_block_wr = (block_wr_fifo_valid & (block_write_count < block_size)) & &(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full});
				IN_DONE = 1'h0;
				clr_blank_done = 1'h0;
				set_blank_done = 1'h0;
			end
			5'h06: begin : scan_seq_ComLL_Output
				data_to_fifo = data_infifo_data_in;
				op_to_fifo = 1'h1;
				addr_to_fifo = segment_addr;
				ID_to_fifo = 16'h0000;
				push_to_outs = data_infifo_valid_in & ~data_infifo_eos_in;
				inc_seg_addr = (data_infifo_valid_in & ~data_infifo_eos_in) & &(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full});
				clr_seg_addr = 1'h0;
				inc_coord_addr = 1'h0;
				clr_coord_addr = 1'h0;
				inc_seg_ctr = 1'h0;
				clr_seg_ctr = 1'h0;
				set_curr_coord = 1'h0;
				clr_curr_coord = 1'h0;
				infifo_pop[0] = data_infifo_valid_in & (data_infifo_eos_in | &(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full}));
				infifo_pop[1] = 1'h0;
				clr_wen_made = 1'h0;
				set_block_size = 1'h0;
				inc_block_write = 1'h0;
				clr_block_write = 1'h0;
				IN_DONE = 1'h0;
				clr_blank_done = 1'h0;
				set_blank_done = 1'h0;
				pop_block_wr = 1'h0;
			end
			5'h07: begin : scan_seq_DONE_Output
				data_to_fifo = 16'h0000;
				op_to_fifo = 1'h0;
				addr_to_fifo = 16'h0000;
				ID_to_fifo = 16'h0000;
				push_to_outs = 1'h0;
				inc_seg_addr = 1'h0;
				clr_seg_addr = 1'h0;
				inc_coord_addr = 1'h0;
				clr_coord_addr = 1'h0;
				inc_seg_ctr = 1'h0;
				clr_seg_ctr = 1'h0;
				set_curr_coord = 1'h0;
				clr_curr_coord = 1'h0;
				infifo_pop[0] = data_done_in;
				infifo_pop[1] = 1'h0;
				clr_wen_made = 1'h0;
				set_block_size = 1'h0;
				inc_block_write = 1'h0;
				clr_block_write = 1'h0;
				set_blank_done = (init_blank & ~blank_done_stick_sticky) & spacc_mode;
				clr_blank_done = ((init_blank & blank_done_stick_sticky) & stop_lvl_new_blank_sticky_sticky) & spacc_mode;
				IN_DONE = 1'h1;
				pop_block_wr = 1'h0;
			end
			5'h08: begin : scan_seq_FINALIZE1_Output
				data_to_fifo = 16'h0000;
				op_to_fifo = 1'h0;
				addr_to_fifo = 16'h0000;
				ID_to_fifo = 16'h0001;
				push_to_outs = 1'h1;
				inc_seg_addr = 1'h0;
				clr_seg_addr = 1'h0;
				inc_coord_addr = 1'h0;
				clr_coord_addr = 1'h0;
				inc_seg_ctr = 1'h0;
				clr_seg_ctr = 1'h0;
				set_curr_coord = 1'h0;
				clr_curr_coord = 1'h0;
				infifo_pop[0] = 1'h0;
				infifo_pop[1] = 1'h0;
				clr_wen_made = 1'h0;
				set_block_size = 1'h0;
				inc_block_write = 1'h0;
				clr_block_write = 1'h0;
				IN_DONE = 1'h0;
				clr_blank_done = 1'h0;
				set_blank_done = 1'h0;
				pop_block_wr = 1'h0;
			end
			5'h09: begin : scan_seq_FINALIZE2_Output
				data_to_fifo = 16'h0000;
				op_to_fifo = 1'h0;
				addr_to_fifo = 16'h0000;
				ID_to_fifo = 16'h0000;
				push_to_outs = 1'h1;
				inc_seg_addr = 1'h0;
				clr_seg_addr = 1'h0;
				inc_coord_addr = 1'h0;
				clr_coord_addr = 1'h0;
				inc_seg_ctr = 1'h0;
				clr_seg_ctr = 1'h0;
				set_curr_coord = 1'h0;
				clr_curr_coord = 1'h0;
				infifo_pop[0] = 1'h0;
				infifo_pop[1] = 1'h0;
				clr_wen_made = 1'h0;
				set_block_size = 1'h0;
				inc_block_write = 1'h0;
				clr_block_write = 1'h0;
				IN_DONE = 1'h0;
				clr_blank_done = 1'h0;
				set_blank_done = 1'h0;
				pop_block_wr = 1'h0;
			end
			5'h0a: begin : scan_seq_LL_Output
				data_to_fifo = 16'h0000;
				op_to_fifo = 1'h0;
				addr_to_fifo = 16'h0000;
				ID_to_fifo = 16'h0000;
				push_to_outs = 1'h0;
				inc_seg_addr = 1'h0;
				clr_seg_addr = 1'h0;
				inc_coord_addr = 1'h0;
				clr_coord_addr = 1'h0;
				inc_seg_ctr = 1'h0;
				clr_seg_ctr = 1'h0;
				set_curr_coord = 1'h0;
				clr_curr_coord = 1'h0;
				infifo_pop[0] = 1'h0;
				infifo_pop[1] = 1'h0;
				clr_wen_made = 1'h0;
				set_block_size = 1'h0;
				inc_block_write = 1'h0;
				clr_block_write = 1'h0;
				IN_DONE = 1'h0;
				clr_blank_done = 1'h0;
				set_blank_done = 1'h0;
				pop_block_wr = 1'h0;
			end
			5'h0b: begin : scan_seq_START_Output
				data_to_fifo = 16'h0000;
				op_to_fifo = 1'h0;
				addr_to_fifo = 16'h0000;
				ID_to_fifo = 16'h0000;
				push_to_outs = 1'h0;
				inc_seg_addr = 1'h0;
				clr_seg_addr = 1'h1;
				inc_coord_addr = 1'h0;
				clr_coord_addr = 1'h1;
				inc_seg_ctr = 1'h0;
				clr_seg_ctr = 1'h1;
				set_curr_coord = 1'h0;
				clr_curr_coord = 1'h1;
				infifo_pop[0] = 1'h0;
				infifo_pop[1] = 1'h0;
				clr_wen_made = 1'h1;
				set_block_size = 1'h0;
				inc_block_write = 1'h0;
				clr_block_write = 1'h1;
				IN_DONE = 1'h0;
				clr_blank_done = 1'h0;
				set_blank_done = 1'h0;
				pop_block_wr = 1'h0;
			end
			5'h0c: begin : scan_seq_UL_Output
				data_to_fifo = 16'h0000;
				op_to_fifo = 1'h0;
				addr_to_fifo = 16'h0000;
				ID_to_fifo = 16'h0000;
				push_to_outs = 1'h0;
				inc_seg_addr = 1'h0;
				clr_seg_addr = 1'h0;
				inc_coord_addr = 1'h0;
				clr_coord_addr = 1'h0;
				inc_seg_ctr = 1'h0;
				clr_seg_ctr = 1'h0;
				set_curr_coord = new_coord;
				clr_curr_coord = 1'h0;
				infifo_pop[0] = 1'h0;
				infifo_pop[1] = 1'h0;
				clr_wen_made = 1'h1;
				set_block_size = 1'h0;
				inc_block_write = 1'h0;
				clr_block_write = 1'h0;
				IN_DONE = 1'h0;
				clr_blank_done = 1'h0;
				set_blank_done = 1'h0;
				pop_block_wr = 1'h0;
			end
			5'h0d: begin : scan_seq_UL_EMIT_COORD_Output
				data_to_fifo = data_infifo_data_in_d1;
				op_to_fifo = 1'h1;
				addr_to_fifo = coord_addr;
				ID_to_fifo = 16'h0001;
				push_to_outs = ~wen_made_sticky & &(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full});
				inc_seg_addr = 1'h0;
				clr_seg_addr = 1'h0;
				inc_coord_addr = ~wen_made_sticky & &(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full});
				clr_coord_addr = 1'h0;
				inc_seg_ctr = ~wen_made_sticky & &(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full});
				clr_seg_ctr = 1'h0;
				set_curr_coord = 1'h0;
				clr_curr_coord = 1'h0;
				infifo_pop[0] = ~new_coord & ~stop_in;
				infifo_pop[1] = 1'h0;
				clr_wen_made = 1'h0;
				set_block_size = 1'h0;
				inc_block_write = 1'h0;
				clr_block_write = 1'h0;
				IN_DONE = 1'h0;
				clr_blank_done = 1'h0;
				set_blank_done = 1'h0;
				pop_block_wr = 1'h0;
			end
			5'h0e: begin : scan_seq_UL_EMIT_SEG_Output
				data_to_fifo = segment_counter;
				op_to_fifo = 1'h1;
				addr_to_fifo = segment_addr;
				ID_to_fifo = 16'h0000;
				push_to_outs = ~wen_made_sticky & &(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full});
				inc_seg_addr = ~wen_made_sticky & &(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full});
				clr_seg_addr = 1'h0;
				inc_coord_addr = 1'h0;
				clr_coord_addr = 1'h0;
				inc_seg_ctr = 1'h0;
				clr_seg_ctr = 1'h0;
				set_curr_coord = 1'h0;
				clr_curr_coord = 1'h1;
				infifo_pop[0] = ((data_infifo_valid_in & data_infifo_eos_in) & ~(init_blank & ~blank_done_stick_sticky)) & ~data_done_in;
				infifo_pop[1] = 1'h0;
				clr_wen_made = 1'h0;
				set_block_size = 1'h0;
				inc_block_write = 1'h0;
				clr_block_write = 1'h0;
				IN_DONE = 1'h0;
				clr_blank_done = 1'h0;
				set_blank_done = 1'h0;
				pop_block_wr = 1'h0;
			end
			5'h0f: begin : scan_seq_UL_WZ_Output
				data_to_fifo = 16'h0000;
				op_to_fifo = 1'h1;
				addr_to_fifo = segment_addr;
				ID_to_fifo = 16'h0000;
				push_to_outs = 1'h1;
				inc_seg_addr = &(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full});
				clr_seg_addr = 1'h0;
				inc_coord_addr = 1'h0;
				clr_coord_addr = 1'h0;
				inc_seg_ctr = 1'h0;
				clr_seg_ctr = 1'h0;
				set_curr_coord = 1'h0;
				clr_curr_coord = 1'h0;
				infifo_pop[0] = 1'h0;
				infifo_pop[1] = 1'h0;
				clr_wen_made = 1'h0;
				set_block_size = 1'h0;
				inc_block_write = 1'h0;
				clr_block_write = 1'h0;
				IN_DONE = 1'h0;
				clr_blank_done = 1'h0;
				set_blank_done = 1'h0;
				pop_block_wr = 1'h0;
			end
			5'h10: begin : scan_seq_UnLL_Output
				data_to_fifo = data_infifo_data_in;
				op_to_fifo = 1'h1;
				addr_to_fifo = addr_infifo_data_in;
				ID_to_fifo = 16'h0000;
				push_to_outs = (data_infifo_valid_in & addr_infifo_valid_in) & ~(data_infifo_eos_in | addr_infifo_eos_in);
				inc_seg_addr = 1'h0;
				clr_seg_addr = 1'h0;
				inc_coord_addr = 1'h0;
				clr_coord_addr = 1'h0;
				inc_seg_ctr = 1'h0;
				clr_seg_ctr = 1'h0;
				set_curr_coord = 1'h0;
				clr_curr_coord = 1'h0;
				infifo_pop[0] = (data_infifo_valid_in & addr_infifo_valid_in) & ((data_infifo_eos_in & addr_infifo_eos_in) | &(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full}));
				infifo_pop[1] = (data_infifo_valid_in & addr_infifo_valid_in) & ((data_infifo_eos_in & addr_infifo_eos_in) | &(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full}));
				clr_wen_made = 1'h0;
				set_block_size = 1'h0;
				inc_block_write = 1'h0;
				clr_block_write = 1'h0;
				IN_DONE = 1'h0;
				clr_blank_done = 1'h0;
				set_blank_done = 1'h0;
				pop_block_wr = 1'h0;
			end
			default: begin : scan_seq_default_Output
				data_to_fifo = 16'h0000;
				op_to_fifo = 1'h0;
				addr_to_fifo = 16'h0000;
				ID_to_fifo = 16'h0000;
				push_to_outs = 1'h0;
				inc_seg_addr = 1'h0;
				clr_seg_addr = 1'h1;
				inc_coord_addr = 1'h0;
				clr_coord_addr = 1'h1;
				inc_seg_ctr = 1'h0;
				clr_seg_ctr = 1'h1;
				set_curr_coord = 1'h0;
				clr_curr_coord = 1'h1;
				infifo_pop[0] = 1'h0;
				infifo_pop[1] = 1'h0;
				clr_wen_made = 1'h1;
				set_block_size = 1'h0;
				inc_block_write = 1'h0;
				clr_block_write = 1'h1;
				IN_DONE = 1'h0;
				clr_blank_done = 1'h0;
				set_blank_done = 1'h0;
				pop_block_wr = 1'h0;
			end
		endcase
	reg_fifo_depth_0_w_17_afd_2 data_input_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(data_infifo_in_packed),
		.flush(flush),
		.pop(infifo_pop[0]),
		.push(data_in_valid),
		.rst_n(rst_n),
		.data_out(data_infifo_out_packed),
		.empty(data_input_fifo_empty),
		.full(data_input_fifo_full)
	);
	reg_fifo_depth_0_w_17_afd_2 addr_input_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(addr_infifo_in_packed),
		.flush(flush),
		.pop(infifo_pop[1]),
		.push(addr_in_valid),
		.rst_n(rst_n),
		.data_out(addr_infifo_out_packed),
		.empty(addr_input_fifo_empty),
		.full(addr_input_fifo_full)
	);
	reg_fifo_depth_0_w_16_afd_2 block_wr_input_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(block_wr_in[15:0]),
		.flush(flush),
		.pop(pop_block_wr),
		.push(block_wr_in_valid),
		.rst_n(rst_n),
		.data_out(block_wr_input_fifo_data_out),
		.empty(block_wr_input_fifo_empty),
		.full(block_wr_input_fifo_full)
	);
	reg_fifo_depth_2_w_17_afd_2 data_out_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(data_out_fifo_data_in),
		.flush(flush),
		.pop(data_out_ready),
		.push(data_out_fifo_push),
		.rst_n(rst_n),
		.data_out(data_out),
		.empty(data_out_fifo_empty),
		.full(data_out_fifo_full)
	);
	reg_fifo_depth_2_w_17_afd_2 addr_out_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(addr_out_fifo_data_in),
		.flush(flush),
		.pop(addr_out_ready),
		.push(addr_out_fifo_push),
		.rst_n(rst_n),
		.data_out(addr_out),
		.empty(addr_out_fifo_empty),
		.full(addr_out_fifo_full)
	);
	reg_fifo_depth_2_w_17_afd_2 ID_out_fifo(
		.clk(gclk),
		.clk_en(clk_en),
		.data_in(ID_out_fifo_data_in),
		.flush(flush),
		.pop(ID_out_ready),
		.push(ID_out_fifo_push),
		.rst_n(rst_n),
		.data_out(ID_out),
		.empty(ID_out_fifo_empty),
		.full(ID_out_fifo_full)
	);
endmodule
module FanoutHash_F95D10B01D02012 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[0]) | I1;
	assign sel2 = (~E2 | ~S2[1]) | I2;
	assign sel3 = (~E3 | ~S3[0]) | I3;
	assign sel4 = (~E4 | ~S4[0]) | I4;
	assign sel5 = (~E5 | ~S5[0]) | I5;
	assign O = ((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5;
endmodule
module FanoutHash_F8E7A0823DC8CDD (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[2]) | I1;
	assign sel2 = (~E2 | ~S2[2]) | I2;
	assign sel3 = (~E3 | ~S3[11]) | I3;
	assign sel4 = (~E4 | ~S4[11]) | I4;
	assign sel5 = (~E5 | ~S5[11]) | I5;
	assign O = ((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5;
endmodule
module FanoutHash_F689C91787363AB (
	E0,
	E1,
	E10,
	E11,
	E12,
	E13,
	E14,
	E15,
	E16,
	E17,
	E18,
	E19,
	E2,
	E20,
	E3,
	E4,
	E5,
	E6,
	E7,
	E8,
	E9,
	I0,
	I1,
	I10,
	I11,
	I12,
	I13,
	I14,
	I15,
	I16,
	I17,
	I18,
	I19,
	I2,
	I20,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	I9,
	S0,
	S1,
	S10,
	S11,
	S12,
	S13,
	S14,
	S15,
	S16,
	S17,
	S18,
	S19,
	S2,
	S20,
	S3,
	S4,
	S5,
	S6,
	S7,
	S8,
	S9,
	O
);
	input wire E0;
	input wire E1;
	input wire E10;
	input wire E11;
	input wire E12;
	input wire E13;
	input wire E14;
	input wire E15;
	input wire E16;
	input wire E17;
	input wire E18;
	input wire E19;
	input wire E2;
	input wire E20;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire E7;
	input wire E8;
	input wire E9;
	input wire I0;
	input wire I1;
	input wire I10;
	input wire I11;
	input wire I12;
	input wire I13;
	input wire I14;
	input wire I15;
	input wire I16;
	input wire I17;
	input wire I18;
	input wire I19;
	input wire I2;
	input wire I20;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire I7;
	input wire I8;
	input wire I9;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S10;
	input wire [7:0] S11;
	input wire [7:0] S12;
	input wire [7:0] S13;
	input wire [7:0] S14;
	input wire [7:0] S15;
	input wire [7:0] S16;
	input wire [7:0] S17;
	input wire [7:0] S18;
	input wire [7:0] S19;
	input wire [7:0] S2;
	input wire [31:0] S20;
	input wire [7:0] S3;
	input wire [7:0] S4;
	input wire [7:0] S5;
	input wire [7:0] S6;
	input wire [7:0] S7;
	input wire [7:0] S8;
	input wire [7:0] S9;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel10;
	wire sel11;
	wire sel12;
	wire sel13;
	wire sel14;
	wire sel15;
	wire sel16;
	wire sel17;
	wire sel18;
	wire sel19;
	wire sel2;
	wire sel20;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	wire sel7;
	wire sel8;
	wire sel9;
	assign sel0 = (~E0 | ~S0[4]) | I0;
	assign sel1 = (~E1 | ~S1[4]) | I1;
	assign sel2 = (~E2 | ~S2[4]) | I2;
	assign sel3 = (~E3 | ~S3[4]) | I3;
	assign sel4 = (~E4 | ~S4[4]) | I4;
	assign sel5 = (~E5 | ~S5[4]) | I5;
	assign sel6 = (~E6 | ~S6[4]) | I6;
	assign sel7 = (~E7 | ~S7[4]) | I7;
	assign sel8 = (~E8 | ~S8[4]) | I8;
	assign sel9 = (~E9 | ~S9[4]) | I9;
	assign sel10 = (~E10 | ~S10[4]) | I10;
	assign sel11 = (~E11 | ~S11[4]) | I11;
	assign sel12 = (~E12 | ~S12[4]) | I12;
	assign sel13 = (~E13 | ~S13[4]) | I13;
	assign sel14 = (~E14 | ~S14[4]) | I14;
	assign sel15 = (~E15 | ~S15[4]) | I15;
	assign sel16 = (~E16 | ~S16[4]) | I16;
	assign sel17 = (~E17 | ~S17[4]) | I17;
	assign sel18 = (~E18 | ~S18[4]) | I18;
	assign sel19 = (~E19 | ~S19[4]) | I19;
	assign sel20 = (~E20 | ~S20[20]) | I20;
	assign O = (((((((((((((((((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6) & sel7) & sel8) & sel9) & sel10) & sel11) & sel12) & sel13) & sel14) & sel15) & sel16) & sel17) & sel18) & sel19) & sel20;
endmodule
module FanoutHash_E70AF988E4250F5 (
	E0,
	E1,
	E10,
	E11,
	E12,
	E13,
	E14,
	E15,
	E16,
	E17,
	E18,
	E19,
	E2,
	E3,
	E4,
	E5,
	E6,
	E7,
	E8,
	E9,
	I0,
	I1,
	I10,
	I11,
	I12,
	I13,
	I14,
	I15,
	I16,
	I17,
	I18,
	I19,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	I9,
	S0,
	S1,
	S10,
	S11,
	S12,
	S13,
	S14,
	S15,
	S16,
	S17,
	S18,
	S19,
	S2,
	S3,
	S4,
	S5,
	S6,
	S7,
	S8,
	S9,
	O
);
	input wire E0;
	input wire E1;
	input wire E10;
	input wire E11;
	input wire E12;
	input wire E13;
	input wire E14;
	input wire E15;
	input wire E16;
	input wire E17;
	input wire E18;
	input wire E19;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire E7;
	input wire E8;
	input wire E9;
	input wire I0;
	input wire I1;
	input wire I10;
	input wire I11;
	input wire I12;
	input wire I13;
	input wire I14;
	input wire I15;
	input wire I16;
	input wire I17;
	input wire I18;
	input wire I19;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire I7;
	input wire I8;
	input wire I9;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S10;
	input wire [7:0] S11;
	input wire [7:0] S12;
	input wire [7:0] S13;
	input wire [7:0] S14;
	input wire [7:0] S15;
	input wire [7:0] S16;
	input wire [7:0] S17;
	input wire [7:0] S18;
	input wire [7:0] S19;
	input wire [7:0] S2;
	input wire [7:0] S3;
	input wire [7:0] S4;
	input wire [7:0] S5;
	input wire [7:0] S6;
	input wire [7:0] S7;
	input wire [7:0] S8;
	input wire [7:0] S9;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel10;
	wire sel11;
	wire sel12;
	wire sel13;
	wire sel14;
	wire sel15;
	wire sel16;
	wire sel17;
	wire sel18;
	wire sel19;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	wire sel7;
	wire sel8;
	wire sel9;
	assign sel0 = (~E0 | ~S0[3]) | I0;
	assign sel1 = (~E1 | ~S1[3]) | I1;
	assign sel2 = (~E2 | ~S2[3]) | I2;
	assign sel3 = (~E3 | ~S3[3]) | I3;
	assign sel4 = (~E4 | ~S4[3]) | I4;
	assign sel5 = (~E5 | ~S5[3]) | I5;
	assign sel6 = (~E6 | ~S6[3]) | I6;
	assign sel7 = (~E7 | ~S7[3]) | I7;
	assign sel8 = (~E8 | ~S8[3]) | I8;
	assign sel9 = (~E9 | ~S9[3]) | I9;
	assign sel10 = (~E10 | ~S10[3]) | I10;
	assign sel11 = (~E11 | ~S11[3]) | I11;
	assign sel12 = (~E12 | ~S12[3]) | I12;
	assign sel13 = (~E13 | ~S13[3]) | I13;
	assign sel14 = (~E14 | ~S14[3]) | I14;
	assign sel15 = (~E15 | ~S15[3]) | I15;
	assign sel16 = (~E16 | ~S16[3]) | I16;
	assign sel17 = (~E17 | ~S17[3]) | I17;
	assign sel18 = (~E18 | ~S18[3]) | I18;
	assign sel19 = (~E19 | ~S19[3]) | I19;
	assign O = ((((((((((((((((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6) & sel7) & sel8) & sel9) & sel10) & sel11) & sel12) & sel13) & sel14) & sel15) & sel16) & sel17) & sel18) & sel19;
endmodule
module FanoutHash_D70CFBE8EA3CE7F (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[0]) | I1;
	assign sel2 = (~E2 | ~S2[2]) | I2;
	assign sel3 = (~E3 | ~S3[14]) | I3;
	assign sel4 = (~E4 | ~S4[14]) | I4;
	assign sel5 = (~E5 | ~S5[14]) | I5;
	assign O = ((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5;
endmodule
module FanoutHash_CE1AA874B742213 (
	E0,
	E1,
	E10,
	E11,
	E12,
	E13,
	E14,
	E15,
	E16,
	E17,
	E18,
	E19,
	E2,
	E3,
	E4,
	E5,
	E6,
	E7,
	E8,
	E9,
	I0,
	I1,
	I10,
	I11,
	I12,
	I13,
	I14,
	I15,
	I16,
	I17,
	I18,
	I19,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	I9,
	S0,
	S1,
	S10,
	S11,
	S12,
	S13,
	S14,
	S15,
	S16,
	S17,
	S18,
	S19,
	S2,
	S3,
	S4,
	S5,
	S6,
	S7,
	S8,
	S9,
	O
);
	input wire E0;
	input wire E1;
	input wire E10;
	input wire E11;
	input wire E12;
	input wire E13;
	input wire E14;
	input wire E15;
	input wire E16;
	input wire E17;
	input wire E18;
	input wire E19;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire E7;
	input wire E8;
	input wire E9;
	input wire I0;
	input wire I1;
	input wire I10;
	input wire I11;
	input wire I12;
	input wire I13;
	input wire I14;
	input wire I15;
	input wire I16;
	input wire I17;
	input wire I18;
	input wire I19;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire I7;
	input wire I8;
	input wire I9;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S10;
	input wire [7:0] S11;
	input wire [7:0] S12;
	input wire [7:0] S13;
	input wire [7:0] S14;
	input wire [7:0] S15;
	input wire [7:0] S16;
	input wire [7:0] S17;
	input wire [7:0] S18;
	input wire [7:0] S19;
	input wire [7:0] S2;
	input wire [7:0] S3;
	input wire [7:0] S4;
	input wire [7:0] S5;
	input wire [7:0] S6;
	input wire [7:0] S7;
	input wire [7:0] S8;
	input wire [7:0] S9;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel10;
	wire sel11;
	wire sel12;
	wire sel13;
	wire sel14;
	wire sel15;
	wire sel16;
	wire sel17;
	wire sel18;
	wire sel19;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	wire sel7;
	wire sel8;
	wire sel9;
	assign sel0 = (~E0 | ~S0[5]) | I0;
	assign sel1 = (~E1 | ~S1[5]) | I1;
	assign sel2 = (~E2 | ~S2[5]) | I2;
	assign sel3 = (~E3 | ~S3[5]) | I3;
	assign sel4 = (~E4 | ~S4[5]) | I4;
	assign sel5 = (~E5 | ~S5[5]) | I5;
	assign sel6 = (~E6 | ~S6[5]) | I6;
	assign sel7 = (~E7 | ~S7[5]) | I7;
	assign sel8 = (~E8 | ~S8[5]) | I8;
	assign sel9 = (~E9 | ~S9[5]) | I9;
	assign sel10 = (~E10 | ~S10[5]) | I10;
	assign sel11 = (~E11 | ~S11[5]) | I11;
	assign sel12 = (~E12 | ~S12[5]) | I12;
	assign sel13 = (~E13 | ~S13[5]) | I13;
	assign sel14 = (~E14 | ~S14[5]) | I14;
	assign sel15 = (~E15 | ~S15[5]) | I15;
	assign sel16 = (~E16 | ~S16[5]) | I16;
	assign sel17 = (~E17 | ~S17[5]) | I17;
	assign sel18 = (~E18 | ~S18[5]) | I18;
	assign sel19 = (~E19 | ~S19[5]) | I19;
	assign O = ((((((((((((((((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6) & sel7) & sel8) & sel9) & sel10) & sel11) & sel12) & sel13) & sel14) & sel15) & sel16) & sel17) & sel18) & sel19;
endmodule
module FanoutHash_AE7392256DF8B0F (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	E7,
	E8,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	S7,
	S8,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire E7;
	input wire E8;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire I7;
	input wire I8;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	input wire [31:0] S7;
	input wire [31:0] S8;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	wire sel7;
	wire sel8;
	assign sel0 = (~E0 | ~S0[1]) | I0;
	assign sel1 = (~E1 | ~S1[1]) | I1;
	assign sel2 = (~E2 | ~S2[2]) | I2;
	assign sel3 = (~E3 | ~S3[17]) | I3;
	assign sel4 = (~E4 | ~S4[17]) | I4;
	assign sel5 = (~E5 | ~S5[17]) | I5;
	assign sel6 = (~E6 | ~S6[17]) | I6;
	assign sel7 = (~E7 | ~S7[17]) | I7;
	assign sel8 = (~E8 | ~S8[17]) | I8;
	assign O = (((((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6) & sel7) & sel8;
endmodule
module FanoutHash_99D793215CEDDD5 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[2]) | I1;
	assign sel2 = (~E2 | ~S2[1]) | I2;
	assign sel3 = (~E3 | ~S3[1]) | I3;
	assign sel4 = (~E4 | ~S4[1]) | I4;
	assign sel5 = (~E5 | ~S5[1]) | I5;
	assign O = ((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5;
endmodule
module FanoutHash_87642A353688B49 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	E7,
	E8,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	S7,
	S8,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire E7;
	input wire E8;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire I7;
	input wire I8;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	input wire [31:0] S7;
	input wire [31:0] S8;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	wire sel7;
	wire sel8;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[0]) | I1;
	assign sel2 = (~E2 | ~S2[0]) | I2;
	assign sel3 = (~E3 | ~S3[3]) | I3;
	assign sel4 = (~E4 | ~S4[3]) | I4;
	assign sel5 = (~E5 | ~S5[3]) | I5;
	assign sel6 = (~E6 | ~S6[3]) | I6;
	assign sel7 = (~E7 | ~S7[3]) | I7;
	assign sel8 = (~E8 | ~S8[3]) | I8;
	assign O = (((((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6) & sel7) & sel8;
endmodule
module FanoutHash_82899D6851EDC11 (
	E0,
	E1,
	E10,
	E11,
	E12,
	E13,
	E14,
	E15,
	E16,
	E17,
	E18,
	E19,
	E2,
	E3,
	E4,
	E5,
	E6,
	E7,
	E8,
	E9,
	I0,
	I1,
	I10,
	I11,
	I12,
	I13,
	I14,
	I15,
	I16,
	I17,
	I18,
	I19,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	I9,
	S0,
	S1,
	S10,
	S11,
	S12,
	S13,
	S14,
	S15,
	S16,
	S17,
	S18,
	S19,
	S2,
	S3,
	S4,
	S5,
	S6,
	S7,
	S8,
	S9,
	O
);
	input wire E0;
	input wire E1;
	input wire E10;
	input wire E11;
	input wire E12;
	input wire E13;
	input wire E14;
	input wire E15;
	input wire E16;
	input wire E17;
	input wire E18;
	input wire E19;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire E7;
	input wire E8;
	input wire E9;
	input wire I0;
	input wire I1;
	input wire I10;
	input wire I11;
	input wire I12;
	input wire I13;
	input wire I14;
	input wire I15;
	input wire I16;
	input wire I17;
	input wire I18;
	input wire I19;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire I7;
	input wire I8;
	input wire I9;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S10;
	input wire [7:0] S11;
	input wire [7:0] S12;
	input wire [7:0] S13;
	input wire [7:0] S14;
	input wire [7:0] S15;
	input wire [7:0] S16;
	input wire [7:0] S17;
	input wire [7:0] S18;
	input wire [7:0] S19;
	input wire [7:0] S2;
	input wire [7:0] S3;
	input wire [7:0] S4;
	input wire [7:0] S5;
	input wire [7:0] S6;
	input wire [7:0] S7;
	input wire [7:0] S8;
	input wire [7:0] S9;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel10;
	wire sel11;
	wire sel12;
	wire sel13;
	wire sel14;
	wire sel15;
	wire sel16;
	wire sel17;
	wire sel18;
	wire sel19;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	wire sel7;
	wire sel8;
	wire sel9;
	assign sel0 = (~E0 | ~S0[4]) | I0;
	assign sel1 = (~E1 | ~S1[4]) | I1;
	assign sel2 = (~E2 | ~S2[4]) | I2;
	assign sel3 = (~E3 | ~S3[4]) | I3;
	assign sel4 = (~E4 | ~S4[4]) | I4;
	assign sel5 = (~E5 | ~S5[4]) | I5;
	assign sel6 = (~E6 | ~S6[4]) | I6;
	assign sel7 = (~E7 | ~S7[4]) | I7;
	assign sel8 = (~E8 | ~S8[4]) | I8;
	assign sel9 = (~E9 | ~S9[4]) | I9;
	assign sel10 = (~E10 | ~S10[4]) | I10;
	assign sel11 = (~E11 | ~S11[4]) | I11;
	assign sel12 = (~E12 | ~S12[4]) | I12;
	assign sel13 = (~E13 | ~S13[4]) | I13;
	assign sel14 = (~E14 | ~S14[4]) | I14;
	assign sel15 = (~E15 | ~S15[4]) | I15;
	assign sel16 = (~E16 | ~S16[4]) | I16;
	assign sel17 = (~E17 | ~S17[4]) | I17;
	assign sel18 = (~E18 | ~S18[4]) | I18;
	assign sel19 = (~E19 | ~S19[4]) | I19;
	assign O = ((((((((((((((((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6) & sel7) & sel8) & sel9) & sel10) & sel11) & sel12) & sel13) & sel14) & sel15) & sel16) & sel17) & sel18) & sel19;
endmodule
module FanoutHash_7FDF2D3240D4A947 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	assign sel0 = (~E0 | ~S0[2]) | I0;
	assign sel1 = (~E1 | ~S1[2]) | I1;
	assign sel2 = (~E2 | ~S2[2]) | I2;
	assign sel3 = (~E3 | ~S3[15]) | I3;
	assign sel4 = (~E4 | ~S4[15]) | I4;
	assign sel5 = (~E5 | ~S5[15]) | I5;
	assign O = ((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5;
endmodule
module FanoutHash_7F4660D1463D9234 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[0]) | I1;
	assign sel2 = (~E2 | ~S2[2]) | I2;
	assign sel3 = (~E3 | ~S3[10]) | I3;
	assign sel4 = (~E4 | ~S4[10]) | I4;
	assign sel5 = (~E5 | ~S5[10]) | I5;
	assign sel6 = (~E6 | ~S6[10]) | I6;
	assign O = (((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6;
endmodule
module FanoutHash_7ED1C80229B84786 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[2]) | I1;
	assign sel2 = (~E2 | ~S2[1]) | I2;
	assign sel3 = (~E3 | ~S3[7]) | I3;
	assign sel4 = (~E4 | ~S4[7]) | I4;
	assign sel5 = (~E5 | ~S5[7]) | I5;
	assign sel6 = (~E6 | ~S6[7]) | I6;
	assign O = (((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6;
endmodule
module FanoutHash_7E22D83B42537D1D (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	E7,
	E8,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	S7,
	S8,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire E7;
	input wire E8;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire I7;
	input wire I8;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	input wire [31:0] S7;
	input wire [31:0] S8;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	wire sel7;
	wire sel8;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[0]) | I1;
	assign sel2 = (~E2 | ~S2[1]) | I2;
	assign sel3 = (~E3 | ~S3[12]) | I3;
	assign sel4 = (~E4 | ~S4[12]) | I4;
	assign sel5 = (~E5 | ~S5[12]) | I5;
	assign sel6 = (~E6 | ~S6[12]) | I6;
	assign sel7 = (~E7 | ~S7[12]) | I7;
	assign sel8 = (~E8 | ~S8[12]) | I8;
	assign O = (((((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6) & sel7) & sel8;
endmodule
module FanoutHash_752C11B748DD905C (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[2]) | I1;
	assign sel2 = (~E2 | ~S2[2]) | I2;
	assign sel3 = (~E3 | ~S3[11]) | I3;
	assign sel4 = (~E4 | ~S4[11]) | I4;
	assign sel5 = (~E5 | ~S5[11]) | I5;
	assign sel6 = (~E6 | ~S6[11]) | I6;
	assign O = (((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6;
endmodule
module FanoutHash_74A3E41836ECED62 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	E7,
	E8,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	S7,
	S8,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire E7;
	input wire E8;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire I7;
	input wire I8;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	input wire [31:0] S7;
	input wire [31:0] S8;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	wire sel7;
	wire sel8;
	assign sel0 = (~E0 | ~S0[1]) | I0;
	assign sel1 = (~E1 | ~S1[1]) | I1;
	assign sel2 = (~E2 | ~S2[0]) | I2;
	assign sel3 = (~E3 | ~S3[8]) | I3;
	assign sel4 = (~E4 | ~S4[8]) | I4;
	assign sel5 = (~E5 | ~S5[8]) | I5;
	assign sel6 = (~E6 | ~S6[8]) | I6;
	assign sel7 = (~E7 | ~S7[8]) | I7;
	assign sel8 = (~E8 | ~S8[8]) | I8;
	assign O = (((((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6) & sel7) & sel8;
endmodule
module FanoutHash_6EB42FA08A9B7B5B (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	assign sel0 = (~E0 | ~S0[1]) | I0;
	assign sel1 = (~E1 | ~S1[1]) | I1;
	assign sel2 = (~E2 | ~S2[0]) | I2;
	assign sel3 = (~E3 | ~S3[8]) | I3;
	assign sel4 = (~E4 | ~S4[8]) | I4;
	assign sel5 = (~E5 | ~S5[8]) | I5;
	assign O = ((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5;
endmodule
module FanoutHash_6E1094CE0D0F6DFA (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	E7,
	E8,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	S7,
	S8,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire E7;
	input wire E8;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire I7;
	input wire I8;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	input wire [31:0] S7;
	input wire [31:0] S8;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	wire sel7;
	wire sel8;
	assign sel0 = (~E0 | ~S0[2]) | I0;
	assign sel1 = (~E1 | ~S1[2]) | I1;
	assign sel2 = (~E2 | ~S2[2]) | I2;
	assign sel3 = (~E3 | ~S3[19]) | I3;
	assign sel4 = (~E4 | ~S4[19]) | I4;
	assign sel5 = (~E5 | ~S5[19]) | I5;
	assign sel6 = (~E6 | ~S6[19]) | I6;
	assign sel7 = (~E7 | ~S7[19]) | I7;
	assign sel8 = (~E8 | ~S8[19]) | I8;
	assign O = (((((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6) & sel7) & sel8;
endmodule
module FanoutHash_69376833A2418E2 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[0]) | I1;
	assign sel2 = (~E2 | ~S2[1]) | I2;
	assign sel3 = (~E3 | ~S3[12]) | I3;
	assign sel4 = (~E4 | ~S4[12]) | I4;
	assign sel5 = (~E5 | ~S5[12]) | I5;
	assign sel6 = (~E6 | ~S6[12]) | I6;
	assign O = (((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6;
endmodule
module FanoutHash_66A75CC8494A4D6B (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	assign sel0 = (~E0 | ~S0[1]) | I0;
	assign sel1 = (~E1 | ~S1[2]) | I1;
	assign sel2 = (~E2 | ~S2[1]) | I2;
	assign sel3 = (~E3 | ~S3[13]) | I3;
	assign sel4 = (~E4 | ~S4[13]) | I4;
	assign sel5 = (~E5 | ~S5[13]) | I5;
	assign sel6 = (~E6 | ~S6[13]) | I6;
	assign O = (((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6;
endmodule
module FanoutHash_660E59B0DDACF452 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	assign sel0 = (~E0 | ~S0[2]) | I0;
	assign sel1 = (~E1 | ~S1[2]) | I1;
	assign sel2 = (~E2 | ~S2[2]) | I2;
	assign sel3 = (~E3 | ~S3[19]) | I3;
	assign sel4 = (~E4 | ~S4[19]) | I4;
	assign sel5 = (~E5 | ~S5[19]) | I5;
	assign O = ((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5;
endmodule
module FanoutHash_65A468071775C7BB (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[0]) | I1;
	assign sel2 = (~E2 | ~S2[0]) | I2;
	assign sel3 = (~E3 | ~S3[3]) | I3;
	assign sel4 = (~E4 | ~S4[3]) | I4;
	assign sel5 = (~E5 | ~S5[3]) | I5;
	assign sel6 = (~E6 | ~S6[3]) | I6;
	assign O = (((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6;
endmodule
module FanoutHash_653384C8EF52B5E3 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	E7,
	E8,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	S7,
	S8,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire E7;
	input wire E8;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire I7;
	input wire I8;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	input wire [31:0] S7;
	input wire [31:0] S8;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	wire sel7;
	wire sel8;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[2]) | I1;
	assign sel2 = (~E2 | ~S2[1]) | I2;
	assign sel3 = (~E3 | ~S3[7]) | I3;
	assign sel4 = (~E4 | ~S4[7]) | I4;
	assign sel5 = (~E5 | ~S5[7]) | I5;
	assign sel6 = (~E6 | ~S6[7]) | I6;
	assign sel7 = (~E7 | ~S7[7]) | I7;
	assign sel8 = (~E8 | ~S8[7]) | I8;
	assign O = (((((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6) & sel7) & sel8;
endmodule
module FanoutHash_5DE101F5B6936D07 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[0]) | I1;
	assign sel2 = (~E2 | ~S2[1]) | I2;
	assign sel3 = (~E3 | ~S3[12]) | I3;
	assign sel4 = (~E4 | ~S4[12]) | I4;
	assign sel5 = (~E5 | ~S5[12]) | I5;
	assign O = ((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5;
endmodule
module FanoutHash_5D7AEC1255CDC1CC (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	assign sel0 = (~E0 | ~S0[1]) | I0;
	assign sel1 = (~E1 | ~S1[1]) | I1;
	assign sel2 = (~E2 | ~S2[2]) | I2;
	assign sel3 = (~E3 | ~S3[18]) | I3;
	assign sel4 = (~E4 | ~S4[18]) | I4;
	assign sel5 = (~E5 | ~S5[18]) | I5;
	assign sel6 = (~E6 | ~S6[18]) | I6;
	assign O = (((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6;
endmodule
module FanoutHash_5CD8077D054B887B (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	E7,
	E8,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	S7,
	S8,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire E7;
	input wire E8;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire I7;
	input wire I8;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	input wire [31:0] S7;
	input wire [31:0] S8;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	wire sel7;
	wire sel8;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[0]) | I1;
	assign sel2 = (~E2 | ~S2[2]) | I2;
	assign sel3 = (~E3 | ~S3[10]) | I3;
	assign sel4 = (~E4 | ~S4[10]) | I4;
	assign sel5 = (~E5 | ~S5[10]) | I5;
	assign sel6 = (~E6 | ~S6[10]) | I6;
	assign sel7 = (~E7 | ~S7[10]) | I7;
	assign sel8 = (~E8 | ~S8[10]) | I8;
	assign O = (((((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6) & sel7) & sel8;
endmodule
module FanoutHash_59B7E37DAE2221E3 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	E7,
	E8,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	S7,
	S8,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire E7;
	input wire E8;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire I7;
	input wire I8;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	input wire [31:0] S7;
	input wire [31:0] S8;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	wire sel7;
	wire sel8;
	assign sel0 = (~E0 | ~S0[1]) | I0;
	assign sel1 = (~E1 | ~S1[2]) | I1;
	assign sel2 = (~E2 | ~S2[1]) | I2;
	assign sel3 = (~E3 | ~S3[13]) | I3;
	assign sel4 = (~E4 | ~S4[13]) | I4;
	assign sel5 = (~E5 | ~S5[13]) | I5;
	assign sel6 = (~E6 | ~S6[13]) | I6;
	assign sel7 = (~E7 | ~S7[13]) | I7;
	assign sel8 = (~E8 | ~S8[13]) | I8;
	assign O = (((((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6) & sel7) & sel8;
endmodule
module FanoutHash_55B00FA90A0098BB (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	E7,
	E8,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	S7,
	S8,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire E7;
	input wire E8;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire I7;
	input wire I8;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	input wire [31:0] S7;
	input wire [31:0] S8;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	wire sel7;
	wire sel8;
	assign sel0 = (~E0 | ~S0[2]) | I0;
	assign sel1 = (~E1 | ~S1[0]) | I1;
	assign sel2 = (~E2 | ~S2[1]) | I2;
	assign sel3 = (~E3 | ~S3[2]) | I3;
	assign sel4 = (~E4 | ~S4[2]) | I4;
	assign sel5 = (~E5 | ~S5[2]) | I5;
	assign sel6 = (~E6 | ~S6[2]) | I6;
	assign sel7 = (~E7 | ~S7[2]) | I7;
	assign sel8 = (~E8 | ~S8[2]) | I8;
	assign O = (((((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6) & sel7) & sel8;
endmodule
module FanoutHash_55169EB19E10AA09 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	E7,
	E8,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	S7,
	S8,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire E7;
	input wire E8;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire I7;
	input wire I8;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	input wire [31:0] S7;
	input wire [31:0] S8;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	wire sel7;
	wire sel8;
	assign sel0 = (~E0 | ~S0[1]) | I0;
	assign sel1 = (~E1 | ~S1[1]) | I1;
	assign sel2 = (~E2 | ~S2[2]) | I2;
	assign sel3 = (~E3 | ~S3[18]) | I3;
	assign sel4 = (~E4 | ~S4[18]) | I4;
	assign sel5 = (~E5 | ~S5[18]) | I5;
	assign sel6 = (~E6 | ~S6[18]) | I6;
	assign sel7 = (~E7 | ~S7[18]) | I7;
	assign sel8 = (~E8 | ~S8[18]) | I8;
	assign O = (((((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6) & sel7) & sel8;
endmodule
module FanoutHash_4FF010386DB0B737 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	assign sel0 = (~E0 | ~S0[1]) | I0;
	assign sel1 = (~E1 | ~S1[1]) | I1;
	assign sel2 = (~E2 | ~S2[1]) | I2;
	assign sel3 = (~E3 | ~S3[5]) | I3;
	assign sel4 = (~E4 | ~S4[5]) | I4;
	assign sel5 = (~E5 | ~S5[5]) | I5;
	assign O = ((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5;
endmodule
module FanoutHash_4FADDC8F90390680 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[1]) | I1;
	assign sel2 = (~E2 | ~S2[0]) | I2;
	assign sel3 = (~E3 | ~S3[4]) | I3;
	assign sel4 = (~E4 | ~S4[4]) | I4;
	assign sel5 = (~E5 | ~S5[4]) | I5;
	assign sel6 = (~E6 | ~S6[4]) | I6;
	assign O = (((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6;
endmodule
module FanoutHash_4F83851A40824F89 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	assign sel0 = (~E0 | ~S0[1]) | I0;
	assign sel1 = (~E1 | ~S1[2]) | I1;
	assign sel2 = (~E2 | ~S2[0]) | I2;
	assign sel3 = (~E3 | ~S3[6]) | I3;
	assign sel4 = (~E4 | ~S4[6]) | I4;
	assign sel5 = (~E5 | ~S5[6]) | I5;
	assign sel6 = (~E6 | ~S6[6]) | I6;
	assign O = (((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6;
endmodule
module FanoutHash_4A74B16B611BA7E4 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	E7,
	E8,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	S7,
	S8,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire E7;
	input wire E8;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire I7;
	input wire I8;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	input wire [31:0] S7;
	input wire [31:0] S8;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	wire sel7;
	wire sel8;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[2]) | I1;
	assign sel2 = (~E2 | ~S2[2]) | I2;
	assign sel3 = (~E3 | ~S3[11]) | I3;
	assign sel4 = (~E4 | ~S4[11]) | I4;
	assign sel5 = (~E5 | ~S5[11]) | I5;
	assign sel6 = (~E6 | ~S6[11]) | I6;
	assign sel7 = (~E7 | ~S7[11]) | I7;
	assign sel8 = (~E8 | ~S8[11]) | I8;
	assign O = (((((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6) & sel7) & sel8;
endmodule
module FanoutHash_47712AAC902ADA2 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[0]) | I1;
	assign sel2 = (~E2 | ~S2[1]) | I2;
	assign sel3 = (~E3 | ~S3[0]) | I3;
	assign sel4 = (~E4 | ~S4[0]) | I4;
	assign sel5 = (~E5 | ~S5[0]) | I5;
	assign sel6 = (~E6 | ~S6[0]) | I6;
	assign O = (((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6;
endmodule
module FanoutHash_4678C6877F96240E (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	assign sel0 = (~E0 | ~S0[2]) | I0;
	assign sel1 = (~E1 | ~S1[0]) | I1;
	assign sel2 = (~E2 | ~S2[1]) | I2;
	assign sel3 = (~E3 | ~S3[2]) | I3;
	assign sel4 = (~E4 | ~S4[2]) | I4;
	assign sel5 = (~E5 | ~S5[2]) | I5;
	assign O = ((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5;
endmodule
module FanoutHash_466EB88CFD0CAD7B (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	assign sel0 = (~E0 | ~S0[1]) | I0;
	assign sel1 = (~E1 | ~S1[1]) | I1;
	assign sel2 = (~E2 | ~S2[1]) | I2;
	assign sel3 = (~E3 | ~S3[5]) | I3;
	assign sel4 = (~E4 | ~S4[5]) | I4;
	assign sel5 = (~E5 | ~S5[5]) | I5;
	assign sel6 = (~E6 | ~S6[5]) | I6;
	assign O = (((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6;
endmodule
module FanoutHash_43D5C80ABD816837 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[0]) | I1;
	assign sel2 = (~E2 | ~S2[2]) | I2;
	assign sel3 = (~E3 | ~S3[14]) | I3;
	assign sel4 = (~E4 | ~S4[14]) | I4;
	assign sel5 = (~E5 | ~S5[14]) | I5;
	assign sel6 = (~E6 | ~S6[14]) | I6;
	assign O = (((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6;
endmodule
module FanoutHash_41D739158D58E184 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	E7,
	E8,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	S7,
	S8,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire E7;
	input wire E8;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire I7;
	input wire I8;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	input wire [31:0] S7;
	input wire [31:0] S8;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	wire sel7;
	wire sel8;
	assign sel0 = (~E0 | ~S0[2]) | I0;
	assign sel1 = (~E1 | ~S1[2]) | I1;
	assign sel2 = (~E2 | ~S2[2]) | I2;
	assign sel3 = (~E3 | ~S3[15]) | I3;
	assign sel4 = (~E4 | ~S4[15]) | I4;
	assign sel5 = (~E5 | ~S5[15]) | I5;
	assign sel6 = (~E6 | ~S6[15]) | I6;
	assign sel7 = (~E7 | ~S7[15]) | I7;
	assign sel8 = (~E8 | ~S8[15]) | I8;
	assign O = (((((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6) & sel7) & sel8;
endmodule
module FanoutHash_3E05574A9CE9CA8A (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	E7,
	E8,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	S7,
	S8,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire E7;
	input wire E8;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire I7;
	input wire I8;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	input wire [31:0] S7;
	input wire [31:0] S8;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	wire sel7;
	wire sel8;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[2]) | I1;
	assign sel2 = (~E2 | ~S2[1]) | I2;
	assign sel3 = (~E3 | ~S3[1]) | I3;
	assign sel4 = (~E4 | ~S4[1]) | I4;
	assign sel5 = (~E5 | ~S5[1]) | I5;
	assign sel6 = (~E6 | ~S6[1]) | I6;
	assign sel7 = (~E7 | ~S7[1]) | I7;
	assign sel8 = (~E8 | ~S8[1]) | I8;
	assign O = (((((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6) & sel7) & sel8;
endmodule
module FanoutHash_3B67229CB02928BA (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	assign sel0 = (~E0 | ~S0[1]) | I0;
	assign sel1 = (~E1 | ~S1[1]) | I1;
	assign sel2 = (~E2 | ~S2[0]) | I2;
	assign sel3 = (~E3 | ~S3[8]) | I3;
	assign sel4 = (~E4 | ~S4[8]) | I4;
	assign sel5 = (~E5 | ~S5[8]) | I5;
	assign sel6 = (~E6 | ~S6[8]) | I6;
	assign O = (((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6;
endmodule
module FanoutHash_3A6A5822E84DCC71 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	E7,
	E8,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	S7,
	S8,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire E7;
	input wire E8;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire I7;
	input wire I8;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	input wire [31:0] S7;
	input wire [31:0] S8;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	wire sel7;
	wire sel8;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[0]) | I1;
	assign sel2 = (~E2 | ~S2[1]) | I2;
	assign sel3 = (~E3 | ~S3[0]) | I3;
	assign sel4 = (~E4 | ~S4[0]) | I4;
	assign sel5 = (~E5 | ~S5[0]) | I5;
	assign sel6 = (~E6 | ~S6[0]) | I6;
	assign sel7 = (~E7 | ~S7[0]) | I7;
	assign sel8 = (~E8 | ~S8[0]) | I8;
	assign O = (((((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6) & sel7) & sel8;
endmodule
module FanoutHash_3A0064632A577CF5 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[0]) | I1;
	assign sel2 = (~E2 | ~S2[0]) | I2;
	assign sel3 = (~E3 | ~S3[3]) | I3;
	assign sel4 = (~E4 | ~S4[3]) | I4;
	assign sel5 = (~E5 | ~S5[3]) | I5;
	assign O = ((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5;
endmodule
module FanoutHash_37E9FE88073C5BAC (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	E7,
	E8,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	S7,
	S8,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire E7;
	input wire E8;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire I7;
	input wire I8;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	input wire [31:0] S7;
	input wire [31:0] S8;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	wire sel7;
	wire sel8;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[1]) | I1;
	assign sel2 = (~E2 | ~S2[0]) | I2;
	assign sel3 = (~E3 | ~S3[4]) | I3;
	assign sel4 = (~E4 | ~S4[4]) | I4;
	assign sel5 = (~E5 | ~S5[4]) | I5;
	assign sel6 = (~E6 | ~S6[4]) | I6;
	assign sel7 = (~E7 | ~S7[4]) | I7;
	assign sel8 = (~E8 | ~S8[4]) | I8;
	assign O = (((((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6) & sel7) & sel8;
endmodule
module FanoutHash_37B926A0CDF82FCC (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[2]) | I1;
	assign sel2 = (~E2 | ~S2[2]) | I2;
	assign sel3 = (~E3 | ~S3[16]) | I3;
	assign sel4 = (~E4 | ~S4[16]) | I4;
	assign sel5 = (~E5 | ~S5[16]) | I5;
	assign O = ((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5;
endmodule
module FanoutHash_330DF95D65589621 (
	E0,
	E1,
	E10,
	E11,
	E12,
	E13,
	E14,
	E15,
	E16,
	E17,
	E18,
	E19,
	E2,
	E20,
	E21,
	E3,
	E4,
	E5,
	E6,
	E7,
	E8,
	E9,
	I0,
	I1,
	I10,
	I11,
	I12,
	I13,
	I14,
	I15,
	I16,
	I17,
	I18,
	I19,
	I2,
	I20,
	I21,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	I9,
	S0,
	S1,
	S10,
	S11,
	S12,
	S13,
	S14,
	S15,
	S16,
	S17,
	S18,
	S19,
	S2,
	S20,
	S21,
	S3,
	S4,
	S5,
	S6,
	S7,
	S8,
	S9,
	O
);
	input wire E0;
	input wire E1;
	input wire E10;
	input wire E11;
	input wire E12;
	input wire E13;
	input wire E14;
	input wire E15;
	input wire E16;
	input wire E17;
	input wire E18;
	input wire E19;
	input wire E2;
	input wire E20;
	input wire E21;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire E7;
	input wire E8;
	input wire E9;
	input wire I0;
	input wire I1;
	input wire I10;
	input wire I11;
	input wire I12;
	input wire I13;
	input wire I14;
	input wire I15;
	input wire I16;
	input wire I17;
	input wire I18;
	input wire I19;
	input wire I2;
	input wire I20;
	input wire I21;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire I7;
	input wire I8;
	input wire I9;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S10;
	input wire [7:0] S11;
	input wire [7:0] S12;
	input wire [7:0] S13;
	input wire [7:0] S14;
	input wire [7:0] S15;
	input wire [7:0] S16;
	input wire [7:0] S17;
	input wire [7:0] S18;
	input wire [7:0] S19;
	input wire [7:0] S2;
	input wire [31:0] S20;
	input wire [31:0] S21;
	input wire [7:0] S3;
	input wire [7:0] S4;
	input wire [7:0] S5;
	input wire [7:0] S6;
	input wire [7:0] S7;
	input wire [7:0] S8;
	input wire [7:0] S9;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel10;
	wire sel11;
	wire sel12;
	wire sel13;
	wire sel14;
	wire sel15;
	wire sel16;
	wire sel17;
	wire sel18;
	wire sel19;
	wire sel2;
	wire sel20;
	wire sel21;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	wire sel7;
	wire sel8;
	wire sel9;
	assign sel0 = (~E0 | ~S0[3]) | I0;
	assign sel1 = (~E1 | ~S1[3]) | I1;
	assign sel2 = (~E2 | ~S2[3]) | I2;
	assign sel3 = (~E3 | ~S3[3]) | I3;
	assign sel4 = (~E4 | ~S4[3]) | I4;
	assign sel5 = (~E5 | ~S5[3]) | I5;
	assign sel6 = (~E6 | ~S6[3]) | I6;
	assign sel7 = (~E7 | ~S7[3]) | I7;
	assign sel8 = (~E8 | ~S8[3]) | I8;
	assign sel9 = (~E9 | ~S9[3]) | I9;
	assign sel10 = (~E10 | ~S10[3]) | I10;
	assign sel11 = (~E11 | ~S11[3]) | I11;
	assign sel12 = (~E12 | ~S12[3]) | I12;
	assign sel13 = (~E13 | ~S13[3]) | I13;
	assign sel14 = (~E14 | ~S14[3]) | I14;
	assign sel15 = (~E15 | ~S15[3]) | I15;
	assign sel16 = (~E16 | ~S16[3]) | I16;
	assign sel17 = (~E17 | ~S17[3]) | I17;
	assign sel18 = (~E18 | ~S18[3]) | I18;
	assign sel19 = (~E19 | ~S19[3]) | I19;
	assign sel20 = (~E20 | ~S20[20]) | I20;
	assign sel21 = (~E21 | ~S21[20]) | I21;
	assign O = ((((((((((((((((((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6) & sel7) & sel8) & sel9) & sel10) & sel11) & sel12) & sel13) & sel14) & sel15) & sel16) & sel17) & sel18) & sel19) & sel20) & sel21;
endmodule
module FanoutHash_31AE65CCDD94603 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	assign sel0 = (~E0 | ~S0[2]) | I0;
	assign sel1 = (~E1 | ~S1[2]) | I1;
	assign sel2 = (~E2 | ~S2[2]) | I2;
	assign sel3 = (~E3 | ~S3[15]) | I3;
	assign sel4 = (~E4 | ~S4[15]) | I4;
	assign sel5 = (~E5 | ~S5[15]) | I5;
	assign sel6 = (~E6 | ~S6[15]) | I6;
	assign O = (((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6;
endmodule
module FanoutHash_31555E0CDC460B97 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[1]) | I1;
	assign sel2 = (~E2 | ~S2[0]) | I2;
	assign sel3 = (~E3 | ~S3[4]) | I3;
	assign sel4 = (~E4 | ~S4[4]) | I4;
	assign sel5 = (~E5 | ~S5[4]) | I5;
	assign O = ((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5;
endmodule
module FanoutHash_308BAC760F688049 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	assign sel0 = (~E0 | ~S0[2]) | I0;
	assign sel1 = (~E1 | ~S1[1]) | I1;
	assign sel2 = (~E2 | ~S2[1]) | I2;
	assign sel3 = (~E3 | ~S3[9]) | I3;
	assign sel4 = (~E4 | ~S4[9]) | I4;
	assign sel5 = (~E5 | ~S5[9]) | I5;
	assign O = ((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5;
endmodule
module FanoutHash_302974B49BE3F0C4 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	assign sel0 = (~E0 | ~S0[2]) | I0;
	assign sel1 = (~E1 | ~S1[0]) | I1;
	assign sel2 = (~E2 | ~S2[1]) | I2;
	assign sel3 = (~E3 | ~S3[2]) | I3;
	assign sel4 = (~E4 | ~S4[2]) | I4;
	assign sel5 = (~E5 | ~S5[2]) | I5;
	assign sel6 = (~E6 | ~S6[2]) | I6;
	assign O = (((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6;
endmodule
module FanoutHash_2F92967E9F56D548 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	E7,
	E8,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	S7,
	S8,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire E7;
	input wire E8;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire I7;
	input wire I8;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	input wire [31:0] S7;
	input wire [31:0] S8;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	wire sel7;
	wire sel8;
	assign sel0 = (~E0 | ~S0[1]) | I0;
	assign sel1 = (~E1 | ~S1[1]) | I1;
	assign sel2 = (~E2 | ~S2[1]) | I2;
	assign sel3 = (~E3 | ~S3[5]) | I3;
	assign sel4 = (~E4 | ~S4[5]) | I4;
	assign sel5 = (~E5 | ~S5[5]) | I5;
	assign sel6 = (~E6 | ~S6[5]) | I6;
	assign sel7 = (~E7 | ~S7[5]) | I7;
	assign sel8 = (~E8 | ~S8[5]) | I8;
	assign O = (((((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6) & sel7) & sel8;
endmodule
module FanoutHash_2CE3041FDDDDEC1A (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	E7,
	E8,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	S7,
	S8,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire E7;
	input wire E8;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire I7;
	input wire I8;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	input wire [31:0] S7;
	input wire [31:0] S8;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	wire sel7;
	wire sel8;
	assign sel0 = (~E0 | ~S0[2]) | I0;
	assign sel1 = (~E1 | ~S1[1]) | I1;
	assign sel2 = (~E2 | ~S2[1]) | I2;
	assign sel3 = (~E3 | ~S3[9]) | I3;
	assign sel4 = (~E4 | ~S4[9]) | I4;
	assign sel5 = (~E5 | ~S5[9]) | I5;
	assign sel6 = (~E6 | ~S6[9]) | I6;
	assign sel7 = (~E7 | ~S7[9]) | I7;
	assign sel8 = (~E8 | ~S8[9]) | I8;
	assign O = (((((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6) & sel7) & sel8;
endmodule
module FanoutHash_28125A548B305607 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	assign sel0 = (~E0 | ~S0[2]) | I0;
	assign sel1 = (~E1 | ~S1[1]) | I1;
	assign sel2 = (~E2 | ~S2[1]) | I2;
	assign sel3 = (~E3 | ~S3[9]) | I3;
	assign sel4 = (~E4 | ~S4[9]) | I4;
	assign sel5 = (~E5 | ~S5[9]) | I5;
	assign sel6 = (~E6 | ~S6[9]) | I6;
	assign O = (((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6;
endmodule
module FanoutHash_2785CE916183C5C (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[2]) | I1;
	assign sel2 = (~E2 | ~S2[1]) | I2;
	assign sel3 = (~E3 | ~S3[1]) | I3;
	assign sel4 = (~E4 | ~S4[1]) | I4;
	assign sel5 = (~E5 | ~S5[1]) | I5;
	assign sel6 = (~E6 | ~S6[1]) | I6;
	assign O = (((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6;
endmodule
module FanoutHash_278348DB702230E6 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[0]) | I1;
	assign sel2 = (~E2 | ~S2[2]) | I2;
	assign sel3 = (~E3 | ~S3[10]) | I3;
	assign sel4 = (~E4 | ~S4[10]) | I4;
	assign sel5 = (~E5 | ~S5[10]) | I5;
	assign O = ((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5;
endmodule
module FanoutHash_276F8381CE025648 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	E7,
	E8,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	S7,
	S8,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire E7;
	input wire E8;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire I7;
	input wire I8;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	input wire [31:0] S7;
	input wire [31:0] S8;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	wire sel7;
	wire sel8;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[0]) | I1;
	assign sel2 = (~E2 | ~S2[2]) | I2;
	assign sel3 = (~E3 | ~S3[14]) | I3;
	assign sel4 = (~E4 | ~S4[14]) | I4;
	assign sel5 = (~E5 | ~S5[14]) | I5;
	assign sel6 = (~E6 | ~S6[14]) | I6;
	assign sel7 = (~E7 | ~S7[14]) | I7;
	assign sel8 = (~E8 | ~S8[14]) | I8;
	assign O = (((((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6) & sel7) & sel8;
endmodule
module FanoutHash_26B6474864379B6A (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	assign sel0 = (~E0 | ~S0[1]) | I0;
	assign sel1 = (~E1 | ~S1[1]) | I1;
	assign sel2 = (~E2 | ~S2[2]) | I2;
	assign sel3 = (~E3 | ~S3[17]) | I3;
	assign sel4 = (~E4 | ~S4[17]) | I4;
	assign sel5 = (~E5 | ~S5[17]) | I5;
	assign sel6 = (~E6 | ~S6[17]) | I6;
	assign O = (((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6;
endmodule
module FanoutHash_245560850976C879 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	E7,
	E8,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	S7,
	S8,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire E7;
	input wire E8;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire I7;
	input wire I8;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	input wire [31:0] S7;
	input wire [31:0] S8;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	wire sel7;
	wire sel8;
	assign sel0 = (~E0 | ~S0[1]) | I0;
	assign sel1 = (~E1 | ~S1[2]) | I1;
	assign sel2 = (~E2 | ~S2[0]) | I2;
	assign sel3 = (~E3 | ~S3[6]) | I3;
	assign sel4 = (~E4 | ~S4[6]) | I4;
	assign sel5 = (~E5 | ~S5[6]) | I5;
	assign sel6 = (~E6 | ~S6[6]) | I6;
	assign sel7 = (~E7 | ~S7[6]) | I7;
	assign sel8 = (~E8 | ~S8[6]) | I8;
	assign O = (((((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6) & sel7) & sel8;
endmodule
module FanoutHash_244497FCED8BEB80 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	E7,
	E8,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	S7,
	S8,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire E7;
	input wire E8;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire I7;
	input wire I8;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	input wire [31:0] S7;
	input wire [31:0] S8;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	wire sel7;
	wire sel8;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[2]) | I1;
	assign sel2 = (~E2 | ~S2[2]) | I2;
	assign sel3 = (~E3 | ~S3[16]) | I3;
	assign sel4 = (~E4 | ~S4[16]) | I4;
	assign sel5 = (~E5 | ~S5[16]) | I5;
	assign sel6 = (~E6 | ~S6[16]) | I6;
	assign sel7 = (~E7 | ~S7[16]) | I7;
	assign sel8 = (~E8 | ~S8[16]) | I8;
	assign O = (((((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6) & sel7) & sel8;
endmodule
module FanoutHash_1EBD0270673B29D7 (
	E0,
	E1,
	E10,
	E11,
	E12,
	E13,
	E14,
	E15,
	E16,
	E17,
	E18,
	E19,
	E2,
	E3,
	E4,
	E5,
	E6,
	E7,
	E8,
	E9,
	I0,
	I1,
	I10,
	I11,
	I12,
	I13,
	I14,
	I15,
	I16,
	I17,
	I18,
	I19,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	I9,
	S0,
	S1,
	S10,
	S11,
	S12,
	S13,
	S14,
	S15,
	S16,
	S17,
	S18,
	S19,
	S2,
	S3,
	S4,
	S5,
	S6,
	S7,
	S8,
	S9,
	O
);
	input wire E0;
	input wire E1;
	input wire E10;
	input wire E11;
	input wire E12;
	input wire E13;
	input wire E14;
	input wire E15;
	input wire E16;
	input wire E17;
	input wire E18;
	input wire E19;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire E7;
	input wire E8;
	input wire E9;
	input wire I0;
	input wire I1;
	input wire I10;
	input wire I11;
	input wire I12;
	input wire I13;
	input wire I14;
	input wire I15;
	input wire I16;
	input wire I17;
	input wire I18;
	input wire I19;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire I7;
	input wire I8;
	input wire I9;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S10;
	input wire [7:0] S11;
	input wire [7:0] S12;
	input wire [7:0] S13;
	input wire [7:0] S14;
	input wire [7:0] S15;
	input wire [7:0] S16;
	input wire [7:0] S17;
	input wire [7:0] S18;
	input wire [7:0] S19;
	input wire [7:0] S2;
	input wire [7:0] S3;
	input wire [7:0] S4;
	input wire [7:0] S5;
	input wire [7:0] S6;
	input wire [7:0] S7;
	input wire [7:0] S8;
	input wire [7:0] S9;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel10;
	wire sel11;
	wire sel12;
	wire sel13;
	wire sel14;
	wire sel15;
	wire sel16;
	wire sel17;
	wire sel18;
	wire sel19;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	wire sel7;
	wire sel8;
	wire sel9;
	assign sel0 = (~E0 | ~S0[6]) | I0;
	assign sel1 = (~E1 | ~S1[6]) | I1;
	assign sel2 = (~E2 | ~S2[6]) | I2;
	assign sel3 = (~E3 | ~S3[6]) | I3;
	assign sel4 = (~E4 | ~S4[6]) | I4;
	assign sel5 = (~E5 | ~S5[6]) | I5;
	assign sel6 = (~E6 | ~S6[6]) | I6;
	assign sel7 = (~E7 | ~S7[6]) | I7;
	assign sel8 = (~E8 | ~S8[6]) | I8;
	assign sel9 = (~E9 | ~S9[6]) | I9;
	assign sel10 = (~E10 | ~S10[6]) | I10;
	assign sel11 = (~E11 | ~S11[6]) | I11;
	assign sel12 = (~E12 | ~S12[6]) | I12;
	assign sel13 = (~E13 | ~S13[6]) | I13;
	assign sel14 = (~E14 | ~S14[6]) | I14;
	assign sel15 = (~E15 | ~S15[6]) | I15;
	assign sel16 = (~E16 | ~S16[6]) | I16;
	assign sel17 = (~E17 | ~S17[6]) | I17;
	assign sel18 = (~E18 | ~S18[6]) | I18;
	assign sel19 = (~E19 | ~S19[6]) | I19;
	assign O = ((((((((((((((((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6) & sel7) & sel8) & sel9) & sel10) & sel11) & sel12) & sel13) & sel14) & sel15) & sel16) & sel17) & sel18) & sel19;
endmodule
module FanoutHash_1B10C32F008C11AC (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	assign sel0 = (~E0 | ~S0[1]) | I0;
	assign sel1 = (~E1 | ~S1[1]) | I1;
	assign sel2 = (~E2 | ~S2[2]) | I2;
	assign sel3 = (~E3 | ~S3[17]) | I3;
	assign sel4 = (~E4 | ~S4[17]) | I4;
	assign sel5 = (~E5 | ~S5[17]) | I5;
	assign O = ((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5;
endmodule
module FanoutHash_1A568579D8E9714B (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[2]) | I1;
	assign sel2 = (~E2 | ~S2[1]) | I2;
	assign sel3 = (~E3 | ~S3[7]) | I3;
	assign sel4 = (~E4 | ~S4[7]) | I4;
	assign sel5 = (~E5 | ~S5[7]) | I5;
	assign O = ((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5;
endmodule
module FanoutHash_184DFC10DAF19BE9 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	assign sel0 = (~E0 | ~S0[0]) | I0;
	assign sel1 = (~E1 | ~S1[2]) | I1;
	assign sel2 = (~E2 | ~S2[2]) | I2;
	assign sel3 = (~E3 | ~S3[16]) | I3;
	assign sel4 = (~E4 | ~S4[16]) | I4;
	assign sel5 = (~E5 | ~S5[16]) | I5;
	assign sel6 = (~E6 | ~S6[16]) | I6;
	assign O = (((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6;
endmodule
module FanoutHash_1816466D6957000 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	E6,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	S6,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire E6;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire I6;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	input wire [31:0] S6;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	wire sel6;
	assign sel0 = (~E0 | ~S0[2]) | I0;
	assign sel1 = (~E1 | ~S1[2]) | I1;
	assign sel2 = (~E2 | ~S2[2]) | I2;
	assign sel3 = (~E3 | ~S3[19]) | I3;
	assign sel4 = (~E4 | ~S4[19]) | I4;
	assign sel5 = (~E5 | ~S5[19]) | I5;
	assign sel6 = (~E6 | ~S6[19]) | I6;
	assign O = (((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5) & sel6;
endmodule
module FanoutHash_14EBE1E8E49CA541 (
	E0,
	E1,
	E2,
	I0,
	I1,
	I2,
	S0,
	S1,
	S2,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire [31:0] S0;
	input wire [31:0] S1;
	input wire [31:0] S2;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	assign sel0 = (~E0 | ~S0[20]) | I0;
	assign sel1 = (~E1 | ~S1[20]) | I1;
	assign sel2 = (~E2 | ~S2[20]) | I2;
	assign O = (sel0 & sel1) & sel2;
endmodule
module FanoutHash_13B77C2790BDE4E2 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	assign sel0 = (~E0 | ~S0[1]) | I0;
	assign sel1 = (~E1 | ~S1[2]) | I1;
	assign sel2 = (~E2 | ~S2[1]) | I2;
	assign sel3 = (~E3 | ~S3[13]) | I3;
	assign sel4 = (~E4 | ~S4[13]) | I4;
	assign sel5 = (~E5 | ~S5[13]) | I5;
	assign O = ((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5;
endmodule
module FanoutHash_11B554A18790BBBC (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	assign sel0 = (~E0 | ~S0[1]) | I0;
	assign sel1 = (~E1 | ~S1[1]) | I1;
	assign sel2 = (~E2 | ~S2[2]) | I2;
	assign sel3 = (~E3 | ~S3[18]) | I3;
	assign sel4 = (~E4 | ~S4[18]) | I4;
	assign sel5 = (~E5 | ~S5[18]) | I5;
	assign O = ((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5;
endmodule
module FanoutHash_1130FCC7DFE98006 (
	E0,
	E1,
	E2,
	E3,
	E4,
	E5,
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	S0,
	S1,
	S2,
	S3,
	S4,
	S5,
	O
);
	input wire E0;
	input wire E1;
	input wire E2;
	input wire E3;
	input wire E4;
	input wire E5;
	input wire I0;
	input wire I1;
	input wire I2;
	input wire I3;
	input wire I4;
	input wire I5;
	input wire [7:0] S0;
	input wire [7:0] S1;
	input wire [7:0] S2;
	input wire [31:0] S3;
	input wire [31:0] S4;
	input wire [31:0] S5;
	output wire O;
	wire sel0;
	wire sel1;
	wire sel2;
	wire sel3;
	wire sel4;
	wire sel5;
	assign sel0 = (~E0 | ~S0[1]) | I0;
	assign sel1 = (~E1 | ~S1[2]) | I1;
	assign sel2 = (~E2 | ~S2[0]) | I2;
	assign sel3 = (~E3 | ~S3[6]) | I3;
	assign sel4 = (~E4 | ~S4[6]) | I4;
	assign sel5 = (~E5 | ~S5[6]) | I5;
	assign O = ((((sel0 & sel1) & sel2) & sel3) & sel4) & sel5;
endmodule
module ExclusiveNodeFanout_H2 (
	I,
	S,
	O
);
	input wire [1:0] I;
	input wire [1:0] S;
	output wire O;
	assign O = (I[0] & S[0]) | (I[1] & S[1]);
endmodule
module Decode98 (
	I,
	O
);
	input [7:0] I;
	output wire O;
	wire [7:0] const_9_8_out;
	wire coreir_eq_8_inst0_out;
	coreir_const #(
		.value(8'h09),
		.width(8)
	) const_9_8(.out(const_9_8_out));
	coreir_eq #(.width(8)) coreir_eq_8_inst0(
		.in0(I),
		.in1(const_9_8_out),
		.out(coreir_eq_8_inst0_out)
	);
	assign O = coreir_eq_8_inst0_out;
endmodule
module Decode88 (
	I,
	O
);
	input [7:0] I;
	output wire O;
	wire [7:0] const_8_8_out;
	wire coreir_eq_8_inst0_out;
	coreir_const #(
		.value(8'h08),
		.width(8)
	) const_8_8(.out(const_8_8_out));
	coreir_eq #(.width(8)) coreir_eq_8_inst0(
		.in0(I),
		.in1(const_8_8_out),
		.out(coreir_eq_8_inst0_out)
	);
	assign O = coreir_eq_8_inst0_out;
endmodule
module Decode78 (
	I,
	O
);
	input [7:0] I;
	output wire O;
	wire [7:0] const_7_8_out;
	wire coreir_eq_8_inst0_out;
	coreir_const #(
		.value(8'h07),
		.width(8)
	) const_7_8(.out(const_7_8_out));
	coreir_eq #(.width(8)) coreir_eq_8_inst0(
		.in0(I),
		.in1(const_7_8_out),
		.out(coreir_eq_8_inst0_out)
	);
	assign O = coreir_eq_8_inst0_out;
endmodule
module Decode68 (
	I,
	O
);
	input [7:0] I;
	output wire O;
	wire [7:0] const_6_8_out;
	wire coreir_eq_8_inst0_out;
	coreir_const #(
		.value(8'h06),
		.width(8)
	) const_6_8(.out(const_6_8_out));
	coreir_eq #(.width(8)) coreir_eq_8_inst0(
		.in0(I),
		.in1(const_6_8_out),
		.out(coreir_eq_8_inst0_out)
	);
	assign O = coreir_eq_8_inst0_out;
endmodule
module Decode58 (
	I,
	O
);
	input [7:0] I;
	output wire O;
	wire [7:0] const_5_8_out;
	wire coreir_eq_8_inst0_out;
	coreir_const #(
		.value(8'h05),
		.width(8)
	) const_5_8(.out(const_5_8_out));
	coreir_eq #(.width(8)) coreir_eq_8_inst0(
		.in0(I),
		.in1(const_5_8_out),
		.out(coreir_eq_8_inst0_out)
	);
	assign O = coreir_eq_8_inst0_out;
endmodule
module Decode48 (
	I,
	O
);
	input [7:0] I;
	output wire O;
	wire [7:0] const_4_8_out;
	wire coreir_eq_8_inst0_out;
	coreir_const #(
		.value(8'h04),
		.width(8)
	) const_4_8(.out(const_4_8_out));
	coreir_eq #(.width(8)) coreir_eq_8_inst0(
		.in0(I),
		.in1(const_4_8_out),
		.out(coreir_eq_8_inst0_out)
	);
	assign O = coreir_eq_8_inst0_out;
endmodule
module Decode38 (
	I,
	O
);
	input [7:0] I;
	output wire O;
	wire [7:0] const_3_8_out;
	wire coreir_eq_8_inst0_out;
	coreir_const #(
		.value(8'h03),
		.width(8)
	) const_3_8(.out(const_3_8_out));
	coreir_eq #(.width(8)) coreir_eq_8_inst0(
		.in0(I),
		.in1(const_3_8_out),
		.out(coreir_eq_8_inst0_out)
	);
	assign O = coreir_eq_8_inst0_out;
endmodule
module Decode28 (
	I,
	O
);
	input [7:0] I;
	output wire O;
	wire [7:0] const_2_8_out;
	wire coreir_eq_8_inst0_out;
	coreir_const #(
		.value(8'h02),
		.width(8)
	) const_2_8(.out(const_2_8_out));
	coreir_eq #(.width(8)) coreir_eq_8_inst0(
		.in0(I),
		.in1(const_2_8_out),
		.out(coreir_eq_8_inst0_out)
	);
	assign O = coreir_eq_8_inst0_out;
endmodule
module Decode18 (
	I,
	O
);
	input [7:0] I;
	output wire O;
	wire [7:0] const_1_8_out;
	wire coreir_eq_8_inst0_out;
	coreir_const #(
		.value(8'h01),
		.width(8)
	) const_1_8(.out(const_1_8_out));
	coreir_eq #(.width(8)) coreir_eq_8_inst0(
		.in0(I),
		.in1(const_1_8_out),
		.out(coreir_eq_8_inst0_out)
	);
	assign O = coreir_eq_8_inst0_out;
endmodule
module Decode158 (
	I,
	O
);
	input [7:0] I;
	output wire O;
	wire [7:0] const_15_8_out;
	wire coreir_eq_8_inst0_out;
	coreir_const #(
		.value(8'h0f),
		.width(8)
	) const_15_8(.out(const_15_8_out));
	coreir_eq #(.width(8)) coreir_eq_8_inst0(
		.in0(I),
		.in1(const_15_8_out),
		.out(coreir_eq_8_inst0_out)
	);
	assign O = coreir_eq_8_inst0_out;
endmodule
module Decode148 (
	I,
	O
);
	input [7:0] I;
	output wire O;
	wire [7:0] const_14_8_out;
	wire coreir_eq_8_inst0_out;
	coreir_const #(
		.value(8'h0e),
		.width(8)
	) const_14_8(.out(const_14_8_out));
	coreir_eq #(.width(8)) coreir_eq_8_inst0(
		.in0(I),
		.in1(const_14_8_out),
		.out(coreir_eq_8_inst0_out)
	);
	assign O = coreir_eq_8_inst0_out;
endmodule
module Decode138 (
	I,
	O
);
	input [7:0] I;
	output wire O;
	wire [7:0] const_13_8_out;
	wire coreir_eq_8_inst0_out;
	coreir_const #(
		.value(8'h0d),
		.width(8)
	) const_13_8(.out(const_13_8_out));
	coreir_eq #(.width(8)) coreir_eq_8_inst0(
		.in0(I),
		.in1(const_13_8_out),
		.out(coreir_eq_8_inst0_out)
	);
	assign O = coreir_eq_8_inst0_out;
endmodule
module Decode128 (
	I,
	O
);
	input [7:0] I;
	output wire O;
	wire [7:0] const_12_8_out;
	wire coreir_eq_8_inst0_out;
	coreir_const #(
		.value(8'h0c),
		.width(8)
	) const_12_8(.out(const_12_8_out));
	coreir_eq #(.width(8)) coreir_eq_8_inst0(
		.in0(I),
		.in1(const_12_8_out),
		.out(coreir_eq_8_inst0_out)
	);
	assign O = coreir_eq_8_inst0_out;
endmodule
module Decode118 (
	I,
	O
);
	input [7:0] I;
	output wire O;
	wire [7:0] const_11_8_out;
	wire coreir_eq_8_inst0_out;
	coreir_const #(
		.value(8'h0b),
		.width(8)
	) const_11_8(.out(const_11_8_out));
	coreir_eq #(.width(8)) coreir_eq_8_inst0(
		.in0(I),
		.in1(const_11_8_out),
		.out(coreir_eq_8_inst0_out)
	);
	assign O = coreir_eq_8_inst0_out;
endmodule
module Decode108 (
	I,
	O
);
	input [7:0] I;
	output wire O;
	wire [7:0] const_10_8_out;
	wire coreir_eq_8_inst0_out;
	coreir_const #(
		.value(8'h0a),
		.width(8)
	) const_10_8(.out(const_10_8_out));
	coreir_eq #(.width(8)) coreir_eq_8_inst0(
		.in0(I),
		.in1(const_10_8_out),
		.out(coreir_eq_8_inst0_out)
	);
	assign O = coreir_eq_8_inst0_out;
endmodule
module Decode08 (
	I,
	O
);
	input [7:0] I;
	output wire O;
	wire [7:0] const_0_8_out;
	wire coreir_eq_8_inst0_out;
	coreir_const #(
		.value(8'h00),
		.width(8)
	) const_0_8(.out(const_0_8_out));
	coreir_eq #(.width(8)) coreir_eq_8_inst0(
		.in0(I),
		.in1(const_0_8_out),
		.out(coreir_eq_8_inst0_out)
	);
	assign O = coreir_eq_8_inst0_out;
endmodule
module ConfigRegister_6_8_32_0 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [5:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [5:0] Register_inst0_O;
	wire [7:0] const_0_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq2 Register_inst0(
		.I(config_data[5:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h00),
		.width(8)
	) const_0_8(.out(const_0_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_0_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_9 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_9_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h09),
		.width(8)
	) const_9_8(.out(const_9_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_9_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_8 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_8_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h08),
		.width(8)
	) const_8_8(.out(const_8_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_8_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_7 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_7_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h07),
		.width(8)
	) const_7_8(.out(const_7_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_7_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_6 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_6_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h06),
		.width(8)
	) const_6_8(.out(const_6_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_6_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_5 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_5_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h05),
		.width(8)
	) const_5_8(.out(const_5_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_5_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_45 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_45_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h2d),
		.width(8)
	) const_45_8(.out(const_45_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_45_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_44 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_44_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h2c),
		.width(8)
	) const_44_8(.out(const_44_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_44_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_43 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_43_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h2b),
		.width(8)
	) const_43_8(.out(const_43_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_43_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_42 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_42_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h2a),
		.width(8)
	) const_42_8(.out(const_42_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_42_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_41 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_41_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h29),
		.width(8)
	) const_41_8(.out(const_41_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_41_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_4 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_4_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h04),
		.width(8)
	) const_4_8(.out(const_4_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_4_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_39 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_39_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h27),
		.width(8)
	) const_39_8(.out(const_39_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_39_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_38 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_38_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h26),
		.width(8)
	) const_38_8(.out(const_38_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_38_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_37 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_37_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h25),
		.width(8)
	) const_37_8(.out(const_37_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_37_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_36 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_36_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h24),
		.width(8)
	) const_36_8(.out(const_36_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_36_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_35 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_35_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h23),
		.width(8)
	) const_35_8(.out(const_35_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_35_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_34 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_34_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h22),
		.width(8)
	) const_34_8(.out(const_34_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_34_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_33 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_33_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h21),
		.width(8)
	) const_33_8(.out(const_33_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_33_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_32 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_32_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h20),
		.width(8)
	) const_32_8(.out(const_32_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_32_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_31 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_31_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h1f),
		.width(8)
	) const_31_8(.out(const_31_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_31_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_30 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_30_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h1e),
		.width(8)
	) const_30_8(.out(const_30_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_30_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_3 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_3_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h03),
		.width(8)
	) const_3_8(.out(const_3_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_3_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_29 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_29_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h1d),
		.width(8)
	) const_29_8(.out(const_29_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_29_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_28 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_28_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h1c),
		.width(8)
	) const_28_8(.out(const_28_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_28_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_27 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_27_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h1b),
		.width(8)
	) const_27_8(.out(const_27_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_27_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_26 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_26_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h1a),
		.width(8)
	) const_26_8(.out(const_26_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_26_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_25 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_25_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h19),
		.width(8)
	) const_25_8(.out(const_25_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_25_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_24 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_24_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h18),
		.width(8)
	) const_24_8(.out(const_24_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_24_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_23 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_23_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h17),
		.width(8)
	) const_23_8(.out(const_23_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_23_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_22 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_22_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h16),
		.width(8)
	) const_22_8(.out(const_22_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_22_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_21 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_21_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h15),
		.width(8)
	) const_21_8(.out(const_21_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_21_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_20 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_20_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h14),
		.width(8)
	) const_20_8(.out(const_20_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_20_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_2 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_2_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h02),
		.width(8)
	) const_2_8(.out(const_2_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_2_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_19 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_19_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h13),
		.width(8)
	) const_19_8(.out(const_19_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_19_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_18 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_18_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h12),
		.width(8)
	) const_18_8(.out(const_18_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_18_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_17 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_17_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h11),
		.width(8)
	) const_17_8(.out(const_17_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_17_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_16 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_16_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h10),
		.width(8)
	) const_16_8(.out(const_16_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_16_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_15 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_15_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h0f),
		.width(8)
	) const_15_8(.out(const_15_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_15_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_14 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_14_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h0e),
		.width(8)
	) const_14_8(.out(const_14_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_14_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_13 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_13_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h0d),
		.width(8)
	) const_13_8(.out(const_13_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_13_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_12 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_12_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h0c),
		.width(8)
	) const_12_8(.out(const_12_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_12_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_11 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_11_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h0b),
		.width(8)
	) const_11_8(.out(const_11_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_11_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_10 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_10_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h0a),
		.width(8)
	) const_10_8(.out(const_10_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_10_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_1 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_1_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h01),
		.width(8)
	) const_1_8(.out(const_1_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_1_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_0 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_0_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h00),
		.width(8)
	) const_0_8(.out(const_0_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_0_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_31_8_32_3 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [30:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [30:0] Register_inst0_O;
	wire [7:0] const_3_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq5 Register_inst0(
		.I(config_data[30:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h03),
		.width(8)
	) const_3_8(.out(const_3_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_3_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_30_8_32_8 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [29:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [29:0] Register_inst0_O;
	wire [7:0] const_8_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data[29:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h08),
		.width(8)
	) const_8_8(.out(const_8_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_8_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_30_8_32_4 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [29:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [29:0] Register_inst0_O;
	wire [7:0] const_4_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data[29:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h04),
		.width(8)
	) const_4_8(.out(const_4_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_4_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_25_8_32_46 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [24:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [24:0] Register_inst0_O;
	wire [7:0] const_46_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq8 Register_inst0(
		.I(config_data[24:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h2e),
		.width(8)
	) const_46_8(.out(const_46_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_46_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_24_8_32_0 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [23:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [23:0] Register_inst0_O;
	wire [7:0] const_0_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq9 Register_inst0(
		.I(config_data[23:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h00),
		.width(8)
	) const_0_8(.out(const_0_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_0_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module IOCoreReadyValid (
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	f2io_1,
	f2io_17,
	f2io_17_ready,
	f2io_17_valid,
	f2io_1_ready,
	f2io_1_valid,
	flush,
	flush_core,
	glb2io_1,
	glb2io_17,
	glb2io_17_ready,
	glb2io_17_valid,
	glb2io_1_ready,
	glb2io_1_valid,
	io2f_1,
	io2f_17,
	io2f_17_ready,
	io2f_17_valid,
	io2f_1_ready,
	io2f_1_valid,
	io2glb_1,
	io2glb_17,
	io2glb_17_ready,
	io2glb_17_valid,
	io2glb_1_ready,
	io2glb_1_valid,
	read_config_data,
	reset,
	stall
);
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	input [0:0] f2io_1;
	input [16:0] f2io_17;
	output wire [0:0] f2io_17_ready;
	input [0:0] f2io_17_valid;
	output wire [0:0] f2io_1_ready;
	input [0:0] f2io_1_valid;
	input [0:0] flush;
	input [0:0] flush_core;
	input [0:0] glb2io_1;
	input [16:0] glb2io_17;
	output wire [0:0] glb2io_17_ready;
	input [0:0] glb2io_17_valid;
	output wire [0:0] glb2io_1_ready;
	input [0:0] glb2io_1_valid;
	output wire [0:0] io2f_1;
	output wire [16:0] io2f_17;
	input [0:0] io2f_17_ready;
	output wire [0:0] io2f_17_valid;
	input [0:0] io2f_1_ready;
	output wire [0:0] io2f_1_valid;
	output wire [0:0] io2glb_1;
	output wire [16:0] io2glb_17;
	input [0:0] io2glb_17_ready;
	output wire [0:0] io2glb_17_valid;
	input [0:0] io2glb_1_ready;
	output wire [0:0] io2glb_1_valid;
	output wire [31:0] read_config_data;
	input reset;
	input [0:0] stall;
	wire [0:0] Invert1_inst0_out;
	wire [0:0] Invert1_inst1_out;
	wire ZextWrapper_24_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_24_32_inst0$self_O_in;
	wire [23:0] config_reg_0_O;
	wire coreir_wrapInAsyncReset_inst0_out;
	wire coreir_wrapOutAsyncReset_inst0_out;
	wire [0:0] f2io_17_valid_reg_sel_value_O;
	wire [0:0] f2io_17_valid_reg_value_value_O;
	wire [0:0] f2io_17_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] f2io_1_reg_sel_value_O;
	wire [0:0] f2io_1_reg_value_value_O;
	wire [0:0] f2io_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] f2io_1_valid_reg_sel_value_O;
	wire [0:0] f2io_1_valid_reg_value_value_O;
	wire [0:0] f2io_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] flush_mux_sel_value_O;
	wire [0:0] flush_reg_sel_value_O;
	wire [0:0] flush_reg_value_value_O;
	wire [0:0] flush_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] glb2io_17_valid_reg_sel_value_O;
	wire [0:0] glb2io_17_valid_reg_value_value_O;
	wire [0:0] glb2io_17_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] glb2io_1_reg_sel_value_O;
	wire [0:0] glb2io_1_reg_value_value_O;
	wire [0:0] glb2io_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] glb2io_1_valid_reg_sel_value_O;
	wire [0:0] glb2io_1_valid_reg_value_value_O;
	wire [0:0] glb2io_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] io2f_17_ready_reg_sel_value_O;
	wire [0:0] io2f_17_ready_reg_value_value_O;
	wire [0:0] io2f_17_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] io2f_1_ready_reg_sel_value_O;
	wire [0:0] io2f_1_ready_reg_value_value_O;
	wire [0:0] io2f_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] io2glb_17_ready_reg_sel_value_O;
	wire [0:0] io2glb_17_ready_reg_value_value_O;
	wire [0:0] io2glb_17_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] io2glb_1_ready_reg_sel_value_O;
	wire [0:0] io2glb_1_ready_reg_value_value_O;
	wire [0:0] io2glb_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] io_core_W_inst0_io2glb_17_valid;
	wire [0:0] io_core_W_inst0_f2io_1_ready;
	wire [0:0] io_core_W_inst0_glb2io_17_ready;
	wire [0:0] io_core_W_inst0_io2glb_1_valid;
	wire [0:0] io_core_W_inst0_io2glb_1;
	wire [0:0] io_core_W_inst0_glb2io_1_ready;
	wire [16:0] io_core_W_inst0_io2glb_17;
	wire [0:0] io_core_W_inst0_io2f_1;
	wire [16:0] io_core_W_inst0_io2f_17;
	wire [0:0] io_core_W_inst0_f2io_17_ready;
	wire [0:0] io_core_W_inst0_io2f_1_valid;
	wire [0:0] io_core_W_inst0_io2f_17_valid;
	wire [0:0] tile_en_value_O;
	coreir_not #(.width(1)) Invert1_inst0(
		.in(coreir_wrapInAsyncReset_inst0_out),
		.out(Invert1_inst0_out)
	);
	coreir_not #(.width(1)) Invert1_inst1(
		.in(stall),
		.out(Invert1_inst1_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_24_32_inst0$bit_const_0_None(.out(ZextWrapper_24_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_24_32_inst0$self_O_out;
	assign ZextWrapper_24_32_inst0$self_O_out = {ZextWrapper_24_32_inst0$bit_const_0_None_out, ZextWrapper_24_32_inst0$bit_const_0_None_out, ZextWrapper_24_32_inst0$bit_const_0_None_out, ZextWrapper_24_32_inst0$bit_const_0_None_out, ZextWrapper_24_32_inst0$bit_const_0_None_out, ZextWrapper_24_32_inst0$bit_const_0_None_out, ZextWrapper_24_32_inst0$bit_const_0_None_out, ZextWrapper_24_32_inst0$bit_const_0_None_out, config_reg_0_O};
	mantle_wire__typeBitIn32 ZextWrapper_24_32_inst0$self_O(
		.in(ZextWrapper_24_32_inst0$self_O_in),
		.out(ZextWrapper_24_32_inst0$self_O_out)
	);
	ConfigRegister_24_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	coreir_wrap coreir_wrapInAsyncReset_inst0(
		.in(reset),
		.out(coreir_wrapInAsyncReset_inst0_out)
	);
	coreir_wrap coreir_wrapOutAsyncReset_inst0(
		.in(Invert1_inst0_out[0]),
		.out(coreir_wrapOutAsyncReset_inst0_out)
	);
	SliceWrapper_24_0_1 f2io_17_valid_reg_sel_value(
		.I(config_reg_0_O),
		.O(f2io_17_valid_reg_sel_value_O)
	);
	SliceWrapper_24_1_2 f2io_17_valid_reg_value_value(
		.I(config_reg_0_O),
		.O(f2io_17_valid_reg_value_value_O)
	);
	coreir_mux #(.width(1)) f2io_17_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(f2io_17_valid),
		.in1(f2io_17_valid_reg_value_value_O),
		.sel(f2io_17_valid_reg_sel_value_O[0]),
		.out(f2io_17_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_24_2_3 f2io_1_reg_sel_value(
		.I(config_reg_0_O),
		.O(f2io_1_reg_sel_value_O)
	);
	SliceWrapper_24_3_4 f2io_1_reg_value_value(
		.I(config_reg_0_O),
		.O(f2io_1_reg_value_value_O)
	);
	coreir_mux #(.width(1)) f2io_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(f2io_1),
		.in1(f2io_1_reg_value_value_O),
		.sel(f2io_1_reg_sel_value_O[0]),
		.out(f2io_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_24_4_5 f2io_1_valid_reg_sel_value(
		.I(config_reg_0_O),
		.O(f2io_1_valid_reg_sel_value_O)
	);
	SliceWrapper_24_5_6 f2io_1_valid_reg_value_value(
		.I(config_reg_0_O),
		.O(f2io_1_valid_reg_value_value_O)
	);
	coreir_mux #(.width(1)) f2io_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(f2io_1_valid),
		.in1(f2io_1_valid_reg_value_value_O),
		.sel(f2io_1_valid_reg_sel_value_O[0]),
		.out(f2io_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(flush_core),
		.in1(flush),
		.sel(flush_mux_sel_value_O[0]),
		.out(flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_24_6_7 flush_mux_sel_value(
		.I(config_reg_0_O),
		.O(flush_mux_sel_value_O)
	);
	SliceWrapper_24_7_8 flush_reg_sel_value(
		.I(config_reg_0_O),
		.O(flush_reg_sel_value_O)
	);
	SliceWrapper_24_8_9 flush_reg_value_value(
		.I(config_reg_0_O),
		.O(flush_reg_value_value_O)
	);
	coreir_mux #(.width(1)) flush_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(flush),
		.in1(flush_reg_value_value_O),
		.sel(flush_reg_sel_value_O[0]),
		.out(flush_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_24_9_10 glb2io_17_valid_reg_sel_value(
		.I(config_reg_0_O),
		.O(glb2io_17_valid_reg_sel_value_O)
	);
	SliceWrapper_24_10_11 glb2io_17_valid_reg_value_value(
		.I(config_reg_0_O),
		.O(glb2io_17_valid_reg_value_value_O)
	);
	coreir_mux #(.width(1)) glb2io_17_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(glb2io_17_valid),
		.in1(glb2io_17_valid_reg_value_value_O),
		.sel(glb2io_17_valid_reg_sel_value_O[0]),
		.out(glb2io_17_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_24_11_12 glb2io_1_reg_sel_value(
		.I(config_reg_0_O),
		.O(glb2io_1_reg_sel_value_O)
	);
	SliceWrapper_24_12_13 glb2io_1_reg_value_value(
		.I(config_reg_0_O),
		.O(glb2io_1_reg_value_value_O)
	);
	coreir_mux #(.width(1)) glb2io_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(glb2io_1),
		.in1(glb2io_1_reg_value_value_O),
		.sel(glb2io_1_reg_sel_value_O[0]),
		.out(glb2io_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_24_13_14 glb2io_1_valid_reg_sel_value(
		.I(config_reg_0_O),
		.O(glb2io_1_valid_reg_sel_value_O)
	);
	SliceWrapper_24_14_15 glb2io_1_valid_reg_value_value(
		.I(config_reg_0_O),
		.O(glb2io_1_valid_reg_value_value_O)
	);
	coreir_mux #(.width(1)) glb2io_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(glb2io_1_valid),
		.in1(glb2io_1_valid_reg_value_value_O),
		.sel(glb2io_1_valid_reg_sel_value_O[0]),
		.out(glb2io_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_24_15_16 io2f_17_ready_reg_sel_value(
		.I(config_reg_0_O),
		.O(io2f_17_ready_reg_sel_value_O)
	);
	SliceWrapper_24_16_17 io2f_17_ready_reg_value_value(
		.I(config_reg_0_O),
		.O(io2f_17_ready_reg_value_value_O)
	);
	coreir_mux #(.width(1)) io2f_17_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(io2f_17_ready),
		.in1(io2f_17_ready_reg_value_value_O),
		.sel(io2f_17_ready_reg_sel_value_O[0]),
		.out(io2f_17_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_24_17_18 io2f_1_ready_reg_sel_value(
		.I(config_reg_0_O),
		.O(io2f_1_ready_reg_sel_value_O)
	);
	SliceWrapper_24_18_19 io2f_1_ready_reg_value_value(
		.I(config_reg_0_O),
		.O(io2f_1_ready_reg_value_value_O)
	);
	coreir_mux #(.width(1)) io2f_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(io2f_1_ready),
		.in1(io2f_1_ready_reg_value_value_O),
		.sel(io2f_1_ready_reg_sel_value_O[0]),
		.out(io2f_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_24_19_20 io2glb_17_ready_reg_sel_value(
		.I(config_reg_0_O),
		.O(io2glb_17_ready_reg_sel_value_O)
	);
	SliceWrapper_24_20_21 io2glb_17_ready_reg_value_value(
		.I(config_reg_0_O),
		.O(io2glb_17_ready_reg_value_value_O)
	);
	coreir_mux #(.width(1)) io2glb_17_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(io2glb_17_ready),
		.in1(io2glb_17_ready_reg_value_value_O),
		.sel(io2glb_17_ready_reg_sel_value_O[0]),
		.out(io2glb_17_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_24_21_22 io2glb_1_ready_reg_sel_value(
		.I(config_reg_0_O),
		.O(io2glb_1_ready_reg_sel_value_O)
	);
	SliceWrapper_24_22_23 io2glb_1_ready_reg_value_value(
		.I(config_reg_0_O),
		.O(io2glb_1_ready_reg_value_value_O)
	);
	coreir_mux #(.width(1)) io2glb_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(io2glb_1_ready),
		.in1(io2glb_1_ready_reg_value_value_O),
		.sel(io2glb_1_ready_reg_sel_value_O[0]),
		.out(io2glb_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	io_core_W io_core_W_inst0(
		.io2glb_1_ready(io2glb_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.io2glb_17_ready(io2glb_17_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.clk_en(Invert1_inst1_out),
		.io2f_1_ready(io2f_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.io2glb_17_valid(io_core_W_inst0_io2glb_17_valid),
		.io2f_17_ready(io2f_17_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.f2io_17(f2io_17),
		.f2io_1_ready(io_core_W_inst0_f2io_1_ready),
		.glb2io_17_ready(io_core_W_inst0_glb2io_17_ready),
		.io2glb_1_valid(io_core_W_inst0_io2glb_1_valid),
		.tile_en(tile_en_value_O),
		.glb2io_17_valid(glb2io_17_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.io2glb_1(io_core_W_inst0_io2glb_1),
		.clk(clk),
		.flush(flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.glb2io_1_valid(glb2io_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.glb2io_1_ready(io_core_W_inst0_glb2io_1_ready),
		.f2io_1(f2io_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.io2glb_17(io_core_W_inst0_io2glb_17),
		.f2io_1_valid(f2io_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.io2f_1(io_core_W_inst0_io2f_1),
		.io2f_17(io_core_W_inst0_io2f_17),
		.f2io_17_ready(io_core_W_inst0_f2io_17_ready),
		.glb2io_17(glb2io_17),
		.io2f_1_valid(io_core_W_inst0_io2f_1_valid),
		.f2io_17_valid(f2io_17_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.glb2io_1(glb2io_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.io2f_17_valid(io_core_W_inst0_io2f_17_valid),
		.rst_n(coreir_wrapOutAsyncReset_inst0_out)
	);
	SliceWrapper_24_23_24 tile_en_value(
		.I(config_reg_0_O),
		.O(tile_en_value_O)
	);
	assign f2io_17_ready = io_core_W_inst0_f2io_17_ready;
	assign f2io_1_ready = io_core_W_inst0_f2io_1_ready;
	assign glb2io_17_ready = io_core_W_inst0_glb2io_17_ready;
	assign glb2io_1_ready = io_core_W_inst0_glb2io_1_ready;
	assign io2f_1 = io_core_W_inst0_io2f_1;
	assign io2f_17 = io_core_W_inst0_io2f_17;
	assign io2f_17_valid = io_core_W_inst0_io2f_17_valid;
	assign io2f_1_valid = io_core_W_inst0_io2f_1_valid;
	assign io2glb_1 = io_core_W_inst0_io2glb_1;
	assign io2glb_17 = io_core_W_inst0_io2glb_17;
	assign io2glb_17_valid = io_core_W_inst0_io2glb_17_valid;
	assign io2glb_1_valid = io_core_W_inst0_io2glb_1_valid;
	assign read_config_data = ZextWrapper_24_32_inst0$self_O_in;
endmodule
module ConfigRegister_23_8_32_5 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [22:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [22:0] Register_inst0_O;
	wire [7:0] const_5_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq6 Register_inst0(
		.I(config_data[22:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h05),
		.width(8)
	) const_5_8(.out(const_5_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_5_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module SB_ID0_5TRACKS_B1_PE (
	PE_input_width_1_num_0_enable,
	PE_input_width_1_num_0_out_sel,
	PE_input_width_1_num_0_ready,
	PE_input_width_1_num_1_enable,
	PE_input_width_1_num_1_out_sel,
	PE_input_width_1_num_1_ready,
	PE_input_width_1_num_2_enable,
	PE_input_width_1_num_2_out_sel,
	PE_input_width_1_num_2_ready,
	PE_output_width_1_num_0,
	PE_output_width_1_num_0_ready_out,
	PE_output_width_1_num_0_valid,
	PondTop_output_width_1_num_0,
	PondTop_output_width_1_num_0_ready_out,
	PondTop_output_width_1_num_0_valid,
	PondTop_output_width_1_num_1,
	PondTop_output_width_1_num_1_ready_out,
	PondTop_output_width_1_num_1_valid,
	SB_T0_EAST_SB_IN_B1,
	SB_T0_EAST_SB_IN_B1_enable,
	SB_T0_EAST_SB_IN_B1_ready_out,
	SB_T0_EAST_SB_IN_B1_valid_in,
	SB_T0_EAST_SB_OUT_B1,
	SB_T0_EAST_SB_OUT_B1_enable,
	SB_T0_EAST_SB_OUT_B1_ready_in,
	SB_T0_EAST_SB_OUT_B1_valid_out,
	SB_T0_NORTH_SB_IN_B1,
	SB_T0_NORTH_SB_IN_B1_enable,
	SB_T0_NORTH_SB_IN_B1_ready_out,
	SB_T0_NORTH_SB_IN_B1_valid_in,
	SB_T0_NORTH_SB_OUT_B1,
	SB_T0_NORTH_SB_OUT_B1_enable,
	SB_T0_NORTH_SB_OUT_B1_ready_in,
	SB_T0_NORTH_SB_OUT_B1_valid_out,
	SB_T0_SOUTH_SB_IN_B1,
	SB_T0_SOUTH_SB_IN_B1_enable,
	SB_T0_SOUTH_SB_IN_B1_ready_out,
	SB_T0_SOUTH_SB_IN_B1_valid_in,
	SB_T0_SOUTH_SB_OUT_B1,
	SB_T0_SOUTH_SB_OUT_B1_enable,
	SB_T0_SOUTH_SB_OUT_B1_ready_in,
	SB_T0_SOUTH_SB_OUT_B1_valid_out,
	SB_T0_WEST_SB_IN_B1,
	SB_T0_WEST_SB_IN_B1_enable,
	SB_T0_WEST_SB_IN_B1_ready_out,
	SB_T0_WEST_SB_IN_B1_valid_in,
	SB_T0_WEST_SB_OUT_B1,
	SB_T0_WEST_SB_OUT_B1_enable,
	SB_T0_WEST_SB_OUT_B1_ready_in,
	SB_T0_WEST_SB_OUT_B1_valid_out,
	SB_T1_EAST_SB_IN_B1,
	SB_T1_EAST_SB_IN_B1_enable,
	SB_T1_EAST_SB_IN_B1_ready_out,
	SB_T1_EAST_SB_IN_B1_valid_in,
	SB_T1_EAST_SB_OUT_B1,
	SB_T1_EAST_SB_OUT_B1_enable,
	SB_T1_EAST_SB_OUT_B1_ready_in,
	SB_T1_EAST_SB_OUT_B1_valid_out,
	SB_T1_NORTH_SB_IN_B1,
	SB_T1_NORTH_SB_IN_B1_enable,
	SB_T1_NORTH_SB_IN_B1_ready_out,
	SB_T1_NORTH_SB_IN_B1_valid_in,
	SB_T1_NORTH_SB_OUT_B1,
	SB_T1_NORTH_SB_OUT_B1_enable,
	SB_T1_NORTH_SB_OUT_B1_ready_in,
	SB_T1_NORTH_SB_OUT_B1_valid_out,
	SB_T1_SOUTH_SB_IN_B1,
	SB_T1_SOUTH_SB_IN_B1_enable,
	SB_T1_SOUTH_SB_IN_B1_ready_out,
	SB_T1_SOUTH_SB_IN_B1_valid_in,
	SB_T1_SOUTH_SB_OUT_B1,
	SB_T1_SOUTH_SB_OUT_B1_enable,
	SB_T1_SOUTH_SB_OUT_B1_ready_in,
	SB_T1_SOUTH_SB_OUT_B1_valid_out,
	SB_T1_WEST_SB_IN_B1,
	SB_T1_WEST_SB_IN_B1_enable,
	SB_T1_WEST_SB_IN_B1_ready_out,
	SB_T1_WEST_SB_IN_B1_valid_in,
	SB_T1_WEST_SB_OUT_B1,
	SB_T1_WEST_SB_OUT_B1_enable,
	SB_T1_WEST_SB_OUT_B1_ready_in,
	SB_T1_WEST_SB_OUT_B1_valid_out,
	SB_T2_EAST_SB_IN_B1,
	SB_T2_EAST_SB_IN_B1_enable,
	SB_T2_EAST_SB_IN_B1_ready_out,
	SB_T2_EAST_SB_IN_B1_valid_in,
	SB_T2_EAST_SB_OUT_B1,
	SB_T2_EAST_SB_OUT_B1_enable,
	SB_T2_EAST_SB_OUT_B1_ready_in,
	SB_T2_EAST_SB_OUT_B1_valid_out,
	SB_T2_NORTH_SB_IN_B1,
	SB_T2_NORTH_SB_IN_B1_enable,
	SB_T2_NORTH_SB_IN_B1_ready_out,
	SB_T2_NORTH_SB_IN_B1_valid_in,
	SB_T2_NORTH_SB_OUT_B1,
	SB_T2_NORTH_SB_OUT_B1_enable,
	SB_T2_NORTH_SB_OUT_B1_ready_in,
	SB_T2_NORTH_SB_OUT_B1_valid_out,
	SB_T2_SOUTH_SB_IN_B1,
	SB_T2_SOUTH_SB_IN_B1_enable,
	SB_T2_SOUTH_SB_IN_B1_ready_out,
	SB_T2_SOUTH_SB_IN_B1_valid_in,
	SB_T2_SOUTH_SB_OUT_B1,
	SB_T2_SOUTH_SB_OUT_B1_enable,
	SB_T2_SOUTH_SB_OUT_B1_ready_in,
	SB_T2_SOUTH_SB_OUT_B1_valid_out,
	SB_T2_WEST_SB_IN_B1,
	SB_T2_WEST_SB_IN_B1_enable,
	SB_T2_WEST_SB_IN_B1_ready_out,
	SB_T2_WEST_SB_IN_B1_valid_in,
	SB_T2_WEST_SB_OUT_B1,
	SB_T2_WEST_SB_OUT_B1_enable,
	SB_T2_WEST_SB_OUT_B1_ready_in,
	SB_T2_WEST_SB_OUT_B1_valid_out,
	SB_T3_EAST_SB_IN_B1,
	SB_T3_EAST_SB_IN_B1_enable,
	SB_T3_EAST_SB_IN_B1_ready_out,
	SB_T3_EAST_SB_IN_B1_valid_in,
	SB_T3_EAST_SB_OUT_B1,
	SB_T3_EAST_SB_OUT_B1_enable,
	SB_T3_EAST_SB_OUT_B1_ready_in,
	SB_T3_EAST_SB_OUT_B1_valid_out,
	SB_T3_NORTH_SB_IN_B1,
	SB_T3_NORTH_SB_IN_B1_enable,
	SB_T3_NORTH_SB_IN_B1_ready_out,
	SB_T3_NORTH_SB_IN_B1_valid_in,
	SB_T3_NORTH_SB_OUT_B1,
	SB_T3_NORTH_SB_OUT_B1_enable,
	SB_T3_NORTH_SB_OUT_B1_ready_in,
	SB_T3_NORTH_SB_OUT_B1_valid_out,
	SB_T3_SOUTH_SB_IN_B1,
	SB_T3_SOUTH_SB_IN_B1_enable,
	SB_T3_SOUTH_SB_IN_B1_ready_out,
	SB_T3_SOUTH_SB_IN_B1_valid_in,
	SB_T3_SOUTH_SB_OUT_B1,
	SB_T3_SOUTH_SB_OUT_B1_enable,
	SB_T3_SOUTH_SB_OUT_B1_ready_in,
	SB_T3_SOUTH_SB_OUT_B1_valid_out,
	SB_T3_WEST_SB_IN_B1,
	SB_T3_WEST_SB_IN_B1_enable,
	SB_T3_WEST_SB_IN_B1_ready_out,
	SB_T3_WEST_SB_IN_B1_valid_in,
	SB_T3_WEST_SB_OUT_B1,
	SB_T3_WEST_SB_OUT_B1_enable,
	SB_T3_WEST_SB_OUT_B1_ready_in,
	SB_T3_WEST_SB_OUT_B1_valid_out,
	SB_T4_EAST_SB_IN_B1,
	SB_T4_EAST_SB_IN_B1_enable,
	SB_T4_EAST_SB_IN_B1_ready_out,
	SB_T4_EAST_SB_IN_B1_valid_in,
	SB_T4_EAST_SB_OUT_B1,
	SB_T4_EAST_SB_OUT_B1_enable,
	SB_T4_EAST_SB_OUT_B1_ready_in,
	SB_T4_EAST_SB_OUT_B1_valid_out,
	SB_T4_NORTH_SB_IN_B1,
	SB_T4_NORTH_SB_IN_B1_enable,
	SB_T4_NORTH_SB_IN_B1_ready_out,
	SB_T4_NORTH_SB_IN_B1_valid_in,
	SB_T4_NORTH_SB_OUT_B1,
	SB_T4_NORTH_SB_OUT_B1_enable,
	SB_T4_NORTH_SB_OUT_B1_ready_in,
	SB_T4_NORTH_SB_OUT_B1_valid_out,
	SB_T4_SOUTH_SB_IN_B1,
	SB_T4_SOUTH_SB_IN_B1_enable,
	SB_T4_SOUTH_SB_IN_B1_ready_out,
	SB_T4_SOUTH_SB_IN_B1_valid_in,
	SB_T4_SOUTH_SB_OUT_B1,
	SB_T4_SOUTH_SB_OUT_B1_enable,
	SB_T4_SOUTH_SB_OUT_B1_ready_in,
	SB_T4_SOUTH_SB_OUT_B1_valid_out,
	SB_T4_WEST_SB_IN_B1,
	SB_T4_WEST_SB_IN_B1_enable,
	SB_T4_WEST_SB_IN_B1_ready_out,
	SB_T4_WEST_SB_IN_B1_valid_in,
	SB_T4_WEST_SB_OUT_B1,
	SB_T4_WEST_SB_OUT_B1_enable,
	SB_T4_WEST_SB_OUT_B1_ready_in,
	SB_T4_WEST_SB_OUT_B1_valid_out,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	read_config_data,
	reset,
	stall
);
	input [0:0] PE_input_width_1_num_0_enable;
	input [31:0] PE_input_width_1_num_0_out_sel;
	input PE_input_width_1_num_0_ready;
	input [0:0] PE_input_width_1_num_1_enable;
	input [31:0] PE_input_width_1_num_1_out_sel;
	input PE_input_width_1_num_1_ready;
	input [0:0] PE_input_width_1_num_2_enable;
	input [31:0] PE_input_width_1_num_2_out_sel;
	input PE_input_width_1_num_2_ready;
	input [0:0] PE_output_width_1_num_0;
	output wire PE_output_width_1_num_0_ready_out;
	input PE_output_width_1_num_0_valid;
	input [0:0] PondTop_output_width_1_num_0;
	output wire PondTop_output_width_1_num_0_ready_out;
	input PondTop_output_width_1_num_0_valid;
	input [0:0] PondTop_output_width_1_num_1;
	output wire PondTop_output_width_1_num_1_ready_out;
	input PondTop_output_width_1_num_1_valid;
	input [0:0] SB_T0_EAST_SB_IN_B1;
	output wire SB_T0_EAST_SB_IN_B1_enable;
	output wire SB_T0_EAST_SB_IN_B1_ready_out;
	input SB_T0_EAST_SB_IN_B1_valid_in;
	output wire [0:0] SB_T0_EAST_SB_OUT_B1;
	output wire SB_T0_EAST_SB_OUT_B1_enable;
	input SB_T0_EAST_SB_OUT_B1_ready_in;
	output wire SB_T0_EAST_SB_OUT_B1_valid_out;
	input [0:0] SB_T0_NORTH_SB_IN_B1;
	output wire SB_T0_NORTH_SB_IN_B1_enable;
	output wire SB_T0_NORTH_SB_IN_B1_ready_out;
	input SB_T0_NORTH_SB_IN_B1_valid_in;
	output wire [0:0] SB_T0_NORTH_SB_OUT_B1;
	output wire SB_T0_NORTH_SB_OUT_B1_enable;
	input SB_T0_NORTH_SB_OUT_B1_ready_in;
	output wire SB_T0_NORTH_SB_OUT_B1_valid_out;
	input [0:0] SB_T0_SOUTH_SB_IN_B1;
	output wire SB_T0_SOUTH_SB_IN_B1_enable;
	output wire SB_T0_SOUTH_SB_IN_B1_ready_out;
	input SB_T0_SOUTH_SB_IN_B1_valid_in;
	output wire [0:0] SB_T0_SOUTH_SB_OUT_B1;
	output wire SB_T0_SOUTH_SB_OUT_B1_enable;
	input SB_T0_SOUTH_SB_OUT_B1_ready_in;
	output wire SB_T0_SOUTH_SB_OUT_B1_valid_out;
	input [0:0] SB_T0_WEST_SB_IN_B1;
	output wire SB_T0_WEST_SB_IN_B1_enable;
	output wire SB_T0_WEST_SB_IN_B1_ready_out;
	input SB_T0_WEST_SB_IN_B1_valid_in;
	output wire [0:0] SB_T0_WEST_SB_OUT_B1;
	output wire SB_T0_WEST_SB_OUT_B1_enable;
	input SB_T0_WEST_SB_OUT_B1_ready_in;
	output wire SB_T0_WEST_SB_OUT_B1_valid_out;
	input [0:0] SB_T1_EAST_SB_IN_B1;
	output wire SB_T1_EAST_SB_IN_B1_enable;
	output wire SB_T1_EAST_SB_IN_B1_ready_out;
	input SB_T1_EAST_SB_IN_B1_valid_in;
	output wire [0:0] SB_T1_EAST_SB_OUT_B1;
	output wire SB_T1_EAST_SB_OUT_B1_enable;
	input SB_T1_EAST_SB_OUT_B1_ready_in;
	output wire SB_T1_EAST_SB_OUT_B1_valid_out;
	input [0:0] SB_T1_NORTH_SB_IN_B1;
	output wire SB_T1_NORTH_SB_IN_B1_enable;
	output wire SB_T1_NORTH_SB_IN_B1_ready_out;
	input SB_T1_NORTH_SB_IN_B1_valid_in;
	output wire [0:0] SB_T1_NORTH_SB_OUT_B1;
	output wire SB_T1_NORTH_SB_OUT_B1_enable;
	input SB_T1_NORTH_SB_OUT_B1_ready_in;
	output wire SB_T1_NORTH_SB_OUT_B1_valid_out;
	input [0:0] SB_T1_SOUTH_SB_IN_B1;
	output wire SB_T1_SOUTH_SB_IN_B1_enable;
	output wire SB_T1_SOUTH_SB_IN_B1_ready_out;
	input SB_T1_SOUTH_SB_IN_B1_valid_in;
	output wire [0:0] SB_T1_SOUTH_SB_OUT_B1;
	output wire SB_T1_SOUTH_SB_OUT_B1_enable;
	input SB_T1_SOUTH_SB_OUT_B1_ready_in;
	output wire SB_T1_SOUTH_SB_OUT_B1_valid_out;
	input [0:0] SB_T1_WEST_SB_IN_B1;
	output wire SB_T1_WEST_SB_IN_B1_enable;
	output wire SB_T1_WEST_SB_IN_B1_ready_out;
	input SB_T1_WEST_SB_IN_B1_valid_in;
	output wire [0:0] SB_T1_WEST_SB_OUT_B1;
	output wire SB_T1_WEST_SB_OUT_B1_enable;
	input SB_T1_WEST_SB_OUT_B1_ready_in;
	output wire SB_T1_WEST_SB_OUT_B1_valid_out;
	input [0:0] SB_T2_EAST_SB_IN_B1;
	output wire SB_T2_EAST_SB_IN_B1_enable;
	output wire SB_T2_EAST_SB_IN_B1_ready_out;
	input SB_T2_EAST_SB_IN_B1_valid_in;
	output wire [0:0] SB_T2_EAST_SB_OUT_B1;
	output wire SB_T2_EAST_SB_OUT_B1_enable;
	input SB_T2_EAST_SB_OUT_B1_ready_in;
	output wire SB_T2_EAST_SB_OUT_B1_valid_out;
	input [0:0] SB_T2_NORTH_SB_IN_B1;
	output wire SB_T2_NORTH_SB_IN_B1_enable;
	output wire SB_T2_NORTH_SB_IN_B1_ready_out;
	input SB_T2_NORTH_SB_IN_B1_valid_in;
	output wire [0:0] SB_T2_NORTH_SB_OUT_B1;
	output wire SB_T2_NORTH_SB_OUT_B1_enable;
	input SB_T2_NORTH_SB_OUT_B1_ready_in;
	output wire SB_T2_NORTH_SB_OUT_B1_valid_out;
	input [0:0] SB_T2_SOUTH_SB_IN_B1;
	output wire SB_T2_SOUTH_SB_IN_B1_enable;
	output wire SB_T2_SOUTH_SB_IN_B1_ready_out;
	input SB_T2_SOUTH_SB_IN_B1_valid_in;
	output wire [0:0] SB_T2_SOUTH_SB_OUT_B1;
	output wire SB_T2_SOUTH_SB_OUT_B1_enable;
	input SB_T2_SOUTH_SB_OUT_B1_ready_in;
	output wire SB_T2_SOUTH_SB_OUT_B1_valid_out;
	input [0:0] SB_T2_WEST_SB_IN_B1;
	output wire SB_T2_WEST_SB_IN_B1_enable;
	output wire SB_T2_WEST_SB_IN_B1_ready_out;
	input SB_T2_WEST_SB_IN_B1_valid_in;
	output wire [0:0] SB_T2_WEST_SB_OUT_B1;
	output wire SB_T2_WEST_SB_OUT_B1_enable;
	input SB_T2_WEST_SB_OUT_B1_ready_in;
	output wire SB_T2_WEST_SB_OUT_B1_valid_out;
	input [0:0] SB_T3_EAST_SB_IN_B1;
	output wire SB_T3_EAST_SB_IN_B1_enable;
	output wire SB_T3_EAST_SB_IN_B1_ready_out;
	input SB_T3_EAST_SB_IN_B1_valid_in;
	output wire [0:0] SB_T3_EAST_SB_OUT_B1;
	output wire SB_T3_EAST_SB_OUT_B1_enable;
	input SB_T3_EAST_SB_OUT_B1_ready_in;
	output wire SB_T3_EAST_SB_OUT_B1_valid_out;
	input [0:0] SB_T3_NORTH_SB_IN_B1;
	output wire SB_T3_NORTH_SB_IN_B1_enable;
	output wire SB_T3_NORTH_SB_IN_B1_ready_out;
	input SB_T3_NORTH_SB_IN_B1_valid_in;
	output wire [0:0] SB_T3_NORTH_SB_OUT_B1;
	output wire SB_T3_NORTH_SB_OUT_B1_enable;
	input SB_T3_NORTH_SB_OUT_B1_ready_in;
	output wire SB_T3_NORTH_SB_OUT_B1_valid_out;
	input [0:0] SB_T3_SOUTH_SB_IN_B1;
	output wire SB_T3_SOUTH_SB_IN_B1_enable;
	output wire SB_T3_SOUTH_SB_IN_B1_ready_out;
	input SB_T3_SOUTH_SB_IN_B1_valid_in;
	output wire [0:0] SB_T3_SOUTH_SB_OUT_B1;
	output wire SB_T3_SOUTH_SB_OUT_B1_enable;
	input SB_T3_SOUTH_SB_OUT_B1_ready_in;
	output wire SB_T3_SOUTH_SB_OUT_B1_valid_out;
	input [0:0] SB_T3_WEST_SB_IN_B1;
	output wire SB_T3_WEST_SB_IN_B1_enable;
	output wire SB_T3_WEST_SB_IN_B1_ready_out;
	input SB_T3_WEST_SB_IN_B1_valid_in;
	output wire [0:0] SB_T3_WEST_SB_OUT_B1;
	output wire SB_T3_WEST_SB_OUT_B1_enable;
	input SB_T3_WEST_SB_OUT_B1_ready_in;
	output wire SB_T3_WEST_SB_OUT_B1_valid_out;
	input [0:0] SB_T4_EAST_SB_IN_B1;
	output wire SB_T4_EAST_SB_IN_B1_enable;
	output wire SB_T4_EAST_SB_IN_B1_ready_out;
	input SB_T4_EAST_SB_IN_B1_valid_in;
	output wire [0:0] SB_T4_EAST_SB_OUT_B1;
	output wire SB_T4_EAST_SB_OUT_B1_enable;
	input SB_T4_EAST_SB_OUT_B1_ready_in;
	output wire SB_T4_EAST_SB_OUT_B1_valid_out;
	input [0:0] SB_T4_NORTH_SB_IN_B1;
	output wire SB_T4_NORTH_SB_IN_B1_enable;
	output wire SB_T4_NORTH_SB_IN_B1_ready_out;
	input SB_T4_NORTH_SB_IN_B1_valid_in;
	output wire [0:0] SB_T4_NORTH_SB_OUT_B1;
	output wire SB_T4_NORTH_SB_OUT_B1_enable;
	input SB_T4_NORTH_SB_OUT_B1_ready_in;
	output wire SB_T4_NORTH_SB_OUT_B1_valid_out;
	input [0:0] SB_T4_SOUTH_SB_IN_B1;
	output wire SB_T4_SOUTH_SB_IN_B1_enable;
	output wire SB_T4_SOUTH_SB_IN_B1_ready_out;
	input SB_T4_SOUTH_SB_IN_B1_valid_in;
	output wire [0:0] SB_T4_SOUTH_SB_OUT_B1;
	output wire SB_T4_SOUTH_SB_OUT_B1_enable;
	input SB_T4_SOUTH_SB_OUT_B1_ready_in;
	output wire SB_T4_SOUTH_SB_OUT_B1_valid_out;
	input [0:0] SB_T4_WEST_SB_IN_B1;
	output wire SB_T4_WEST_SB_IN_B1_enable;
	output wire SB_T4_WEST_SB_IN_B1_ready_out;
	input SB_T4_WEST_SB_IN_B1_valid_in;
	output wire [0:0] SB_T4_WEST_SB_OUT_B1;
	output wire SB_T4_WEST_SB_OUT_B1_enable;
	input SB_T4_WEST_SB_OUT_B1_ready_in;
	output wire SB_T4_WEST_SB_OUT_B1_valid_out;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output wire [31:0] read_config_data;
	input reset;
	input [0:0] stall;
	wire [0:0] CB_PE_output_width_1_num_0_fan_in_O;
	wire [0:0] CB_PondTop_output_width_1_num_0_fan_in_O;
	wire [0:0] CB_PondTop_output_width_1_num_1_fan_in_O;
	wire [0:0] Invert1_inst0_out;
	wire [0:0] MUX_SB_T0_EAST_SB_OUT_B1_O;
	wire MUX_SB_T0_EAST_SB_OUT_B1_ready_out;
	wire MUX_SB_T0_EAST_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T0_EAST_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T0_NORTH_SB_OUT_B1_O;
	wire MUX_SB_T0_NORTH_SB_OUT_B1_ready_out;
	wire MUX_SB_T0_NORTH_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T0_NORTH_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T0_SOUTH_SB_OUT_B1_O;
	wire MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out;
	wire MUX_SB_T0_SOUTH_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T0_WEST_SB_OUT_B1_O;
	wire MUX_SB_T0_WEST_SB_OUT_B1_ready_out;
	wire MUX_SB_T0_WEST_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T0_WEST_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T1_EAST_SB_OUT_B1_O;
	wire MUX_SB_T1_EAST_SB_OUT_B1_ready_out;
	wire MUX_SB_T1_EAST_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T1_EAST_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T1_NORTH_SB_OUT_B1_O;
	wire MUX_SB_T1_NORTH_SB_OUT_B1_ready_out;
	wire MUX_SB_T1_NORTH_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T1_NORTH_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T1_SOUTH_SB_OUT_B1_O;
	wire MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out;
	wire MUX_SB_T1_SOUTH_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T1_WEST_SB_OUT_B1_O;
	wire MUX_SB_T1_WEST_SB_OUT_B1_ready_out;
	wire MUX_SB_T1_WEST_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T1_WEST_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T2_EAST_SB_OUT_B1_O;
	wire MUX_SB_T2_EAST_SB_OUT_B1_ready_out;
	wire MUX_SB_T2_EAST_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T2_EAST_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T2_NORTH_SB_OUT_B1_O;
	wire MUX_SB_T2_NORTH_SB_OUT_B1_ready_out;
	wire MUX_SB_T2_NORTH_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T2_NORTH_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T2_SOUTH_SB_OUT_B1_O;
	wire MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out;
	wire MUX_SB_T2_SOUTH_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T2_WEST_SB_OUT_B1_O;
	wire MUX_SB_T2_WEST_SB_OUT_B1_ready_out;
	wire MUX_SB_T2_WEST_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T2_WEST_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T3_EAST_SB_OUT_B1_O;
	wire MUX_SB_T3_EAST_SB_OUT_B1_ready_out;
	wire MUX_SB_T3_EAST_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T3_EAST_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T3_NORTH_SB_OUT_B1_O;
	wire MUX_SB_T3_NORTH_SB_OUT_B1_ready_out;
	wire MUX_SB_T3_NORTH_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T3_NORTH_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T3_SOUTH_SB_OUT_B1_O;
	wire MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out;
	wire MUX_SB_T3_SOUTH_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T3_WEST_SB_OUT_B1_O;
	wire MUX_SB_T3_WEST_SB_OUT_B1_ready_out;
	wire MUX_SB_T3_WEST_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T3_WEST_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T4_EAST_SB_OUT_B1_O;
	wire MUX_SB_T4_EAST_SB_OUT_B1_ready_out;
	wire MUX_SB_T4_EAST_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T4_EAST_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T4_NORTH_SB_OUT_B1_O;
	wire MUX_SB_T4_NORTH_SB_OUT_B1_ready_out;
	wire MUX_SB_T4_NORTH_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T4_NORTH_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T4_SOUTH_SB_OUT_B1_O;
	wire MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out;
	wire MUX_SB_T4_SOUTH_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T4_WEST_SB_OUT_B1_O;
	wire MUX_SB_T4_WEST_SB_OUT_B1_ready_out;
	wire MUX_SB_T4_WEST_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T4_WEST_SB_OUT_B1_out_sel;
	wire [0:0] REG_T0_EAST_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T0_EAST_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T0_EAST_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T0_EAST_B1_end_value_O;
	wire [0:0] REG_T0_EAST_B1_fifo_value_O;
	wire [0:0] REG_T0_EAST_B1_start_value_O;
	wire [0:0] REG_T0_NORTH_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T0_NORTH_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T0_NORTH_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T0_NORTH_B1_end_value_O;
	wire [0:0] REG_T0_NORTH_B1_fifo_value_O;
	wire [0:0] REG_T0_NORTH_B1_start_value_O;
	wire [0:0] REG_T0_SOUTH_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T0_SOUTH_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T0_SOUTH_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T0_SOUTH_B1_end_value_O;
	wire [0:0] REG_T0_SOUTH_B1_fifo_value_O;
	wire [0:0] REG_T0_SOUTH_B1_start_value_O;
	wire [0:0] REG_T0_WEST_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T0_WEST_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T0_WEST_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T0_WEST_B1_end_value_O;
	wire [0:0] REG_T0_WEST_B1_fifo_value_O;
	wire [0:0] REG_T0_WEST_B1_start_value_O;
	wire [0:0] REG_T1_EAST_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T1_EAST_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T1_EAST_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T1_EAST_B1_end_value_O;
	wire [0:0] REG_T1_EAST_B1_fifo_value_O;
	wire [0:0] REG_T1_EAST_B1_start_value_O;
	wire [0:0] REG_T1_NORTH_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T1_NORTH_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T1_NORTH_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T1_NORTH_B1_end_value_O;
	wire [0:0] REG_T1_NORTH_B1_fifo_value_O;
	wire [0:0] REG_T1_NORTH_B1_start_value_O;
	wire [0:0] REG_T1_SOUTH_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T1_SOUTH_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T1_SOUTH_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T1_SOUTH_B1_end_value_O;
	wire [0:0] REG_T1_SOUTH_B1_fifo_value_O;
	wire [0:0] REG_T1_SOUTH_B1_start_value_O;
	wire [0:0] REG_T1_WEST_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T1_WEST_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T1_WEST_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T1_WEST_B1_end_value_O;
	wire [0:0] REG_T1_WEST_B1_fifo_value_O;
	wire [0:0] REG_T1_WEST_B1_start_value_O;
	wire [0:0] REG_T2_EAST_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T2_EAST_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T2_EAST_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T2_EAST_B1_end_value_O;
	wire [0:0] REG_T2_EAST_B1_fifo_value_O;
	wire [0:0] REG_T2_EAST_B1_start_value_O;
	wire [0:0] REG_T2_NORTH_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T2_NORTH_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T2_NORTH_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T2_NORTH_B1_end_value_O;
	wire [0:0] REG_T2_NORTH_B1_fifo_value_O;
	wire [0:0] REG_T2_NORTH_B1_start_value_O;
	wire [0:0] REG_T2_SOUTH_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T2_SOUTH_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T2_SOUTH_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T2_SOUTH_B1_end_value_O;
	wire [0:0] REG_T2_SOUTH_B1_fifo_value_O;
	wire [0:0] REG_T2_SOUTH_B1_start_value_O;
	wire [0:0] REG_T2_WEST_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T2_WEST_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T2_WEST_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T2_WEST_B1_end_value_O;
	wire [0:0] REG_T2_WEST_B1_fifo_value_O;
	wire [0:0] REG_T2_WEST_B1_start_value_O;
	wire [0:0] REG_T3_EAST_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T3_EAST_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T3_EAST_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T3_EAST_B1_end_value_O;
	wire [0:0] REG_T3_EAST_B1_fifo_value_O;
	wire [0:0] REG_T3_EAST_B1_start_value_O;
	wire [0:0] REG_T3_NORTH_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T3_NORTH_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T3_NORTH_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T3_NORTH_B1_end_value_O;
	wire [0:0] REG_T3_NORTH_B1_fifo_value_O;
	wire [0:0] REG_T3_NORTH_B1_start_value_O;
	wire [0:0] REG_T3_SOUTH_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T3_SOUTH_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T3_SOUTH_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T3_SOUTH_B1_end_value_O;
	wire [0:0] REG_T3_SOUTH_B1_fifo_value_O;
	wire [0:0] REG_T3_SOUTH_B1_start_value_O;
	wire [0:0] REG_T3_WEST_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T3_WEST_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T3_WEST_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T3_WEST_B1_end_value_O;
	wire [0:0] REG_T3_WEST_B1_fifo_value_O;
	wire [0:0] REG_T3_WEST_B1_start_value_O;
	wire [0:0] REG_T4_EAST_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T4_EAST_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T4_EAST_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T4_EAST_B1_end_value_O;
	wire [0:0] REG_T4_EAST_B1_fifo_value_O;
	wire [0:0] REG_T4_EAST_B1_start_value_O;
	wire [0:0] REG_T4_NORTH_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T4_NORTH_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T4_NORTH_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T4_NORTH_B1_end_value_O;
	wire [0:0] REG_T4_NORTH_B1_fifo_value_O;
	wire [0:0] REG_T4_NORTH_B1_start_value_O;
	wire [0:0] REG_T4_SOUTH_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T4_SOUTH_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T4_SOUTH_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T4_SOUTH_B1_end_value_O;
	wire [0:0] REG_T4_SOUTH_B1_fifo_value_O;
	wire [0:0] REG_T4_SOUTH_B1_start_value_O;
	wire [0:0] REG_T4_WEST_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T4_WEST_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T4_WEST_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T4_WEST_B1_end_value_O;
	wire [0:0] REG_T4_WEST_B1_fifo_value_O;
	wire [0:0] REG_T4_WEST_B1_start_value_O;
	wire [0:0] RMUX_T0_EAST_B1_O;
	wire RMUX_T0_EAST_B1_ready_out;
	wire RMUX_T0_EAST_B1_valid_out;
	wire [1:0] RMUX_T0_EAST_B1_out_sel;
	wire [0:0] RMUX_T0_EAST_B1_sel_value_O;
	wire [0:0] RMUX_T0_NORTH_B1_O;
	wire RMUX_T0_NORTH_B1_ready_out;
	wire RMUX_T0_NORTH_B1_valid_out;
	wire [1:0] RMUX_T0_NORTH_B1_out_sel;
	wire [0:0] RMUX_T0_NORTH_B1_sel_value_O;
	wire [0:0] RMUX_T0_SOUTH_B1_O;
	wire RMUX_T0_SOUTH_B1_ready_out;
	wire RMUX_T0_SOUTH_B1_valid_out;
	wire [1:0] RMUX_T0_SOUTH_B1_out_sel;
	wire [0:0] RMUX_T0_SOUTH_B1_sel_value_O;
	wire [0:0] RMUX_T0_WEST_B1_O;
	wire RMUX_T0_WEST_B1_ready_out;
	wire RMUX_T0_WEST_B1_valid_out;
	wire [1:0] RMUX_T0_WEST_B1_out_sel;
	wire [0:0] RMUX_T0_WEST_B1_sel_value_O;
	wire [0:0] RMUX_T1_EAST_B1_O;
	wire RMUX_T1_EAST_B1_ready_out;
	wire RMUX_T1_EAST_B1_valid_out;
	wire [1:0] RMUX_T1_EAST_B1_out_sel;
	wire [0:0] RMUX_T1_EAST_B1_sel_value_O;
	wire [0:0] RMUX_T1_NORTH_B1_O;
	wire RMUX_T1_NORTH_B1_ready_out;
	wire RMUX_T1_NORTH_B1_valid_out;
	wire [1:0] RMUX_T1_NORTH_B1_out_sel;
	wire [0:0] RMUX_T1_NORTH_B1_sel_value_O;
	wire [0:0] RMUX_T1_SOUTH_B1_O;
	wire RMUX_T1_SOUTH_B1_ready_out;
	wire RMUX_T1_SOUTH_B1_valid_out;
	wire [1:0] RMUX_T1_SOUTH_B1_out_sel;
	wire [0:0] RMUX_T1_SOUTH_B1_sel_value_O;
	wire [0:0] RMUX_T1_WEST_B1_O;
	wire RMUX_T1_WEST_B1_ready_out;
	wire RMUX_T1_WEST_B1_valid_out;
	wire [1:0] RMUX_T1_WEST_B1_out_sel;
	wire [0:0] RMUX_T1_WEST_B1_sel_value_O;
	wire [0:0] RMUX_T2_EAST_B1_O;
	wire RMUX_T2_EAST_B1_ready_out;
	wire RMUX_T2_EAST_B1_valid_out;
	wire [1:0] RMUX_T2_EAST_B1_out_sel;
	wire [0:0] RMUX_T2_EAST_B1_sel_value_O;
	wire [0:0] RMUX_T2_NORTH_B1_O;
	wire RMUX_T2_NORTH_B1_ready_out;
	wire RMUX_T2_NORTH_B1_valid_out;
	wire [1:0] RMUX_T2_NORTH_B1_out_sel;
	wire [0:0] RMUX_T2_NORTH_B1_sel_value_O;
	wire [0:0] RMUX_T2_SOUTH_B1_O;
	wire RMUX_T2_SOUTH_B1_ready_out;
	wire RMUX_T2_SOUTH_B1_valid_out;
	wire [1:0] RMUX_T2_SOUTH_B1_out_sel;
	wire [0:0] RMUX_T2_SOUTH_B1_sel_value_O;
	wire [0:0] RMUX_T2_WEST_B1_O;
	wire RMUX_T2_WEST_B1_ready_out;
	wire RMUX_T2_WEST_B1_valid_out;
	wire [1:0] RMUX_T2_WEST_B1_out_sel;
	wire [0:0] RMUX_T2_WEST_B1_sel_value_O;
	wire [0:0] RMUX_T3_EAST_B1_O;
	wire RMUX_T3_EAST_B1_ready_out;
	wire RMUX_T3_EAST_B1_valid_out;
	wire [1:0] RMUX_T3_EAST_B1_out_sel;
	wire [0:0] RMUX_T3_EAST_B1_sel_value_O;
	wire [0:0] RMUX_T3_NORTH_B1_O;
	wire RMUX_T3_NORTH_B1_ready_out;
	wire RMUX_T3_NORTH_B1_valid_out;
	wire [1:0] RMUX_T3_NORTH_B1_out_sel;
	wire [0:0] RMUX_T3_NORTH_B1_sel_value_O;
	wire [0:0] RMUX_T3_SOUTH_B1_O;
	wire RMUX_T3_SOUTH_B1_ready_out;
	wire RMUX_T3_SOUTH_B1_valid_out;
	wire [1:0] RMUX_T3_SOUTH_B1_out_sel;
	wire [0:0] RMUX_T3_SOUTH_B1_sel_value_O;
	wire [0:0] RMUX_T3_WEST_B1_O;
	wire RMUX_T3_WEST_B1_ready_out;
	wire RMUX_T3_WEST_B1_valid_out;
	wire [1:0] RMUX_T3_WEST_B1_out_sel;
	wire [0:0] RMUX_T3_WEST_B1_sel_value_O;
	wire [0:0] RMUX_T4_EAST_B1_O;
	wire RMUX_T4_EAST_B1_ready_out;
	wire RMUX_T4_EAST_B1_valid_out;
	wire [1:0] RMUX_T4_EAST_B1_out_sel;
	wire [0:0] RMUX_T4_EAST_B1_sel_value_O;
	wire [0:0] RMUX_T4_NORTH_B1_O;
	wire RMUX_T4_NORTH_B1_ready_out;
	wire RMUX_T4_NORTH_B1_valid_out;
	wire [1:0] RMUX_T4_NORTH_B1_out_sel;
	wire [0:0] RMUX_T4_NORTH_B1_sel_value_O;
	wire [0:0] RMUX_T4_SOUTH_B1_O;
	wire RMUX_T4_SOUTH_B1_ready_out;
	wire RMUX_T4_SOUTH_B1_valid_out;
	wire [1:0] RMUX_T4_SOUTH_B1_out_sel;
	wire [0:0] RMUX_T4_SOUTH_B1_sel_value_O;
	wire [0:0] RMUX_T4_WEST_B1_O;
	wire RMUX_T4_WEST_B1_ready_out;
	wire RMUX_T4_WEST_B1_valid_out;
	wire [1:0] RMUX_T4_WEST_B1_out_sel;
	wire [0:0] RMUX_T4_WEST_B1_sel_value_O;
	wire [0:0] SB_T0_EAST_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T0_EAST_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T0_EAST_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T0_EAST_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T0_EAST_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T0_NORTH_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T0_NORTH_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T0_NORTH_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T0_NORTH_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T0_NORTH_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T0_SOUTH_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T0_SOUTH_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T0_SOUTH_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T0_SOUTH_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T0_SOUTH_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T0_WEST_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T0_WEST_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T0_WEST_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T0_WEST_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T0_WEST_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T1_EAST_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T1_EAST_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T1_EAST_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T1_EAST_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T1_EAST_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T1_NORTH_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T1_NORTH_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T1_NORTH_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T1_NORTH_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T1_NORTH_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T1_SOUTH_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T1_SOUTH_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T1_SOUTH_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T1_SOUTH_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T1_SOUTH_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T1_WEST_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T1_WEST_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T1_WEST_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T1_WEST_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T1_WEST_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T2_EAST_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T2_EAST_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T2_EAST_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T2_EAST_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T2_EAST_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T2_NORTH_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T2_NORTH_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T2_NORTH_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T2_NORTH_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T2_NORTH_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T2_SOUTH_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T2_SOUTH_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T2_SOUTH_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T2_SOUTH_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T2_SOUTH_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T2_WEST_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T2_WEST_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T2_WEST_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T2_WEST_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T2_WEST_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T3_EAST_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T3_EAST_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T3_EAST_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T3_EAST_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T3_EAST_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T3_NORTH_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T3_NORTH_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T3_NORTH_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T3_NORTH_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T3_NORTH_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T3_SOUTH_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T3_SOUTH_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T3_SOUTH_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T3_SOUTH_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T3_SOUTH_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T3_WEST_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T3_WEST_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T3_WEST_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T3_WEST_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T3_WEST_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T4_EAST_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T4_EAST_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T4_EAST_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T4_EAST_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T4_EAST_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T4_NORTH_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T4_NORTH_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T4_NORTH_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T4_NORTH_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T4_NORTH_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T4_SOUTH_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T4_SOUTH_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T4_SOUTH_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T4_SOUTH_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T4_SOUTH_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T4_WEST_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T4_WEST_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T4_WEST_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T4_WEST_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T4_WEST_SB_OUT_B1_sel_value_O;
	wire [0:0] WIRE_SB_T0_EAST_SB_IN_B1_O;
	wire WIRE_SB_T0_EAST_SB_IN_B1_ready_out;
	wire WIRE_SB_T0_EAST_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T0_NORTH_SB_IN_B1_O;
	wire WIRE_SB_T0_NORTH_SB_IN_B1_ready_out;
	wire WIRE_SB_T0_NORTH_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T0_SOUTH_SB_IN_B1_O;
	wire WIRE_SB_T0_SOUTH_SB_IN_B1_ready_out;
	wire WIRE_SB_T0_SOUTH_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T0_WEST_SB_IN_B1_O;
	wire WIRE_SB_T0_WEST_SB_IN_B1_ready_out;
	wire WIRE_SB_T0_WEST_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T1_EAST_SB_IN_B1_O;
	wire WIRE_SB_T1_EAST_SB_IN_B1_ready_out;
	wire WIRE_SB_T1_EAST_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T1_NORTH_SB_IN_B1_O;
	wire WIRE_SB_T1_NORTH_SB_IN_B1_ready_out;
	wire WIRE_SB_T1_NORTH_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T1_SOUTH_SB_IN_B1_O;
	wire WIRE_SB_T1_SOUTH_SB_IN_B1_ready_out;
	wire WIRE_SB_T1_SOUTH_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T1_WEST_SB_IN_B1_O;
	wire WIRE_SB_T1_WEST_SB_IN_B1_ready_out;
	wire WIRE_SB_T1_WEST_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T2_EAST_SB_IN_B1_O;
	wire WIRE_SB_T2_EAST_SB_IN_B1_ready_out;
	wire WIRE_SB_T2_EAST_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T2_NORTH_SB_IN_B1_O;
	wire WIRE_SB_T2_NORTH_SB_IN_B1_ready_out;
	wire WIRE_SB_T2_NORTH_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T2_SOUTH_SB_IN_B1_O;
	wire WIRE_SB_T2_SOUTH_SB_IN_B1_ready_out;
	wire WIRE_SB_T2_SOUTH_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T2_WEST_SB_IN_B1_O;
	wire WIRE_SB_T2_WEST_SB_IN_B1_ready_out;
	wire WIRE_SB_T2_WEST_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T3_EAST_SB_IN_B1_O;
	wire WIRE_SB_T3_EAST_SB_IN_B1_ready_out;
	wire WIRE_SB_T3_EAST_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T3_NORTH_SB_IN_B1_O;
	wire WIRE_SB_T3_NORTH_SB_IN_B1_ready_out;
	wire WIRE_SB_T3_NORTH_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T3_SOUTH_SB_IN_B1_O;
	wire WIRE_SB_T3_SOUTH_SB_IN_B1_ready_out;
	wire WIRE_SB_T3_SOUTH_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T3_WEST_SB_IN_B1_O;
	wire WIRE_SB_T3_WEST_SB_IN_B1_ready_out;
	wire WIRE_SB_T3_WEST_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T4_EAST_SB_IN_B1_O;
	wire WIRE_SB_T4_EAST_SB_IN_B1_ready_out;
	wire WIRE_SB_T4_EAST_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T4_NORTH_SB_IN_B1_O;
	wire WIRE_SB_T4_NORTH_SB_IN_B1_ready_out;
	wire WIRE_SB_T4_NORTH_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T4_SOUTH_SB_IN_B1_O;
	wire WIRE_SB_T4_SOUTH_SB_IN_B1_ready_out;
	wire WIRE_SB_T4_SOUTH_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T4_WEST_SB_IN_B1_O;
	wire WIRE_SB_T4_WEST_SB_IN_B1_ready_out;
	wire WIRE_SB_T4_WEST_SB_IN_B1_valid_out;
	wire ZextWrapper_23_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_23_32_inst0$self_O_in;
	wire ZextWrapper_30_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_30_32_inst0$self_O_in;
	wire ZextWrapper_31_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_31_32_inst0$self_O_in;
	wire [0:0] and1_inst0_out;
	wire [0:0] and1_inst1_out;
	wire [0:0] and1_inst10_out;
	wire [0:0] and1_inst11_out;
	wire [0:0] and1_inst12_out;
	wire [0:0] and1_inst13_out;
	wire [0:0] and1_inst14_out;
	wire [0:0] and1_inst15_out;
	wire [0:0] and1_inst16_out;
	wire [0:0] and1_inst17_out;
	wire [0:0] and1_inst18_out;
	wire [0:0] and1_inst19_out;
	wire [0:0] and1_inst2_out;
	wire [0:0] and1_inst3_out;
	wire [0:0] and1_inst4_out;
	wire [0:0] and1_inst5_out;
	wire [0:0] and1_inst6_out;
	wire [0:0] and1_inst7_out;
	wire [0:0] and1_inst8_out;
	wire [0:0] and1_inst9_out;
	wire [31:0] config_reg_0_O;
	wire [31:0] config_reg_1_O;
	wire [31:0] config_reg_2_O;
	wire [30:0] config_reg_3_O;
	wire [29:0] config_reg_4_O;
	wire [22:0] config_reg_5_O;
	wire [0:0] const_0_1_out;
	wire [31:0] const_0_32_out;
	wire [0:0] const_1_1_out;
	wire coreir_eq_1_inst0_out;
	wire coreir_eq_1_inst1_out;
	wire coreir_eq_1_inst10_out;
	wire coreir_eq_1_inst11_out;
	wire coreir_eq_1_inst12_out;
	wire coreir_eq_1_inst13_out;
	wire coreir_eq_1_inst14_out;
	wire coreir_eq_1_inst15_out;
	wire coreir_eq_1_inst16_out;
	wire coreir_eq_1_inst17_out;
	wire coreir_eq_1_inst18_out;
	wire coreir_eq_1_inst19_out;
	wire coreir_eq_1_inst2_out;
	wire coreir_eq_1_inst3_out;
	wire coreir_eq_1_inst4_out;
	wire coreir_eq_1_inst5_out;
	wire coreir_eq_1_inst6_out;
	wire coreir_eq_1_inst7_out;
	wire coreir_eq_1_inst8_out;
	wire coreir_eq_1_inst9_out;
	wire [31:0] mux_aoi_6_32_inst0_O;
	wire [7:0] mux_aoi_6_32_inst0_out_sel;
	wire [7:0] self_config_config_addr_out;
	FanoutHash_E70AF988E4250F5 CB_PE_output_width_1_num_0_fan_in(
		.I13(MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out),
		.E8(SB_T2_NORTH_SB_OUT_B1_enable_value_O),
		.E17(SB_T4_SOUTH_SB_OUT_B1_enable_value_O),
		.I15(MUX_SB_T3_WEST_SB_OUT_B1_ready_out),
		.I12(MUX_SB_T3_NORTH_SB_OUT_B1_ready_out),
		.E6(SB_T1_EAST_SB_OUT_B1_enable_value_O),
		.I9(MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out),
		.I16(MUX_SB_T4_NORTH_SB_OUT_B1_ready_out),
		.E3(SB_T0_WEST_SB_OUT_B1_enable_value_O),
		.S14(MUX_SB_T3_EAST_SB_OUT_B1_out_sel),
		.E10(SB_T2_EAST_SB_OUT_B1_enable_value_O),
		.I5(MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out),
		.S6(MUX_SB_T1_EAST_SB_OUT_B1_out_sel),
		.E0(SB_T0_NORTH_SB_OUT_B1_enable_value_O),
		.E18(SB_T4_EAST_SB_OUT_B1_enable_value_O),
		.I19(MUX_SB_T4_WEST_SB_OUT_B1_ready_out),
		.I10(MUX_SB_T2_EAST_SB_OUT_B1_ready_out),
		.S5(MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel),
		.I6(MUX_SB_T1_EAST_SB_OUT_B1_ready_out),
		.I8(MUX_SB_T2_NORTH_SB_OUT_B1_ready_out),
		.S3(MUX_SB_T0_WEST_SB_OUT_B1_out_sel),
		.S10(MUX_SB_T2_EAST_SB_OUT_B1_out_sel),
		.E16(SB_T4_NORTH_SB_OUT_B1_enable_value_O),
		.S4(MUX_SB_T1_NORTH_SB_OUT_B1_out_sel),
		.E11(SB_T2_WEST_SB_OUT_B1_enable_value_O),
		.S19(MUX_SB_T4_WEST_SB_OUT_B1_out_sel),
		.E15(SB_T3_WEST_SB_OUT_B1_enable_value_O),
		.E19(SB_T4_WEST_SB_OUT_B1_enable_value_O),
		.I3(MUX_SB_T0_WEST_SB_OUT_B1_ready_out),
		.I4(MUX_SB_T1_NORTH_SB_OUT_B1_ready_out),
		.S1(MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel),
		.E13(SB_T3_SOUTH_SB_OUT_B1_enable_value_O),
		.S0(MUX_SB_T0_NORTH_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T0_EAST_SB_OUT_B1_out_sel),
		.I11(MUX_SB_T2_WEST_SB_OUT_B1_ready_out),
		.S8(MUX_SB_T2_NORTH_SB_OUT_B1_out_sel),
		.E2(SB_T0_EAST_SB_OUT_B1_enable_value_O),
		.E14(SB_T3_EAST_SB_OUT_B1_enable_value_O),
		.S17(MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel),
		.E5(SB_T1_SOUTH_SB_OUT_B1_enable_value_O),
		.E4(SB_T1_NORTH_SB_OUT_B1_enable_value_O),
		.I1(MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out),
		.I2(MUX_SB_T0_EAST_SB_OUT_B1_ready_out),
		.I17(MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out),
		.O(CB_PE_output_width_1_num_0_fan_in_O),
		.E9(SB_T2_SOUTH_SB_OUT_B1_enable_value_O),
		.S13(MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel),
		.S11(MUX_SB_T2_WEST_SB_OUT_B1_out_sel),
		.S7(MUX_SB_T1_WEST_SB_OUT_B1_out_sel),
		.E1(SB_T0_SOUTH_SB_OUT_B1_enable_value_O),
		.S15(MUX_SB_T3_WEST_SB_OUT_B1_out_sel),
		.S9(MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel),
		.S18(MUX_SB_T4_EAST_SB_OUT_B1_out_sel),
		.S12(MUX_SB_T3_NORTH_SB_OUT_B1_out_sel),
		.I14(MUX_SB_T3_EAST_SB_OUT_B1_ready_out),
		.I7(MUX_SB_T1_WEST_SB_OUT_B1_ready_out),
		.S16(MUX_SB_T4_NORTH_SB_OUT_B1_out_sel),
		.E12(SB_T3_NORTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T0_NORTH_SB_OUT_B1_ready_out),
		.E7(SB_T1_WEST_SB_OUT_B1_enable_value_O),
		.I18(MUX_SB_T4_EAST_SB_OUT_B1_ready_out)
	);
	FanoutHash_F689C91787363AB CB_PondTop_output_width_1_num_0_fan_in(
		.I13(MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out),
		.E8(SB_T2_NORTH_SB_OUT_B1_enable_value_O),
		.E17(SB_T4_SOUTH_SB_OUT_B1_enable_value_O),
		.I15(MUX_SB_T3_WEST_SB_OUT_B1_ready_out),
		.I12(MUX_SB_T3_NORTH_SB_OUT_B1_ready_out),
		.E6(SB_T1_EAST_SB_OUT_B1_enable_value_O),
		.I9(MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out),
		.I16(MUX_SB_T4_NORTH_SB_OUT_B1_ready_out),
		.E3(SB_T0_WEST_SB_OUT_B1_enable_value_O),
		.S14(MUX_SB_T3_EAST_SB_OUT_B1_out_sel),
		.E10(SB_T2_EAST_SB_OUT_B1_enable_value_O),
		.I20(PE_input_width_1_num_0_ready),
		.I5(MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out),
		.S6(MUX_SB_T1_EAST_SB_OUT_B1_out_sel),
		.E0(SB_T0_NORTH_SB_OUT_B1_enable_value_O),
		.E18(SB_T4_EAST_SB_OUT_B1_enable_value_O),
		.I19(MUX_SB_T4_WEST_SB_OUT_B1_ready_out),
		.I10(MUX_SB_T2_EAST_SB_OUT_B1_ready_out),
		.S5(MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel),
		.I6(MUX_SB_T1_EAST_SB_OUT_B1_ready_out),
		.I8(MUX_SB_T2_NORTH_SB_OUT_B1_ready_out),
		.S3(MUX_SB_T0_WEST_SB_OUT_B1_out_sel),
		.S10(MUX_SB_T2_EAST_SB_OUT_B1_out_sel),
		.E16(SB_T4_NORTH_SB_OUT_B1_enable_value_O),
		.S4(MUX_SB_T1_NORTH_SB_OUT_B1_out_sel),
		.E11(SB_T2_WEST_SB_OUT_B1_enable_value_O),
		.S19(MUX_SB_T4_WEST_SB_OUT_B1_out_sel),
		.E15(SB_T3_WEST_SB_OUT_B1_enable_value_O),
		.E19(SB_T4_WEST_SB_OUT_B1_enable_value_O),
		.I3(MUX_SB_T0_WEST_SB_OUT_B1_ready_out),
		.I4(MUX_SB_T1_NORTH_SB_OUT_B1_ready_out),
		.S1(MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel),
		.E13(SB_T3_SOUTH_SB_OUT_B1_enable_value_O),
		.S0(MUX_SB_T0_NORTH_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T0_EAST_SB_OUT_B1_out_sel),
		.I11(MUX_SB_T2_WEST_SB_OUT_B1_ready_out),
		.S8(MUX_SB_T2_NORTH_SB_OUT_B1_out_sel),
		.E2(SB_T0_EAST_SB_OUT_B1_enable_value_O),
		.E14(SB_T3_EAST_SB_OUT_B1_enable_value_O),
		.S17(MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel),
		.E5(SB_T1_SOUTH_SB_OUT_B1_enable_value_O),
		.E4(SB_T1_NORTH_SB_OUT_B1_enable_value_O),
		.I1(MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out),
		.I2(MUX_SB_T0_EAST_SB_OUT_B1_ready_out),
		.I17(MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out),
		.O(CB_PondTop_output_width_1_num_0_fan_in_O),
		.E9(SB_T2_SOUTH_SB_OUT_B1_enable_value_O),
		.S13(MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel),
		.S11(MUX_SB_T2_WEST_SB_OUT_B1_out_sel),
		.S20(PE_input_width_1_num_0_out_sel),
		.S7(MUX_SB_T1_WEST_SB_OUT_B1_out_sel),
		.E1(SB_T0_SOUTH_SB_OUT_B1_enable_value_O),
		.E20(PE_input_width_1_num_0_enable),
		.S15(MUX_SB_T3_WEST_SB_OUT_B1_out_sel),
		.S9(MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel),
		.S18(MUX_SB_T4_EAST_SB_OUT_B1_out_sel),
		.S12(MUX_SB_T3_NORTH_SB_OUT_B1_out_sel),
		.I14(MUX_SB_T3_EAST_SB_OUT_B1_ready_out),
		.I7(MUX_SB_T1_WEST_SB_OUT_B1_ready_out),
		.S16(MUX_SB_T4_NORTH_SB_OUT_B1_out_sel),
		.E12(SB_T3_NORTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T0_NORTH_SB_OUT_B1_ready_out),
		.E7(SB_T1_WEST_SB_OUT_B1_enable_value_O),
		.I18(MUX_SB_T4_EAST_SB_OUT_B1_ready_out)
	);
	FanoutHash_CE1AA874B742213 CB_PondTop_output_width_1_num_1_fan_in(
		.I13(MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out),
		.E8(SB_T2_NORTH_SB_OUT_B1_enable_value_O),
		.E17(SB_T4_SOUTH_SB_OUT_B1_enable_value_O),
		.I15(MUX_SB_T3_WEST_SB_OUT_B1_ready_out),
		.I12(MUX_SB_T3_NORTH_SB_OUT_B1_ready_out),
		.E6(SB_T1_EAST_SB_OUT_B1_enable_value_O),
		.I9(MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out),
		.I16(MUX_SB_T4_NORTH_SB_OUT_B1_ready_out),
		.E3(SB_T0_WEST_SB_OUT_B1_enable_value_O),
		.S14(MUX_SB_T3_EAST_SB_OUT_B1_out_sel),
		.E10(SB_T2_EAST_SB_OUT_B1_enable_value_O),
		.I5(MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out),
		.S6(MUX_SB_T1_EAST_SB_OUT_B1_out_sel),
		.E0(SB_T0_NORTH_SB_OUT_B1_enable_value_O),
		.E18(SB_T4_EAST_SB_OUT_B1_enable_value_O),
		.I19(MUX_SB_T4_WEST_SB_OUT_B1_ready_out),
		.I10(MUX_SB_T2_EAST_SB_OUT_B1_ready_out),
		.S5(MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel),
		.I6(MUX_SB_T1_EAST_SB_OUT_B1_ready_out),
		.I8(MUX_SB_T2_NORTH_SB_OUT_B1_ready_out),
		.S3(MUX_SB_T0_WEST_SB_OUT_B1_out_sel),
		.S10(MUX_SB_T2_EAST_SB_OUT_B1_out_sel),
		.E16(SB_T4_NORTH_SB_OUT_B1_enable_value_O),
		.S4(MUX_SB_T1_NORTH_SB_OUT_B1_out_sel),
		.E11(SB_T2_WEST_SB_OUT_B1_enable_value_O),
		.S19(MUX_SB_T4_WEST_SB_OUT_B1_out_sel),
		.E15(SB_T3_WEST_SB_OUT_B1_enable_value_O),
		.E19(SB_T4_WEST_SB_OUT_B1_enable_value_O),
		.I3(MUX_SB_T0_WEST_SB_OUT_B1_ready_out),
		.I4(MUX_SB_T1_NORTH_SB_OUT_B1_ready_out),
		.S1(MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel),
		.E13(SB_T3_SOUTH_SB_OUT_B1_enable_value_O),
		.S0(MUX_SB_T0_NORTH_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T0_EAST_SB_OUT_B1_out_sel),
		.I11(MUX_SB_T2_WEST_SB_OUT_B1_ready_out),
		.S8(MUX_SB_T2_NORTH_SB_OUT_B1_out_sel),
		.E2(SB_T0_EAST_SB_OUT_B1_enable_value_O),
		.E14(SB_T3_EAST_SB_OUT_B1_enable_value_O),
		.S17(MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel),
		.E5(SB_T1_SOUTH_SB_OUT_B1_enable_value_O),
		.E4(SB_T1_NORTH_SB_OUT_B1_enable_value_O),
		.I1(MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out),
		.I2(MUX_SB_T0_EAST_SB_OUT_B1_ready_out),
		.I17(MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out),
		.O(CB_PondTop_output_width_1_num_1_fan_in_O),
		.E9(SB_T2_SOUTH_SB_OUT_B1_enable_value_O),
		.S13(MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel),
		.S11(MUX_SB_T2_WEST_SB_OUT_B1_out_sel),
		.S7(MUX_SB_T1_WEST_SB_OUT_B1_out_sel),
		.E1(SB_T0_SOUTH_SB_OUT_B1_enable_value_O),
		.S15(MUX_SB_T3_WEST_SB_OUT_B1_out_sel),
		.S9(MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel),
		.S18(MUX_SB_T4_EAST_SB_OUT_B1_out_sel),
		.S12(MUX_SB_T3_NORTH_SB_OUT_B1_out_sel),
		.I14(MUX_SB_T3_EAST_SB_OUT_B1_ready_out),
		.I7(MUX_SB_T1_WEST_SB_OUT_B1_ready_out),
		.S16(MUX_SB_T4_NORTH_SB_OUT_B1_out_sel),
		.E12(SB_T3_NORTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T0_NORTH_SB_OUT_B1_ready_out),
		.E7(SB_T1_WEST_SB_OUT_B1_enable_value_O),
		.I18(MUX_SB_T4_EAST_SB_OUT_B1_ready_out)
	);
	coreir_not #(.width(1)) Invert1_inst0(
		.in(stall),
		.out(Invert1_inst0_out)
	);
	wire [5:0] MUX_SB_T0_EAST_SB_OUT_B1_I;
	assign MUX_SB_T0_EAST_SB_OUT_B1_I[5+:1] = PondTop_output_width_1_num_1;
	assign MUX_SB_T0_EAST_SB_OUT_B1_I[4+:1] = PondTop_output_width_1_num_0;
	assign MUX_SB_T0_EAST_SB_OUT_B1_I[3+:1] = PE_output_width_1_num_0;
	assign MUX_SB_T0_EAST_SB_OUT_B1_I[2+:1] = WIRE_SB_T4_NORTH_SB_IN_B1_O;
	assign MUX_SB_T0_EAST_SB_OUT_B1_I[1+:1] = WIRE_SB_T3_SOUTH_SB_IN_B1_O;
	assign MUX_SB_T0_EAST_SB_OUT_B1_I[0+:1] = WIRE_SB_T0_WEST_SB_IN_B1_O;
	wire [5:0] MUX_SB_T0_EAST_SB_OUT_B1_valid_in;
	assign MUX_SB_T0_EAST_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid, PondTop_output_width_1_num_0_valid, PE_output_width_1_num_0_valid, WIRE_SB_T4_NORTH_SB_IN_B1_valid_out, WIRE_SB_T3_SOUTH_SB_IN_B1_valid_out, WIRE_SB_T0_WEST_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T0_EAST_SB_OUT_B1(
		.I(MUX_SB_T0_EAST_SB_OUT_B1_I),
		.O(MUX_SB_T0_EAST_SB_OUT_B1_O),
		.ready_in(SB_T0_EAST_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T0_EAST_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T0_EAST_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T0_EAST_SB_OUT_B1_valid_out),
		.S(SB_T0_EAST_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T0_EAST_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T0_NORTH_SB_OUT_B1_I;
	assign MUX_SB_T0_NORTH_SB_OUT_B1_I[5+:1] = PondTop_output_width_1_num_1;
	assign MUX_SB_T0_NORTH_SB_OUT_B1_I[4+:1] = PondTop_output_width_1_num_0;
	assign MUX_SB_T0_NORTH_SB_OUT_B1_I[3+:1] = PE_output_width_1_num_0;
	assign MUX_SB_T0_NORTH_SB_OUT_B1_I[2+:1] = WIRE_SB_T0_SOUTH_SB_IN_B1_O;
	assign MUX_SB_T0_NORTH_SB_OUT_B1_I[1+:1] = WIRE_SB_T1_EAST_SB_IN_B1_O;
	assign MUX_SB_T0_NORTH_SB_OUT_B1_I[0+:1] = WIRE_SB_T0_WEST_SB_IN_B1_O;
	wire [5:0] MUX_SB_T0_NORTH_SB_OUT_B1_valid_in;
	assign MUX_SB_T0_NORTH_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid, PondTop_output_width_1_num_0_valid, PE_output_width_1_num_0_valid, WIRE_SB_T0_SOUTH_SB_IN_B1_valid_out, WIRE_SB_T1_EAST_SB_IN_B1_valid_out, WIRE_SB_T0_WEST_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T0_NORTH_SB_OUT_B1(
		.I(MUX_SB_T0_NORTH_SB_OUT_B1_I),
		.O(MUX_SB_T0_NORTH_SB_OUT_B1_O),
		.ready_in(SB_T0_NORTH_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T0_NORTH_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T0_NORTH_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T0_NORTH_SB_OUT_B1_valid_out),
		.S(SB_T0_NORTH_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T0_NORTH_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T0_SOUTH_SB_OUT_B1_I;
	assign MUX_SB_T0_SOUTH_SB_OUT_B1_I[5+:1] = PondTop_output_width_1_num_1;
	assign MUX_SB_T0_SOUTH_SB_OUT_B1_I[4+:1] = PondTop_output_width_1_num_0;
	assign MUX_SB_T0_SOUTH_SB_OUT_B1_I[3+:1] = PE_output_width_1_num_0;
	assign MUX_SB_T0_SOUTH_SB_OUT_B1_I[2+:1] = WIRE_SB_T1_WEST_SB_IN_B1_O;
	assign MUX_SB_T0_SOUTH_SB_OUT_B1_I[1+:1] = WIRE_SB_T0_NORTH_SB_IN_B1_O;
	assign MUX_SB_T0_SOUTH_SB_OUT_B1_I[0+:1] = WIRE_SB_T3_EAST_SB_IN_B1_O;
	wire [5:0] MUX_SB_T0_SOUTH_SB_OUT_B1_valid_in;
	assign MUX_SB_T0_SOUTH_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid, PondTop_output_width_1_num_0_valid, PE_output_width_1_num_0_valid, WIRE_SB_T1_WEST_SB_IN_B1_valid_out, WIRE_SB_T0_NORTH_SB_IN_B1_valid_out, WIRE_SB_T3_EAST_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T0_SOUTH_SB_OUT_B1(
		.I(MUX_SB_T0_SOUTH_SB_OUT_B1_I),
		.O(MUX_SB_T0_SOUTH_SB_OUT_B1_O),
		.ready_in(SB_T0_SOUTH_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T0_SOUTH_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T0_SOUTH_SB_OUT_B1_valid_out),
		.S(SB_T0_SOUTH_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T0_WEST_SB_OUT_B1_I;
	assign MUX_SB_T0_WEST_SB_OUT_B1_I[5+:1] = PondTop_output_width_1_num_1;
	assign MUX_SB_T0_WEST_SB_OUT_B1_I[4+:1] = PondTop_output_width_1_num_0;
	assign MUX_SB_T0_WEST_SB_OUT_B1_I[3+:1] = PE_output_width_1_num_0;
	assign MUX_SB_T0_WEST_SB_OUT_B1_I[2+:1] = WIRE_SB_T0_EAST_SB_IN_B1_O;
	assign MUX_SB_T0_WEST_SB_OUT_B1_I[1+:1] = WIRE_SB_T4_SOUTH_SB_IN_B1_O;
	assign MUX_SB_T0_WEST_SB_OUT_B1_I[0+:1] = WIRE_SB_T0_NORTH_SB_IN_B1_O;
	wire [5:0] MUX_SB_T0_WEST_SB_OUT_B1_valid_in;
	assign MUX_SB_T0_WEST_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid, PondTop_output_width_1_num_0_valid, PE_output_width_1_num_0_valid, WIRE_SB_T0_EAST_SB_IN_B1_valid_out, WIRE_SB_T4_SOUTH_SB_IN_B1_valid_out, WIRE_SB_T0_NORTH_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T0_WEST_SB_OUT_B1(
		.I(MUX_SB_T0_WEST_SB_OUT_B1_I),
		.O(MUX_SB_T0_WEST_SB_OUT_B1_O),
		.ready_in(SB_T0_WEST_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T0_WEST_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T0_WEST_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T0_WEST_SB_OUT_B1_valid_out),
		.S(SB_T0_WEST_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T0_WEST_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T1_EAST_SB_OUT_B1_I;
	assign MUX_SB_T1_EAST_SB_OUT_B1_I[5+:1] = PondTop_output_width_1_num_1;
	assign MUX_SB_T1_EAST_SB_OUT_B1_I[4+:1] = PondTop_output_width_1_num_0;
	assign MUX_SB_T1_EAST_SB_OUT_B1_I[3+:1] = PE_output_width_1_num_0;
	assign MUX_SB_T1_EAST_SB_OUT_B1_I[2+:1] = WIRE_SB_T2_SOUTH_SB_IN_B1_O;
	assign MUX_SB_T1_EAST_SB_OUT_B1_I[1+:1] = WIRE_SB_T1_WEST_SB_IN_B1_O;
	assign MUX_SB_T1_EAST_SB_OUT_B1_I[0+:1] = WIRE_SB_T0_NORTH_SB_IN_B1_O;
	wire [5:0] MUX_SB_T1_EAST_SB_OUT_B1_valid_in;
	assign MUX_SB_T1_EAST_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid, PondTop_output_width_1_num_0_valid, PE_output_width_1_num_0_valid, WIRE_SB_T2_SOUTH_SB_IN_B1_valid_out, WIRE_SB_T1_WEST_SB_IN_B1_valid_out, WIRE_SB_T0_NORTH_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T1_EAST_SB_OUT_B1(
		.I(MUX_SB_T1_EAST_SB_OUT_B1_I),
		.O(MUX_SB_T1_EAST_SB_OUT_B1_O),
		.ready_in(SB_T1_EAST_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T1_EAST_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T1_EAST_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T1_EAST_SB_OUT_B1_valid_out),
		.S(SB_T1_EAST_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T1_EAST_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T1_NORTH_SB_OUT_B1_I;
	assign MUX_SB_T1_NORTH_SB_OUT_B1_I[5+:1] = PondTop_output_width_1_num_1;
	assign MUX_SB_T1_NORTH_SB_OUT_B1_I[4+:1] = PondTop_output_width_1_num_0;
	assign MUX_SB_T1_NORTH_SB_OUT_B1_I[3+:1] = PE_output_width_1_num_0;
	assign MUX_SB_T1_NORTH_SB_OUT_B1_I[2+:1] = WIRE_SB_T4_WEST_SB_IN_B1_O;
	assign MUX_SB_T1_NORTH_SB_OUT_B1_I[1+:1] = WIRE_SB_T1_SOUTH_SB_IN_B1_O;
	assign MUX_SB_T1_NORTH_SB_OUT_B1_I[0+:1] = WIRE_SB_T2_EAST_SB_IN_B1_O;
	wire [5:0] MUX_SB_T1_NORTH_SB_OUT_B1_valid_in;
	assign MUX_SB_T1_NORTH_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid, PondTop_output_width_1_num_0_valid, PE_output_width_1_num_0_valid, WIRE_SB_T4_WEST_SB_IN_B1_valid_out, WIRE_SB_T1_SOUTH_SB_IN_B1_valid_out, WIRE_SB_T2_EAST_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T1_NORTH_SB_OUT_B1(
		.I(MUX_SB_T1_NORTH_SB_OUT_B1_I),
		.O(MUX_SB_T1_NORTH_SB_OUT_B1_O),
		.ready_in(SB_T1_NORTH_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T1_NORTH_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T1_NORTH_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T1_NORTH_SB_OUT_B1_valid_out),
		.S(SB_T1_NORTH_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T1_NORTH_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T1_SOUTH_SB_OUT_B1_I;
	assign MUX_SB_T1_SOUTH_SB_OUT_B1_I[5+:1] = PondTop_output_width_1_num_1;
	assign MUX_SB_T1_SOUTH_SB_OUT_B1_I[4+:1] = PondTop_output_width_1_num_0;
	assign MUX_SB_T1_SOUTH_SB_OUT_B1_I[3+:1] = PE_output_width_1_num_0;
	assign MUX_SB_T1_SOUTH_SB_OUT_B1_I[2+:1] = WIRE_SB_T2_WEST_SB_IN_B1_O;
	assign MUX_SB_T1_SOUTH_SB_OUT_B1_I[1+:1] = WIRE_SB_T1_NORTH_SB_IN_B1_O;
	assign MUX_SB_T1_SOUTH_SB_OUT_B1_I[0+:1] = WIRE_SB_T2_EAST_SB_IN_B1_O;
	wire [5:0] MUX_SB_T1_SOUTH_SB_OUT_B1_valid_in;
	assign MUX_SB_T1_SOUTH_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid, PondTop_output_width_1_num_0_valid, PE_output_width_1_num_0_valid, WIRE_SB_T2_WEST_SB_IN_B1_valid_out, WIRE_SB_T1_NORTH_SB_IN_B1_valid_out, WIRE_SB_T2_EAST_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T1_SOUTH_SB_OUT_B1(
		.I(MUX_SB_T1_SOUTH_SB_OUT_B1_I),
		.O(MUX_SB_T1_SOUTH_SB_OUT_B1_O),
		.ready_in(SB_T1_SOUTH_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T1_SOUTH_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T1_SOUTH_SB_OUT_B1_valid_out),
		.S(SB_T1_SOUTH_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T1_WEST_SB_OUT_B1_I;
	assign MUX_SB_T1_WEST_SB_OUT_B1_I[5+:1] = PondTop_output_width_1_num_1;
	assign MUX_SB_T1_WEST_SB_OUT_B1_I[4+:1] = PondTop_output_width_1_num_0;
	assign MUX_SB_T1_WEST_SB_OUT_B1_I[3+:1] = PE_output_width_1_num_0;
	assign MUX_SB_T1_WEST_SB_OUT_B1_I[2+:1] = WIRE_SB_T1_EAST_SB_IN_B1_O;
	assign MUX_SB_T1_WEST_SB_OUT_B1_I[1+:1] = WIRE_SB_T0_SOUTH_SB_IN_B1_O;
	assign MUX_SB_T1_WEST_SB_OUT_B1_I[0+:1] = WIRE_SB_T4_NORTH_SB_IN_B1_O;
	wire [5:0] MUX_SB_T1_WEST_SB_OUT_B1_valid_in;
	assign MUX_SB_T1_WEST_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid, PondTop_output_width_1_num_0_valid, PE_output_width_1_num_0_valid, WIRE_SB_T1_EAST_SB_IN_B1_valid_out, WIRE_SB_T0_SOUTH_SB_IN_B1_valid_out, WIRE_SB_T4_NORTH_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T1_WEST_SB_OUT_B1(
		.I(MUX_SB_T1_WEST_SB_OUT_B1_I),
		.O(MUX_SB_T1_WEST_SB_OUT_B1_O),
		.ready_in(SB_T1_WEST_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T1_WEST_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T1_WEST_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T1_WEST_SB_OUT_B1_valid_out),
		.S(SB_T1_WEST_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T1_WEST_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T2_EAST_SB_OUT_B1_I;
	assign MUX_SB_T2_EAST_SB_OUT_B1_I[5+:1] = PondTop_output_width_1_num_1;
	assign MUX_SB_T2_EAST_SB_OUT_B1_I[4+:1] = PondTop_output_width_1_num_0;
	assign MUX_SB_T2_EAST_SB_OUT_B1_I[3+:1] = PE_output_width_1_num_0;
	assign MUX_SB_T2_EAST_SB_OUT_B1_I[2+:1] = WIRE_SB_T2_WEST_SB_IN_B1_O;
	assign MUX_SB_T2_EAST_SB_OUT_B1_I[1+:1] = WIRE_SB_T1_SOUTH_SB_IN_B1_O;
	assign MUX_SB_T2_EAST_SB_OUT_B1_I[0+:1] = WIRE_SB_T1_NORTH_SB_IN_B1_O;
	wire [5:0] MUX_SB_T2_EAST_SB_OUT_B1_valid_in;
	assign MUX_SB_T2_EAST_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid, PondTop_output_width_1_num_0_valid, PE_output_width_1_num_0_valid, WIRE_SB_T2_WEST_SB_IN_B1_valid_out, WIRE_SB_T1_SOUTH_SB_IN_B1_valid_out, WIRE_SB_T1_NORTH_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T2_EAST_SB_OUT_B1(
		.I(MUX_SB_T2_EAST_SB_OUT_B1_I),
		.O(MUX_SB_T2_EAST_SB_OUT_B1_O),
		.ready_in(SB_T2_EAST_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T2_EAST_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T2_EAST_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T2_EAST_SB_OUT_B1_valid_out),
		.S(SB_T2_EAST_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T2_EAST_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T2_NORTH_SB_OUT_B1_I;
	assign MUX_SB_T2_NORTH_SB_OUT_B1_I[5+:1] = PondTop_output_width_1_num_1;
	assign MUX_SB_T2_NORTH_SB_OUT_B1_I[4+:1] = PondTop_output_width_1_num_0;
	assign MUX_SB_T2_NORTH_SB_OUT_B1_I[3+:1] = PE_output_width_1_num_0;
	assign MUX_SB_T2_NORTH_SB_OUT_B1_I[2+:1] = WIRE_SB_T3_WEST_SB_IN_B1_O;
	assign MUX_SB_T2_NORTH_SB_OUT_B1_I[1+:1] = WIRE_SB_T2_SOUTH_SB_IN_B1_O;
	assign MUX_SB_T2_NORTH_SB_OUT_B1_I[0+:1] = WIRE_SB_T3_EAST_SB_IN_B1_O;
	wire [5:0] MUX_SB_T2_NORTH_SB_OUT_B1_valid_in;
	assign MUX_SB_T2_NORTH_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid, PondTop_output_width_1_num_0_valid, PE_output_width_1_num_0_valid, WIRE_SB_T3_WEST_SB_IN_B1_valid_out, WIRE_SB_T2_SOUTH_SB_IN_B1_valid_out, WIRE_SB_T3_EAST_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T2_NORTH_SB_OUT_B1(
		.I(MUX_SB_T2_NORTH_SB_OUT_B1_I),
		.O(MUX_SB_T2_NORTH_SB_OUT_B1_O),
		.ready_in(SB_T2_NORTH_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T2_NORTH_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T2_NORTH_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T2_NORTH_SB_OUT_B1_valid_out),
		.S(SB_T2_NORTH_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T2_NORTH_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T2_SOUTH_SB_OUT_B1_I;
	assign MUX_SB_T2_SOUTH_SB_OUT_B1_I[5+:1] = PondTop_output_width_1_num_1;
	assign MUX_SB_T2_SOUTH_SB_OUT_B1_I[4+:1] = PondTop_output_width_1_num_0;
	assign MUX_SB_T2_SOUTH_SB_OUT_B1_I[3+:1] = PE_output_width_1_num_0;
	assign MUX_SB_T2_SOUTH_SB_OUT_B1_I[2+:1] = WIRE_SB_T3_WEST_SB_IN_B1_O;
	assign MUX_SB_T2_SOUTH_SB_OUT_B1_I[1+:1] = WIRE_SB_T2_NORTH_SB_IN_B1_O;
	assign MUX_SB_T2_SOUTH_SB_OUT_B1_I[0+:1] = WIRE_SB_T1_EAST_SB_IN_B1_O;
	wire [5:0] MUX_SB_T2_SOUTH_SB_OUT_B1_valid_in;
	assign MUX_SB_T2_SOUTH_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid, PondTop_output_width_1_num_0_valid, PE_output_width_1_num_0_valid, WIRE_SB_T3_WEST_SB_IN_B1_valid_out, WIRE_SB_T2_NORTH_SB_IN_B1_valid_out, WIRE_SB_T1_EAST_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T2_SOUTH_SB_OUT_B1(
		.I(MUX_SB_T2_SOUTH_SB_OUT_B1_I),
		.O(MUX_SB_T2_SOUTH_SB_OUT_B1_O),
		.ready_in(SB_T2_SOUTH_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T2_SOUTH_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T2_SOUTH_SB_OUT_B1_valid_out),
		.S(SB_T2_SOUTH_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T2_WEST_SB_OUT_B1_I;
	assign MUX_SB_T2_WEST_SB_OUT_B1_I[5+:1] = PondTop_output_width_1_num_1;
	assign MUX_SB_T2_WEST_SB_OUT_B1_I[4+:1] = PondTop_output_width_1_num_0;
	assign MUX_SB_T2_WEST_SB_OUT_B1_I[3+:1] = PE_output_width_1_num_0;
	assign MUX_SB_T2_WEST_SB_OUT_B1_I[2+:1] = WIRE_SB_T2_EAST_SB_IN_B1_O;
	assign MUX_SB_T2_WEST_SB_OUT_B1_I[1+:1] = WIRE_SB_T1_SOUTH_SB_IN_B1_O;
	assign MUX_SB_T2_WEST_SB_OUT_B1_I[0+:1] = WIRE_SB_T3_NORTH_SB_IN_B1_O;
	wire [5:0] MUX_SB_T2_WEST_SB_OUT_B1_valid_in;
	assign MUX_SB_T2_WEST_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid, PondTop_output_width_1_num_0_valid, PE_output_width_1_num_0_valid, WIRE_SB_T2_EAST_SB_IN_B1_valid_out, WIRE_SB_T1_SOUTH_SB_IN_B1_valid_out, WIRE_SB_T3_NORTH_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T2_WEST_SB_OUT_B1(
		.I(MUX_SB_T2_WEST_SB_OUT_B1_I),
		.O(MUX_SB_T2_WEST_SB_OUT_B1_O),
		.ready_in(SB_T2_WEST_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T2_WEST_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T2_WEST_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T2_WEST_SB_OUT_B1_valid_out),
		.S(SB_T2_WEST_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T2_WEST_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T3_EAST_SB_OUT_B1_I;
	assign MUX_SB_T3_EAST_SB_OUT_B1_I[5+:1] = PondTop_output_width_1_num_1;
	assign MUX_SB_T3_EAST_SB_OUT_B1_I[4+:1] = PondTop_output_width_1_num_0;
	assign MUX_SB_T3_EAST_SB_OUT_B1_I[3+:1] = PE_output_width_1_num_0;
	assign MUX_SB_T3_EAST_SB_OUT_B1_I[2+:1] = WIRE_SB_T3_WEST_SB_IN_B1_O;
	assign MUX_SB_T3_EAST_SB_OUT_B1_I[1+:1] = WIRE_SB_T2_NORTH_SB_IN_B1_O;
	assign MUX_SB_T3_EAST_SB_OUT_B1_I[0+:1] = WIRE_SB_T0_SOUTH_SB_IN_B1_O;
	wire [5:0] MUX_SB_T3_EAST_SB_OUT_B1_valid_in;
	assign MUX_SB_T3_EAST_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid, PondTop_output_width_1_num_0_valid, PE_output_width_1_num_0_valid, WIRE_SB_T3_WEST_SB_IN_B1_valid_out, WIRE_SB_T2_NORTH_SB_IN_B1_valid_out, WIRE_SB_T0_SOUTH_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T3_EAST_SB_OUT_B1(
		.I(MUX_SB_T3_EAST_SB_OUT_B1_I),
		.O(MUX_SB_T3_EAST_SB_OUT_B1_O),
		.ready_in(SB_T3_EAST_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T3_EAST_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T3_EAST_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T3_EAST_SB_OUT_B1_valid_out),
		.S(SB_T3_EAST_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T3_EAST_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T3_NORTH_SB_OUT_B1_I;
	assign MUX_SB_T3_NORTH_SB_OUT_B1_I[5+:1] = PondTop_output_width_1_num_1;
	assign MUX_SB_T3_NORTH_SB_OUT_B1_I[4+:1] = PondTop_output_width_1_num_0;
	assign MUX_SB_T3_NORTH_SB_OUT_B1_I[3+:1] = PE_output_width_1_num_0;
	assign MUX_SB_T3_NORTH_SB_OUT_B1_I[2+:1] = WIRE_SB_T3_SOUTH_SB_IN_B1_O;
	assign MUX_SB_T3_NORTH_SB_OUT_B1_I[1+:1] = WIRE_SB_T4_EAST_SB_IN_B1_O;
	assign MUX_SB_T3_NORTH_SB_OUT_B1_I[0+:1] = WIRE_SB_T2_WEST_SB_IN_B1_O;
	wire [5:0] MUX_SB_T3_NORTH_SB_OUT_B1_valid_in;
	assign MUX_SB_T3_NORTH_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid, PondTop_output_width_1_num_0_valid, PE_output_width_1_num_0_valid, WIRE_SB_T3_SOUTH_SB_IN_B1_valid_out, WIRE_SB_T4_EAST_SB_IN_B1_valid_out, WIRE_SB_T2_WEST_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T3_NORTH_SB_OUT_B1(
		.I(MUX_SB_T3_NORTH_SB_OUT_B1_I),
		.O(MUX_SB_T3_NORTH_SB_OUT_B1_O),
		.ready_in(SB_T3_NORTH_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T3_NORTH_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T3_NORTH_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T3_NORTH_SB_OUT_B1_valid_out),
		.S(SB_T3_NORTH_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T3_NORTH_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T3_SOUTH_SB_OUT_B1_I;
	assign MUX_SB_T3_SOUTH_SB_OUT_B1_I[5+:1] = PondTop_output_width_1_num_1;
	assign MUX_SB_T3_SOUTH_SB_OUT_B1_I[4+:1] = PondTop_output_width_1_num_0;
	assign MUX_SB_T3_SOUTH_SB_OUT_B1_I[3+:1] = PE_output_width_1_num_0;
	assign MUX_SB_T3_SOUTH_SB_OUT_B1_I[2+:1] = WIRE_SB_T4_WEST_SB_IN_B1_O;
	assign MUX_SB_T3_SOUTH_SB_OUT_B1_I[1+:1] = WIRE_SB_T3_NORTH_SB_IN_B1_O;
	assign MUX_SB_T3_SOUTH_SB_OUT_B1_I[0+:1] = WIRE_SB_T0_EAST_SB_IN_B1_O;
	wire [5:0] MUX_SB_T3_SOUTH_SB_OUT_B1_valid_in;
	assign MUX_SB_T3_SOUTH_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid, PondTop_output_width_1_num_0_valid, PE_output_width_1_num_0_valid, WIRE_SB_T4_WEST_SB_IN_B1_valid_out, WIRE_SB_T3_NORTH_SB_IN_B1_valid_out, WIRE_SB_T0_EAST_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T3_SOUTH_SB_OUT_B1(
		.I(MUX_SB_T3_SOUTH_SB_OUT_B1_I),
		.O(MUX_SB_T3_SOUTH_SB_OUT_B1_O),
		.ready_in(SB_T3_SOUTH_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T3_SOUTH_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T3_SOUTH_SB_OUT_B1_valid_out),
		.S(SB_T3_SOUTH_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T3_WEST_SB_OUT_B1_I;
	assign MUX_SB_T3_WEST_SB_OUT_B1_I[5+:1] = PondTop_output_width_1_num_1;
	assign MUX_SB_T3_WEST_SB_OUT_B1_I[4+:1] = PondTop_output_width_1_num_0;
	assign MUX_SB_T3_WEST_SB_OUT_B1_I[3+:1] = PE_output_width_1_num_0;
	assign MUX_SB_T3_WEST_SB_OUT_B1_I[2+:1] = WIRE_SB_T3_EAST_SB_IN_B1_O;
	assign MUX_SB_T3_WEST_SB_OUT_B1_I[1+:1] = WIRE_SB_T2_SOUTH_SB_IN_B1_O;
	assign MUX_SB_T3_WEST_SB_OUT_B1_I[0+:1] = WIRE_SB_T2_NORTH_SB_IN_B1_O;
	wire [5:0] MUX_SB_T3_WEST_SB_OUT_B1_valid_in;
	assign MUX_SB_T3_WEST_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid, PondTop_output_width_1_num_0_valid, PE_output_width_1_num_0_valid, WIRE_SB_T3_EAST_SB_IN_B1_valid_out, WIRE_SB_T2_SOUTH_SB_IN_B1_valid_out, WIRE_SB_T2_NORTH_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T3_WEST_SB_OUT_B1(
		.I(MUX_SB_T3_WEST_SB_OUT_B1_I),
		.O(MUX_SB_T3_WEST_SB_OUT_B1_O),
		.ready_in(SB_T3_WEST_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T3_WEST_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T3_WEST_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T3_WEST_SB_OUT_B1_valid_out),
		.S(SB_T3_WEST_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T3_WEST_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T4_EAST_SB_OUT_B1_I;
	assign MUX_SB_T4_EAST_SB_OUT_B1_I[5+:1] = PondTop_output_width_1_num_1;
	assign MUX_SB_T4_EAST_SB_OUT_B1_I[4+:1] = PondTop_output_width_1_num_0;
	assign MUX_SB_T4_EAST_SB_OUT_B1_I[3+:1] = PE_output_width_1_num_0;
	assign MUX_SB_T4_EAST_SB_OUT_B1_I[2+:1] = WIRE_SB_T4_WEST_SB_IN_B1_O;
	assign MUX_SB_T4_EAST_SB_OUT_B1_I[1+:1] = WIRE_SB_T4_SOUTH_SB_IN_B1_O;
	assign MUX_SB_T4_EAST_SB_OUT_B1_I[0+:1] = WIRE_SB_T3_NORTH_SB_IN_B1_O;
	wire [5:0] MUX_SB_T4_EAST_SB_OUT_B1_valid_in;
	assign MUX_SB_T4_EAST_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid, PondTop_output_width_1_num_0_valid, PE_output_width_1_num_0_valid, WIRE_SB_T4_WEST_SB_IN_B1_valid_out, WIRE_SB_T4_SOUTH_SB_IN_B1_valid_out, WIRE_SB_T3_NORTH_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T4_EAST_SB_OUT_B1(
		.I(MUX_SB_T4_EAST_SB_OUT_B1_I),
		.O(MUX_SB_T4_EAST_SB_OUT_B1_O),
		.ready_in(SB_T4_EAST_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T4_EAST_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T4_EAST_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T4_EAST_SB_OUT_B1_valid_out),
		.S(SB_T4_EAST_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T4_EAST_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T4_NORTH_SB_OUT_B1_I;
	assign MUX_SB_T4_NORTH_SB_OUT_B1_I[5+:1] = PondTop_output_width_1_num_1;
	assign MUX_SB_T4_NORTH_SB_OUT_B1_I[4+:1] = PondTop_output_width_1_num_0;
	assign MUX_SB_T4_NORTH_SB_OUT_B1_I[3+:1] = PE_output_width_1_num_0;
	assign MUX_SB_T4_NORTH_SB_OUT_B1_I[2+:1] = WIRE_SB_T4_SOUTH_SB_IN_B1_O;
	assign MUX_SB_T4_NORTH_SB_OUT_B1_I[1+:1] = WIRE_SB_T0_EAST_SB_IN_B1_O;
	assign MUX_SB_T4_NORTH_SB_OUT_B1_I[0+:1] = WIRE_SB_T1_WEST_SB_IN_B1_O;
	wire [5:0] MUX_SB_T4_NORTH_SB_OUT_B1_valid_in;
	assign MUX_SB_T4_NORTH_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid, PondTop_output_width_1_num_0_valid, PE_output_width_1_num_0_valid, WIRE_SB_T4_SOUTH_SB_IN_B1_valid_out, WIRE_SB_T0_EAST_SB_IN_B1_valid_out, WIRE_SB_T1_WEST_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T4_NORTH_SB_OUT_B1(
		.I(MUX_SB_T4_NORTH_SB_OUT_B1_I),
		.O(MUX_SB_T4_NORTH_SB_OUT_B1_O),
		.ready_in(SB_T4_NORTH_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T4_NORTH_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T4_NORTH_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T4_NORTH_SB_OUT_B1_valid_out),
		.S(SB_T4_NORTH_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T4_NORTH_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T4_SOUTH_SB_OUT_B1_I;
	assign MUX_SB_T4_SOUTH_SB_OUT_B1_I[5+:1] = PondTop_output_width_1_num_1;
	assign MUX_SB_T4_SOUTH_SB_OUT_B1_I[4+:1] = PondTop_output_width_1_num_0;
	assign MUX_SB_T4_SOUTH_SB_OUT_B1_I[3+:1] = PE_output_width_1_num_0;
	assign MUX_SB_T4_SOUTH_SB_OUT_B1_I[2+:1] = WIRE_SB_T4_NORTH_SB_IN_B1_O;
	assign MUX_SB_T4_SOUTH_SB_OUT_B1_I[1+:1] = WIRE_SB_T4_EAST_SB_IN_B1_O;
	assign MUX_SB_T4_SOUTH_SB_OUT_B1_I[0+:1] = WIRE_SB_T0_WEST_SB_IN_B1_O;
	wire [5:0] MUX_SB_T4_SOUTH_SB_OUT_B1_valid_in;
	assign MUX_SB_T4_SOUTH_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid, PondTop_output_width_1_num_0_valid, PE_output_width_1_num_0_valid, WIRE_SB_T4_NORTH_SB_IN_B1_valid_out, WIRE_SB_T4_EAST_SB_IN_B1_valid_out, WIRE_SB_T0_WEST_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T4_SOUTH_SB_OUT_B1(
		.I(MUX_SB_T4_SOUTH_SB_OUT_B1_I),
		.O(MUX_SB_T4_SOUTH_SB_OUT_B1_O),
		.ready_in(SB_T4_SOUTH_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T4_SOUTH_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T4_SOUTH_SB_OUT_B1_valid_out),
		.S(SB_T4_SOUTH_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T4_WEST_SB_OUT_B1_I;
	assign MUX_SB_T4_WEST_SB_OUT_B1_I[5+:1] = PondTop_output_width_1_num_1;
	assign MUX_SB_T4_WEST_SB_OUT_B1_I[4+:1] = PondTop_output_width_1_num_0;
	assign MUX_SB_T4_WEST_SB_OUT_B1_I[3+:1] = PE_output_width_1_num_0;
	assign MUX_SB_T4_WEST_SB_OUT_B1_I[2+:1] = WIRE_SB_T4_EAST_SB_IN_B1_O;
	assign MUX_SB_T4_WEST_SB_OUT_B1_I[1+:1] = WIRE_SB_T3_SOUTH_SB_IN_B1_O;
	assign MUX_SB_T4_WEST_SB_OUT_B1_I[0+:1] = WIRE_SB_T1_NORTH_SB_IN_B1_O;
	wire [5:0] MUX_SB_T4_WEST_SB_OUT_B1_valid_in;
	assign MUX_SB_T4_WEST_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid, PondTop_output_width_1_num_0_valid, PE_output_width_1_num_0_valid, WIRE_SB_T4_EAST_SB_IN_B1_valid_out, WIRE_SB_T3_SOUTH_SB_IN_B1_valid_out, WIRE_SB_T1_NORTH_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T4_WEST_SB_OUT_B1(
		.I(MUX_SB_T4_WEST_SB_OUT_B1_I),
		.O(MUX_SB_T4_WEST_SB_OUT_B1_O),
		.ready_in(SB_T4_WEST_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T4_WEST_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T4_WEST_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T4_WEST_SB_OUT_B1_valid_out),
		.S(SB_T4_WEST_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T4_WEST_SB_OUT_B1_out_sel)
	);
	SplitFifo_1 REG_T0_EAST_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T0_EAST_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T0_EAST_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T0_EAST_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T0_EAST_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst2_out[0]),
		.end_fifo(REG_T0_EAST_B1_end_value_O[0]),
		.valid0(MUX_SB_T0_EAST_SB_OUT_B1_valid_out),
		.valid1(REG_T0_EAST_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T0_EAST_B1_ready_out),
		.fifo_en(REG_T0_EAST_B1_fifo_value_O[0])
	);
	SliceWrapper_32_0_1 REG_T0_EAST_B1_end_value(
		.I(config_reg_0_O),
		.O(REG_T0_EAST_B1_end_value_O)
	);
	SliceWrapper_32_1_2 REG_T0_EAST_B1_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T0_EAST_B1_fifo_value_O)
	);
	SliceWrapper_32_2_3 REG_T0_EAST_B1_start_value(
		.I(config_reg_0_O),
		.O(REG_T0_EAST_B1_start_value_O)
	);
	SplitFifo_1 REG_T0_NORTH_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T0_NORTH_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T0_NORTH_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T0_NORTH_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T0_NORTH_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst0_out[0]),
		.end_fifo(REG_T0_NORTH_B1_end_value_O[0]),
		.valid0(MUX_SB_T0_NORTH_SB_OUT_B1_valid_out),
		.valid1(REG_T0_NORTH_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T0_NORTH_B1_ready_out),
		.fifo_en(REG_T0_NORTH_B1_fifo_value_O[0])
	);
	SliceWrapper_32_3_4 REG_T0_NORTH_B1_end_value(
		.I(config_reg_0_O),
		.O(REG_T0_NORTH_B1_end_value_O)
	);
	SliceWrapper_32_4_5 REG_T0_NORTH_B1_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T0_NORTH_B1_fifo_value_O)
	);
	SliceWrapper_32_5_6 REG_T0_NORTH_B1_start_value(
		.I(config_reg_0_O),
		.O(REG_T0_NORTH_B1_start_value_O)
	);
	SplitFifo_1 REG_T0_SOUTH_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T0_SOUTH_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T0_SOUTH_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T0_SOUTH_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T0_SOUTH_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst1_out[0]),
		.end_fifo(REG_T0_SOUTH_B1_end_value_O[0]),
		.valid0(MUX_SB_T0_SOUTH_SB_OUT_B1_valid_out),
		.valid1(REG_T0_SOUTH_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T0_SOUTH_B1_ready_out),
		.fifo_en(REG_T0_SOUTH_B1_fifo_value_O[0])
	);
	SliceWrapper_32_6_7 REG_T0_SOUTH_B1_end_value(
		.I(config_reg_0_O),
		.O(REG_T0_SOUTH_B1_end_value_O)
	);
	SliceWrapper_32_7_8 REG_T0_SOUTH_B1_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T0_SOUTH_B1_fifo_value_O)
	);
	SliceWrapper_32_8_9 REG_T0_SOUTH_B1_start_value(
		.I(config_reg_0_O),
		.O(REG_T0_SOUTH_B1_start_value_O)
	);
	SplitFifo_1 REG_T0_WEST_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T0_WEST_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T0_WEST_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T0_WEST_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T0_WEST_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst3_out[0]),
		.end_fifo(REG_T0_WEST_B1_end_value_O[0]),
		.valid0(MUX_SB_T0_WEST_SB_OUT_B1_valid_out),
		.valid1(REG_T0_WEST_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T0_WEST_B1_ready_out),
		.fifo_en(REG_T0_WEST_B1_fifo_value_O[0])
	);
	SliceWrapper_32_9_10 REG_T0_WEST_B1_end_value(
		.I(config_reg_0_O),
		.O(REG_T0_WEST_B1_end_value_O)
	);
	SliceWrapper_32_10_11 REG_T0_WEST_B1_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T0_WEST_B1_fifo_value_O)
	);
	SliceWrapper_32_11_12 REG_T0_WEST_B1_start_value(
		.I(config_reg_0_O),
		.O(REG_T0_WEST_B1_start_value_O)
	);
	SplitFifo_1 REG_T1_EAST_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T1_EAST_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T1_EAST_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T1_EAST_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T1_EAST_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst6_out[0]),
		.end_fifo(REG_T1_EAST_B1_end_value_O[0]),
		.valid0(MUX_SB_T1_EAST_SB_OUT_B1_valid_out),
		.valid1(REG_T1_EAST_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T1_EAST_B1_ready_out),
		.fifo_en(REG_T1_EAST_B1_fifo_value_O[0])
	);
	SliceWrapper_32_12_13 REG_T1_EAST_B1_end_value(
		.I(config_reg_0_O),
		.O(REG_T1_EAST_B1_end_value_O)
	);
	SliceWrapper_32_13_14 REG_T1_EAST_B1_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T1_EAST_B1_fifo_value_O)
	);
	SliceWrapper_32_14_15 REG_T1_EAST_B1_start_value(
		.I(config_reg_0_O),
		.O(REG_T1_EAST_B1_start_value_O)
	);
	SplitFifo_1 REG_T1_NORTH_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T1_NORTH_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T1_NORTH_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T1_NORTH_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T1_NORTH_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst4_out[0]),
		.end_fifo(REG_T1_NORTH_B1_end_value_O[0]),
		.valid0(MUX_SB_T1_NORTH_SB_OUT_B1_valid_out),
		.valid1(REG_T1_NORTH_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T1_NORTH_B1_ready_out),
		.fifo_en(REG_T1_NORTH_B1_fifo_value_O[0])
	);
	SliceWrapper_32_15_16 REG_T1_NORTH_B1_end_value(
		.I(config_reg_0_O),
		.O(REG_T1_NORTH_B1_end_value_O)
	);
	SliceWrapper_32_16_17 REG_T1_NORTH_B1_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T1_NORTH_B1_fifo_value_O)
	);
	SliceWrapper_32_17_18 REG_T1_NORTH_B1_start_value(
		.I(config_reg_0_O),
		.O(REG_T1_NORTH_B1_start_value_O)
	);
	SplitFifo_1 REG_T1_SOUTH_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T1_SOUTH_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T1_SOUTH_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T1_SOUTH_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T1_SOUTH_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst5_out[0]),
		.end_fifo(REG_T1_SOUTH_B1_end_value_O[0]),
		.valid0(MUX_SB_T1_SOUTH_SB_OUT_B1_valid_out),
		.valid1(REG_T1_SOUTH_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T1_SOUTH_B1_ready_out),
		.fifo_en(REG_T1_SOUTH_B1_fifo_value_O[0])
	);
	SliceWrapper_32_18_19 REG_T1_SOUTH_B1_end_value(
		.I(config_reg_0_O),
		.O(REG_T1_SOUTH_B1_end_value_O)
	);
	SliceWrapper_32_19_20 REG_T1_SOUTH_B1_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T1_SOUTH_B1_fifo_value_O)
	);
	SliceWrapper_32_20_21 REG_T1_SOUTH_B1_start_value(
		.I(config_reg_0_O),
		.O(REG_T1_SOUTH_B1_start_value_O)
	);
	SplitFifo_1 REG_T1_WEST_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T1_WEST_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T1_WEST_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T1_WEST_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T1_WEST_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst7_out[0]),
		.end_fifo(REG_T1_WEST_B1_end_value_O[0]),
		.valid0(MUX_SB_T1_WEST_SB_OUT_B1_valid_out),
		.valid1(REG_T1_WEST_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T1_WEST_B1_ready_out),
		.fifo_en(REG_T1_WEST_B1_fifo_value_O[0])
	);
	SliceWrapper_32_21_22 REG_T1_WEST_B1_end_value(
		.I(config_reg_0_O),
		.O(REG_T1_WEST_B1_end_value_O)
	);
	SliceWrapper_32_22_23 REG_T1_WEST_B1_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T1_WEST_B1_fifo_value_O)
	);
	SliceWrapper_32_23_24 REG_T1_WEST_B1_start_value(
		.I(config_reg_0_O),
		.O(REG_T1_WEST_B1_start_value_O)
	);
	SplitFifo_1 REG_T2_EAST_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T2_EAST_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T2_EAST_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T2_EAST_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T2_EAST_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst10_out[0]),
		.end_fifo(REG_T2_EAST_B1_end_value_O[0]),
		.valid0(MUX_SB_T2_EAST_SB_OUT_B1_valid_out),
		.valid1(REG_T2_EAST_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T2_EAST_B1_ready_out),
		.fifo_en(REG_T2_EAST_B1_fifo_value_O[0])
	);
	SliceWrapper_32_24_25 REG_T2_EAST_B1_end_value(
		.I(config_reg_0_O),
		.O(REG_T2_EAST_B1_end_value_O)
	);
	SliceWrapper_32_25_26 REG_T2_EAST_B1_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T2_EAST_B1_fifo_value_O)
	);
	SliceWrapper_32_26_27 REG_T2_EAST_B1_start_value(
		.I(config_reg_0_O),
		.O(REG_T2_EAST_B1_start_value_O)
	);
	SplitFifo_1 REG_T2_NORTH_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T2_NORTH_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T2_NORTH_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T2_NORTH_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T2_NORTH_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst8_out[0]),
		.end_fifo(REG_T2_NORTH_B1_end_value_O[0]),
		.valid0(MUX_SB_T2_NORTH_SB_OUT_B1_valid_out),
		.valid1(REG_T2_NORTH_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T2_NORTH_B1_ready_out),
		.fifo_en(REG_T2_NORTH_B1_fifo_value_O[0])
	);
	SliceWrapper_32_27_28 REG_T2_NORTH_B1_end_value(
		.I(config_reg_0_O),
		.O(REG_T2_NORTH_B1_end_value_O)
	);
	SliceWrapper_32_28_29 REG_T2_NORTH_B1_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T2_NORTH_B1_fifo_value_O)
	);
	SliceWrapper_32_29_30 REG_T2_NORTH_B1_start_value(
		.I(config_reg_0_O),
		.O(REG_T2_NORTH_B1_start_value_O)
	);
	SplitFifo_1 REG_T2_SOUTH_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T2_SOUTH_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T2_SOUTH_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T2_SOUTH_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T2_SOUTH_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst9_out[0]),
		.end_fifo(REG_T2_SOUTH_B1_end_value_O[0]),
		.valid0(MUX_SB_T2_SOUTH_SB_OUT_B1_valid_out),
		.valid1(REG_T2_SOUTH_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T2_SOUTH_B1_ready_out),
		.fifo_en(REG_T2_SOUTH_B1_fifo_value_O[0])
	);
	SliceWrapper_32_30_31 REG_T2_SOUTH_B1_end_value(
		.I(config_reg_0_O),
		.O(REG_T2_SOUTH_B1_end_value_O)
	);
	SliceWrapper_32_31_32 REG_T2_SOUTH_B1_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T2_SOUTH_B1_fifo_value_O)
	);
	SliceWrapper_32_0_1 REG_T2_SOUTH_B1_start_value(
		.I(config_reg_1_O),
		.O(REG_T2_SOUTH_B1_start_value_O)
	);
	SplitFifo_1 REG_T2_WEST_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T2_WEST_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T2_WEST_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T2_WEST_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T2_WEST_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst11_out[0]),
		.end_fifo(REG_T2_WEST_B1_end_value_O[0]),
		.valid0(MUX_SB_T2_WEST_SB_OUT_B1_valid_out),
		.valid1(REG_T2_WEST_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T2_WEST_B1_ready_out),
		.fifo_en(REG_T2_WEST_B1_fifo_value_O[0])
	);
	SliceWrapper_32_1_2 REG_T2_WEST_B1_end_value(
		.I(config_reg_1_O),
		.O(REG_T2_WEST_B1_end_value_O)
	);
	SliceWrapper_32_2_3 REG_T2_WEST_B1_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T2_WEST_B1_fifo_value_O)
	);
	SliceWrapper_32_3_4 REG_T2_WEST_B1_start_value(
		.I(config_reg_1_O),
		.O(REG_T2_WEST_B1_start_value_O)
	);
	SplitFifo_1 REG_T3_EAST_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T3_EAST_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T3_EAST_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T3_EAST_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T3_EAST_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst14_out[0]),
		.end_fifo(REG_T3_EAST_B1_end_value_O[0]),
		.valid0(MUX_SB_T3_EAST_SB_OUT_B1_valid_out),
		.valid1(REG_T3_EAST_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T3_EAST_B1_ready_out),
		.fifo_en(REG_T3_EAST_B1_fifo_value_O[0])
	);
	SliceWrapper_32_4_5 REG_T3_EAST_B1_end_value(
		.I(config_reg_1_O),
		.O(REG_T3_EAST_B1_end_value_O)
	);
	SliceWrapper_32_5_6 REG_T3_EAST_B1_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T3_EAST_B1_fifo_value_O)
	);
	SliceWrapper_32_6_7 REG_T3_EAST_B1_start_value(
		.I(config_reg_1_O),
		.O(REG_T3_EAST_B1_start_value_O)
	);
	SplitFifo_1 REG_T3_NORTH_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T3_NORTH_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T3_NORTH_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T3_NORTH_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T3_NORTH_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst12_out[0]),
		.end_fifo(REG_T3_NORTH_B1_end_value_O[0]),
		.valid0(MUX_SB_T3_NORTH_SB_OUT_B1_valid_out),
		.valid1(REG_T3_NORTH_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T3_NORTH_B1_ready_out),
		.fifo_en(REG_T3_NORTH_B1_fifo_value_O[0])
	);
	SliceWrapper_32_7_8 REG_T3_NORTH_B1_end_value(
		.I(config_reg_1_O),
		.O(REG_T3_NORTH_B1_end_value_O)
	);
	SliceWrapper_32_8_9 REG_T3_NORTH_B1_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T3_NORTH_B1_fifo_value_O)
	);
	SliceWrapper_32_9_10 REG_T3_NORTH_B1_start_value(
		.I(config_reg_1_O),
		.O(REG_T3_NORTH_B1_start_value_O)
	);
	SplitFifo_1 REG_T3_SOUTH_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T3_SOUTH_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T3_SOUTH_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T3_SOUTH_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T3_SOUTH_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst13_out[0]),
		.end_fifo(REG_T3_SOUTH_B1_end_value_O[0]),
		.valid0(MUX_SB_T3_SOUTH_SB_OUT_B1_valid_out),
		.valid1(REG_T3_SOUTH_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T3_SOUTH_B1_ready_out),
		.fifo_en(REG_T3_SOUTH_B1_fifo_value_O[0])
	);
	SliceWrapper_32_10_11 REG_T3_SOUTH_B1_end_value(
		.I(config_reg_1_O),
		.O(REG_T3_SOUTH_B1_end_value_O)
	);
	SliceWrapper_32_11_12 REG_T3_SOUTH_B1_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T3_SOUTH_B1_fifo_value_O)
	);
	SliceWrapper_32_12_13 REG_T3_SOUTH_B1_start_value(
		.I(config_reg_1_O),
		.O(REG_T3_SOUTH_B1_start_value_O)
	);
	SplitFifo_1 REG_T3_WEST_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T3_WEST_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T3_WEST_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T3_WEST_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T3_WEST_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst15_out[0]),
		.end_fifo(REG_T3_WEST_B1_end_value_O[0]),
		.valid0(MUX_SB_T3_WEST_SB_OUT_B1_valid_out),
		.valid1(REG_T3_WEST_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T3_WEST_B1_ready_out),
		.fifo_en(REG_T3_WEST_B1_fifo_value_O[0])
	);
	SliceWrapper_32_13_14 REG_T3_WEST_B1_end_value(
		.I(config_reg_1_O),
		.O(REG_T3_WEST_B1_end_value_O)
	);
	SliceWrapper_32_14_15 REG_T3_WEST_B1_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T3_WEST_B1_fifo_value_O)
	);
	SliceWrapper_32_15_16 REG_T3_WEST_B1_start_value(
		.I(config_reg_1_O),
		.O(REG_T3_WEST_B1_start_value_O)
	);
	SplitFifo_1 REG_T4_EAST_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T4_EAST_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T4_EAST_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T4_EAST_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T4_EAST_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst18_out[0]),
		.end_fifo(REG_T4_EAST_B1_end_value_O[0]),
		.valid0(MUX_SB_T4_EAST_SB_OUT_B1_valid_out),
		.valid1(REG_T4_EAST_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T4_EAST_B1_ready_out),
		.fifo_en(REG_T4_EAST_B1_fifo_value_O[0])
	);
	SliceWrapper_32_16_17 REG_T4_EAST_B1_end_value(
		.I(config_reg_1_O),
		.O(REG_T4_EAST_B1_end_value_O)
	);
	SliceWrapper_32_17_18 REG_T4_EAST_B1_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T4_EAST_B1_fifo_value_O)
	);
	SliceWrapper_32_18_19 REG_T4_EAST_B1_start_value(
		.I(config_reg_1_O),
		.O(REG_T4_EAST_B1_start_value_O)
	);
	SplitFifo_1 REG_T4_NORTH_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T4_NORTH_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T4_NORTH_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T4_NORTH_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T4_NORTH_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst16_out[0]),
		.end_fifo(REG_T4_NORTH_B1_end_value_O[0]),
		.valid0(MUX_SB_T4_NORTH_SB_OUT_B1_valid_out),
		.valid1(REG_T4_NORTH_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T4_NORTH_B1_ready_out),
		.fifo_en(REG_T4_NORTH_B1_fifo_value_O[0])
	);
	SliceWrapper_32_19_20 REG_T4_NORTH_B1_end_value(
		.I(config_reg_1_O),
		.O(REG_T4_NORTH_B1_end_value_O)
	);
	SliceWrapper_32_20_21 REG_T4_NORTH_B1_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T4_NORTH_B1_fifo_value_O)
	);
	SliceWrapper_32_21_22 REG_T4_NORTH_B1_start_value(
		.I(config_reg_1_O),
		.O(REG_T4_NORTH_B1_start_value_O)
	);
	SplitFifo_1 REG_T4_SOUTH_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T4_SOUTH_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T4_SOUTH_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T4_SOUTH_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T4_SOUTH_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst17_out[0]),
		.end_fifo(REG_T4_SOUTH_B1_end_value_O[0]),
		.valid0(MUX_SB_T4_SOUTH_SB_OUT_B1_valid_out),
		.valid1(REG_T4_SOUTH_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T4_SOUTH_B1_ready_out),
		.fifo_en(REG_T4_SOUTH_B1_fifo_value_O[0])
	);
	SliceWrapper_32_22_23 REG_T4_SOUTH_B1_end_value(
		.I(config_reg_1_O),
		.O(REG_T4_SOUTH_B1_end_value_O)
	);
	SliceWrapper_32_23_24 REG_T4_SOUTH_B1_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T4_SOUTH_B1_fifo_value_O)
	);
	SliceWrapper_32_24_25 REG_T4_SOUTH_B1_start_value(
		.I(config_reg_1_O),
		.O(REG_T4_SOUTH_B1_start_value_O)
	);
	SplitFifo_1 REG_T4_WEST_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T4_WEST_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T4_WEST_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T4_WEST_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T4_WEST_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst19_out[0]),
		.end_fifo(REG_T4_WEST_B1_end_value_O[0]),
		.valid0(MUX_SB_T4_WEST_SB_OUT_B1_valid_out),
		.valid1(REG_T4_WEST_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T4_WEST_B1_ready_out),
		.fifo_en(REG_T4_WEST_B1_fifo_value_O[0])
	);
	SliceWrapper_32_25_26 REG_T4_WEST_B1_end_value(
		.I(config_reg_1_O),
		.O(REG_T4_WEST_B1_end_value_O)
	);
	SliceWrapper_32_26_27 REG_T4_WEST_B1_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T4_WEST_B1_fifo_value_O)
	);
	SliceWrapper_32_27_28 REG_T4_WEST_B1_start_value(
		.I(config_reg_1_O),
		.O(REG_T4_WEST_B1_start_value_O)
	);
	wire [1:0] RMUX_T0_EAST_B1_I;
	assign RMUX_T0_EAST_B1_I[1+:1] = REG_T0_EAST_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T0_EAST_B1_I[0+:1] = MUX_SB_T0_EAST_SB_OUT_B1_O;
	wire [1:0] RMUX_T0_EAST_B1_valid_in;
	assign RMUX_T0_EAST_B1_valid_in = {REG_T0_EAST_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T0_EAST_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T0_EAST_B1(
		.I(RMUX_T0_EAST_B1_I),
		.O(RMUX_T0_EAST_B1_O),
		.ready_in(SB_T0_EAST_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T0_EAST_B1_ready_out),
		.valid_in(RMUX_T0_EAST_B1_valid_in),
		.valid_out(RMUX_T0_EAST_B1_valid_out),
		.S(RMUX_T0_EAST_B1_sel_value_O),
		.out_sel(RMUX_T0_EAST_B1_out_sel)
	);
	SliceWrapper_32_28_29 RMUX_T0_EAST_B1_sel_value(
		.I(config_reg_1_O),
		.O(RMUX_T0_EAST_B1_sel_value_O)
	);
	wire [1:0] RMUX_T0_NORTH_B1_I;
	assign RMUX_T0_NORTH_B1_I[1+:1] = REG_T0_NORTH_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T0_NORTH_B1_I[0+:1] = MUX_SB_T0_NORTH_SB_OUT_B1_O;
	wire [1:0] RMUX_T0_NORTH_B1_valid_in;
	assign RMUX_T0_NORTH_B1_valid_in = {REG_T0_NORTH_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T0_NORTH_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T0_NORTH_B1(
		.I(RMUX_T0_NORTH_B1_I),
		.O(RMUX_T0_NORTH_B1_O),
		.ready_in(SB_T0_NORTH_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T0_NORTH_B1_ready_out),
		.valid_in(RMUX_T0_NORTH_B1_valid_in),
		.valid_out(RMUX_T0_NORTH_B1_valid_out),
		.S(RMUX_T0_NORTH_B1_sel_value_O),
		.out_sel(RMUX_T0_NORTH_B1_out_sel)
	);
	SliceWrapper_32_29_30 RMUX_T0_NORTH_B1_sel_value(
		.I(config_reg_1_O),
		.O(RMUX_T0_NORTH_B1_sel_value_O)
	);
	wire [1:0] RMUX_T0_SOUTH_B1_I;
	assign RMUX_T0_SOUTH_B1_I[1+:1] = REG_T0_SOUTH_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T0_SOUTH_B1_I[0+:1] = MUX_SB_T0_SOUTH_SB_OUT_B1_O;
	wire [1:0] RMUX_T0_SOUTH_B1_valid_in;
	assign RMUX_T0_SOUTH_B1_valid_in = {REG_T0_SOUTH_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T0_SOUTH_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T0_SOUTH_B1(
		.I(RMUX_T0_SOUTH_B1_I),
		.O(RMUX_T0_SOUTH_B1_O),
		.ready_in(SB_T0_SOUTH_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T0_SOUTH_B1_ready_out),
		.valid_in(RMUX_T0_SOUTH_B1_valid_in),
		.valid_out(RMUX_T0_SOUTH_B1_valid_out),
		.S(RMUX_T0_SOUTH_B1_sel_value_O),
		.out_sel(RMUX_T0_SOUTH_B1_out_sel)
	);
	SliceWrapper_32_30_31 RMUX_T0_SOUTH_B1_sel_value(
		.I(config_reg_1_O),
		.O(RMUX_T0_SOUTH_B1_sel_value_O)
	);
	wire [1:0] RMUX_T0_WEST_B1_I;
	assign RMUX_T0_WEST_B1_I[1+:1] = REG_T0_WEST_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T0_WEST_B1_I[0+:1] = MUX_SB_T0_WEST_SB_OUT_B1_O;
	wire [1:0] RMUX_T0_WEST_B1_valid_in;
	assign RMUX_T0_WEST_B1_valid_in = {REG_T0_WEST_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T0_WEST_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T0_WEST_B1(
		.I(RMUX_T0_WEST_B1_I),
		.O(RMUX_T0_WEST_B1_O),
		.ready_in(SB_T0_WEST_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T0_WEST_B1_ready_out),
		.valid_in(RMUX_T0_WEST_B1_valid_in),
		.valid_out(RMUX_T0_WEST_B1_valid_out),
		.S(RMUX_T0_WEST_B1_sel_value_O),
		.out_sel(RMUX_T0_WEST_B1_out_sel)
	);
	SliceWrapper_32_31_32 RMUX_T0_WEST_B1_sel_value(
		.I(config_reg_1_O),
		.O(RMUX_T0_WEST_B1_sel_value_O)
	);
	wire [1:0] RMUX_T1_EAST_B1_I;
	assign RMUX_T1_EAST_B1_I[1+:1] = REG_T1_EAST_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T1_EAST_B1_I[0+:1] = MUX_SB_T1_EAST_SB_OUT_B1_O;
	wire [1:0] RMUX_T1_EAST_B1_valid_in;
	assign RMUX_T1_EAST_B1_valid_in = {REG_T1_EAST_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T1_EAST_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T1_EAST_B1(
		.I(RMUX_T1_EAST_B1_I),
		.O(RMUX_T1_EAST_B1_O),
		.ready_in(SB_T1_EAST_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T1_EAST_B1_ready_out),
		.valid_in(RMUX_T1_EAST_B1_valid_in),
		.valid_out(RMUX_T1_EAST_B1_valid_out),
		.S(RMUX_T1_EAST_B1_sel_value_O),
		.out_sel(RMUX_T1_EAST_B1_out_sel)
	);
	SliceWrapper_32_0_1 RMUX_T1_EAST_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T1_EAST_B1_sel_value_O)
	);
	wire [1:0] RMUX_T1_NORTH_B1_I;
	assign RMUX_T1_NORTH_B1_I[1+:1] = REG_T1_NORTH_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T1_NORTH_B1_I[0+:1] = MUX_SB_T1_NORTH_SB_OUT_B1_O;
	wire [1:0] RMUX_T1_NORTH_B1_valid_in;
	assign RMUX_T1_NORTH_B1_valid_in = {REG_T1_NORTH_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T1_NORTH_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T1_NORTH_B1(
		.I(RMUX_T1_NORTH_B1_I),
		.O(RMUX_T1_NORTH_B1_O),
		.ready_in(SB_T1_NORTH_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T1_NORTH_B1_ready_out),
		.valid_in(RMUX_T1_NORTH_B1_valid_in),
		.valid_out(RMUX_T1_NORTH_B1_valid_out),
		.S(RMUX_T1_NORTH_B1_sel_value_O),
		.out_sel(RMUX_T1_NORTH_B1_out_sel)
	);
	SliceWrapper_32_1_2 RMUX_T1_NORTH_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T1_NORTH_B1_sel_value_O)
	);
	wire [1:0] RMUX_T1_SOUTH_B1_I;
	assign RMUX_T1_SOUTH_B1_I[1+:1] = REG_T1_SOUTH_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T1_SOUTH_B1_I[0+:1] = MUX_SB_T1_SOUTH_SB_OUT_B1_O;
	wire [1:0] RMUX_T1_SOUTH_B1_valid_in;
	assign RMUX_T1_SOUTH_B1_valid_in = {REG_T1_SOUTH_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T1_SOUTH_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T1_SOUTH_B1(
		.I(RMUX_T1_SOUTH_B1_I),
		.O(RMUX_T1_SOUTH_B1_O),
		.ready_in(SB_T1_SOUTH_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T1_SOUTH_B1_ready_out),
		.valid_in(RMUX_T1_SOUTH_B1_valid_in),
		.valid_out(RMUX_T1_SOUTH_B1_valid_out),
		.S(RMUX_T1_SOUTH_B1_sel_value_O),
		.out_sel(RMUX_T1_SOUTH_B1_out_sel)
	);
	SliceWrapper_32_2_3 RMUX_T1_SOUTH_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T1_SOUTH_B1_sel_value_O)
	);
	wire [1:0] RMUX_T1_WEST_B1_I;
	assign RMUX_T1_WEST_B1_I[1+:1] = REG_T1_WEST_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T1_WEST_B1_I[0+:1] = MUX_SB_T1_WEST_SB_OUT_B1_O;
	wire [1:0] RMUX_T1_WEST_B1_valid_in;
	assign RMUX_T1_WEST_B1_valid_in = {REG_T1_WEST_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T1_WEST_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T1_WEST_B1(
		.I(RMUX_T1_WEST_B1_I),
		.O(RMUX_T1_WEST_B1_O),
		.ready_in(SB_T1_WEST_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T1_WEST_B1_ready_out),
		.valid_in(RMUX_T1_WEST_B1_valid_in),
		.valid_out(RMUX_T1_WEST_B1_valid_out),
		.S(RMUX_T1_WEST_B1_sel_value_O),
		.out_sel(RMUX_T1_WEST_B1_out_sel)
	);
	SliceWrapper_32_3_4 RMUX_T1_WEST_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T1_WEST_B1_sel_value_O)
	);
	wire [1:0] RMUX_T2_EAST_B1_I;
	assign RMUX_T2_EAST_B1_I[1+:1] = REG_T2_EAST_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T2_EAST_B1_I[0+:1] = MUX_SB_T2_EAST_SB_OUT_B1_O;
	wire [1:0] RMUX_T2_EAST_B1_valid_in;
	assign RMUX_T2_EAST_B1_valid_in = {REG_T2_EAST_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T2_EAST_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T2_EAST_B1(
		.I(RMUX_T2_EAST_B1_I),
		.O(RMUX_T2_EAST_B1_O),
		.ready_in(SB_T2_EAST_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T2_EAST_B1_ready_out),
		.valid_in(RMUX_T2_EAST_B1_valid_in),
		.valid_out(RMUX_T2_EAST_B1_valid_out),
		.S(RMUX_T2_EAST_B1_sel_value_O),
		.out_sel(RMUX_T2_EAST_B1_out_sel)
	);
	SliceWrapper_32_4_5 RMUX_T2_EAST_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T2_EAST_B1_sel_value_O)
	);
	wire [1:0] RMUX_T2_NORTH_B1_I;
	assign RMUX_T2_NORTH_B1_I[1+:1] = REG_T2_NORTH_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T2_NORTH_B1_I[0+:1] = MUX_SB_T2_NORTH_SB_OUT_B1_O;
	wire [1:0] RMUX_T2_NORTH_B1_valid_in;
	assign RMUX_T2_NORTH_B1_valid_in = {REG_T2_NORTH_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T2_NORTH_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T2_NORTH_B1(
		.I(RMUX_T2_NORTH_B1_I),
		.O(RMUX_T2_NORTH_B1_O),
		.ready_in(SB_T2_NORTH_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T2_NORTH_B1_ready_out),
		.valid_in(RMUX_T2_NORTH_B1_valid_in),
		.valid_out(RMUX_T2_NORTH_B1_valid_out),
		.S(RMUX_T2_NORTH_B1_sel_value_O),
		.out_sel(RMUX_T2_NORTH_B1_out_sel)
	);
	SliceWrapper_32_5_6 RMUX_T2_NORTH_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T2_NORTH_B1_sel_value_O)
	);
	wire [1:0] RMUX_T2_SOUTH_B1_I;
	assign RMUX_T2_SOUTH_B1_I[1+:1] = REG_T2_SOUTH_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T2_SOUTH_B1_I[0+:1] = MUX_SB_T2_SOUTH_SB_OUT_B1_O;
	wire [1:0] RMUX_T2_SOUTH_B1_valid_in;
	assign RMUX_T2_SOUTH_B1_valid_in = {REG_T2_SOUTH_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T2_SOUTH_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T2_SOUTH_B1(
		.I(RMUX_T2_SOUTH_B1_I),
		.O(RMUX_T2_SOUTH_B1_O),
		.ready_in(SB_T2_SOUTH_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T2_SOUTH_B1_ready_out),
		.valid_in(RMUX_T2_SOUTH_B1_valid_in),
		.valid_out(RMUX_T2_SOUTH_B1_valid_out),
		.S(RMUX_T2_SOUTH_B1_sel_value_O),
		.out_sel(RMUX_T2_SOUTH_B1_out_sel)
	);
	SliceWrapper_32_6_7 RMUX_T2_SOUTH_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T2_SOUTH_B1_sel_value_O)
	);
	wire [1:0] RMUX_T2_WEST_B1_I;
	assign RMUX_T2_WEST_B1_I[1+:1] = REG_T2_WEST_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T2_WEST_B1_I[0+:1] = MUX_SB_T2_WEST_SB_OUT_B1_O;
	wire [1:0] RMUX_T2_WEST_B1_valid_in;
	assign RMUX_T2_WEST_B1_valid_in = {REG_T2_WEST_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T2_WEST_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T2_WEST_B1(
		.I(RMUX_T2_WEST_B1_I),
		.O(RMUX_T2_WEST_B1_O),
		.ready_in(SB_T2_WEST_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T2_WEST_B1_ready_out),
		.valid_in(RMUX_T2_WEST_B1_valid_in),
		.valid_out(RMUX_T2_WEST_B1_valid_out),
		.S(RMUX_T2_WEST_B1_sel_value_O),
		.out_sel(RMUX_T2_WEST_B1_out_sel)
	);
	SliceWrapper_32_7_8 RMUX_T2_WEST_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T2_WEST_B1_sel_value_O)
	);
	wire [1:0] RMUX_T3_EAST_B1_I;
	assign RMUX_T3_EAST_B1_I[1+:1] = REG_T3_EAST_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T3_EAST_B1_I[0+:1] = MUX_SB_T3_EAST_SB_OUT_B1_O;
	wire [1:0] RMUX_T3_EAST_B1_valid_in;
	assign RMUX_T3_EAST_B1_valid_in = {REG_T3_EAST_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T3_EAST_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T3_EAST_B1(
		.I(RMUX_T3_EAST_B1_I),
		.O(RMUX_T3_EAST_B1_O),
		.ready_in(SB_T3_EAST_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T3_EAST_B1_ready_out),
		.valid_in(RMUX_T3_EAST_B1_valid_in),
		.valid_out(RMUX_T3_EAST_B1_valid_out),
		.S(RMUX_T3_EAST_B1_sel_value_O),
		.out_sel(RMUX_T3_EAST_B1_out_sel)
	);
	SliceWrapper_32_8_9 RMUX_T3_EAST_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T3_EAST_B1_sel_value_O)
	);
	wire [1:0] RMUX_T3_NORTH_B1_I;
	assign RMUX_T3_NORTH_B1_I[1+:1] = REG_T3_NORTH_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T3_NORTH_B1_I[0+:1] = MUX_SB_T3_NORTH_SB_OUT_B1_O;
	wire [1:0] RMUX_T3_NORTH_B1_valid_in;
	assign RMUX_T3_NORTH_B1_valid_in = {REG_T3_NORTH_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T3_NORTH_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T3_NORTH_B1(
		.I(RMUX_T3_NORTH_B1_I),
		.O(RMUX_T3_NORTH_B1_O),
		.ready_in(SB_T3_NORTH_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T3_NORTH_B1_ready_out),
		.valid_in(RMUX_T3_NORTH_B1_valid_in),
		.valid_out(RMUX_T3_NORTH_B1_valid_out),
		.S(RMUX_T3_NORTH_B1_sel_value_O),
		.out_sel(RMUX_T3_NORTH_B1_out_sel)
	);
	SliceWrapper_32_9_10 RMUX_T3_NORTH_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T3_NORTH_B1_sel_value_O)
	);
	wire [1:0] RMUX_T3_SOUTH_B1_I;
	assign RMUX_T3_SOUTH_B1_I[1+:1] = REG_T3_SOUTH_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T3_SOUTH_B1_I[0+:1] = MUX_SB_T3_SOUTH_SB_OUT_B1_O;
	wire [1:0] RMUX_T3_SOUTH_B1_valid_in;
	assign RMUX_T3_SOUTH_B1_valid_in = {REG_T3_SOUTH_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T3_SOUTH_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T3_SOUTH_B1(
		.I(RMUX_T3_SOUTH_B1_I),
		.O(RMUX_T3_SOUTH_B1_O),
		.ready_in(SB_T3_SOUTH_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T3_SOUTH_B1_ready_out),
		.valid_in(RMUX_T3_SOUTH_B1_valid_in),
		.valid_out(RMUX_T3_SOUTH_B1_valid_out),
		.S(RMUX_T3_SOUTH_B1_sel_value_O),
		.out_sel(RMUX_T3_SOUTH_B1_out_sel)
	);
	SliceWrapper_32_10_11 RMUX_T3_SOUTH_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T3_SOUTH_B1_sel_value_O)
	);
	wire [1:0] RMUX_T3_WEST_B1_I;
	assign RMUX_T3_WEST_B1_I[1+:1] = REG_T3_WEST_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T3_WEST_B1_I[0+:1] = MUX_SB_T3_WEST_SB_OUT_B1_O;
	wire [1:0] RMUX_T3_WEST_B1_valid_in;
	assign RMUX_T3_WEST_B1_valid_in = {REG_T3_WEST_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T3_WEST_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T3_WEST_B1(
		.I(RMUX_T3_WEST_B1_I),
		.O(RMUX_T3_WEST_B1_O),
		.ready_in(SB_T3_WEST_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T3_WEST_B1_ready_out),
		.valid_in(RMUX_T3_WEST_B1_valid_in),
		.valid_out(RMUX_T3_WEST_B1_valid_out),
		.S(RMUX_T3_WEST_B1_sel_value_O),
		.out_sel(RMUX_T3_WEST_B1_out_sel)
	);
	SliceWrapper_32_11_12 RMUX_T3_WEST_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T3_WEST_B1_sel_value_O)
	);
	wire [1:0] RMUX_T4_EAST_B1_I;
	assign RMUX_T4_EAST_B1_I[1+:1] = REG_T4_EAST_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T4_EAST_B1_I[0+:1] = MUX_SB_T4_EAST_SB_OUT_B1_O;
	wire [1:0] RMUX_T4_EAST_B1_valid_in;
	assign RMUX_T4_EAST_B1_valid_in = {REG_T4_EAST_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T4_EAST_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T4_EAST_B1(
		.I(RMUX_T4_EAST_B1_I),
		.O(RMUX_T4_EAST_B1_O),
		.ready_in(SB_T4_EAST_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T4_EAST_B1_ready_out),
		.valid_in(RMUX_T4_EAST_B1_valid_in),
		.valid_out(RMUX_T4_EAST_B1_valid_out),
		.S(RMUX_T4_EAST_B1_sel_value_O),
		.out_sel(RMUX_T4_EAST_B1_out_sel)
	);
	SliceWrapper_32_12_13 RMUX_T4_EAST_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T4_EAST_B1_sel_value_O)
	);
	wire [1:0] RMUX_T4_NORTH_B1_I;
	assign RMUX_T4_NORTH_B1_I[1+:1] = REG_T4_NORTH_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T4_NORTH_B1_I[0+:1] = MUX_SB_T4_NORTH_SB_OUT_B1_O;
	wire [1:0] RMUX_T4_NORTH_B1_valid_in;
	assign RMUX_T4_NORTH_B1_valid_in = {REG_T4_NORTH_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T4_NORTH_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T4_NORTH_B1(
		.I(RMUX_T4_NORTH_B1_I),
		.O(RMUX_T4_NORTH_B1_O),
		.ready_in(SB_T4_NORTH_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T4_NORTH_B1_ready_out),
		.valid_in(RMUX_T4_NORTH_B1_valid_in),
		.valid_out(RMUX_T4_NORTH_B1_valid_out),
		.S(RMUX_T4_NORTH_B1_sel_value_O),
		.out_sel(RMUX_T4_NORTH_B1_out_sel)
	);
	SliceWrapper_32_13_14 RMUX_T4_NORTH_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T4_NORTH_B1_sel_value_O)
	);
	wire [1:0] RMUX_T4_SOUTH_B1_I;
	assign RMUX_T4_SOUTH_B1_I[1+:1] = REG_T4_SOUTH_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T4_SOUTH_B1_I[0+:1] = MUX_SB_T4_SOUTH_SB_OUT_B1_O;
	wire [1:0] RMUX_T4_SOUTH_B1_valid_in;
	assign RMUX_T4_SOUTH_B1_valid_in = {REG_T4_SOUTH_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T4_SOUTH_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T4_SOUTH_B1(
		.I(RMUX_T4_SOUTH_B1_I),
		.O(RMUX_T4_SOUTH_B1_O),
		.ready_in(SB_T4_SOUTH_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T4_SOUTH_B1_ready_out),
		.valid_in(RMUX_T4_SOUTH_B1_valid_in),
		.valid_out(RMUX_T4_SOUTH_B1_valid_out),
		.S(RMUX_T4_SOUTH_B1_sel_value_O),
		.out_sel(RMUX_T4_SOUTH_B1_out_sel)
	);
	SliceWrapper_32_14_15 RMUX_T4_SOUTH_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T4_SOUTH_B1_sel_value_O)
	);
	wire [1:0] RMUX_T4_WEST_B1_I;
	assign RMUX_T4_WEST_B1_I[1+:1] = REG_T4_WEST_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T4_WEST_B1_I[0+:1] = MUX_SB_T4_WEST_SB_OUT_B1_O;
	wire [1:0] RMUX_T4_WEST_B1_valid_in;
	assign RMUX_T4_WEST_B1_valid_in = {REG_T4_WEST_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T4_WEST_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T4_WEST_B1(
		.I(RMUX_T4_WEST_B1_I),
		.O(RMUX_T4_WEST_B1_O),
		.ready_in(SB_T4_WEST_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T4_WEST_B1_ready_out),
		.valid_in(RMUX_T4_WEST_B1_valid_in),
		.valid_out(RMUX_T4_WEST_B1_valid_out),
		.S(RMUX_T4_WEST_B1_sel_value_O),
		.out_sel(RMUX_T4_WEST_B1_out_sel)
	);
	SliceWrapper_32_15_16 RMUX_T4_WEST_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T4_WEST_B1_sel_value_O)
	);
	SliceWrapper_32_16_17 SB_T0_EAST_SB_IN_B1_enable_value(
		.I(config_reg_2_O),
		.O(SB_T0_EAST_SB_IN_B1_enable_value_O)
	);
	FanoutHash_302974B49BE3F0C4 SB_T0_EAST_SB_IN_B1_fan_in(
		.E6(const_0_1_out),
		.E3(PE_input_width_1_num_0_enable),
		.I5(PE_input_width_1_num_2_ready),
		.S6(const_0_32_out),
		.E0(SB_T0_WEST_SB_OUT_B1_enable_value_O),
		.S5(PE_input_width_1_num_2_out_sel),
		.I6(const_0_1_out),
		.S3(PE_input_width_1_num_0_out_sel),
		.S4(PE_input_width_1_num_1_out_sel),
		.I3(PE_input_width_1_num_0_ready),
		.I4(PE_input_width_1_num_1_ready),
		.S1(MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T0_WEST_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T4_NORTH_SB_OUT_B1_out_sel),
		.E2(SB_T4_NORTH_SB_OUT_B1_enable_value_O),
		.E5(PE_input_width_1_num_2_enable),
		.E4(PE_input_width_1_num_1_enable),
		.I2(MUX_SB_T4_NORTH_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out),
		.O(SB_T0_EAST_SB_IN_B1_fan_in_O),
		.E1(SB_T3_SOUTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T0_WEST_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T0_EAST_SB_OUT_B1_FANOUT_I;
	assign SB_T0_EAST_SB_OUT_B1_FANOUT_I = {REG_T0_EAST_B1$SplitFifo_1_inst0_ready0[0], RMUX_T0_EAST_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T0_EAST_SB_OUT_B1_FANOUT(
		.O(SB_T0_EAST_SB_OUT_B1_FANOUT_O),
		.I(SB_T0_EAST_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T0_EAST_B1_out_sel)
	);
	SliceWrapper_32_17_18 SB_T0_EAST_SB_OUT_B1_enable_value(
		.I(config_reg_2_O),
		.O(SB_T0_EAST_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_32_18_21 SB_T0_EAST_SB_OUT_B1_sel_value(
		.I(config_reg_2_O),
		.O(SB_T0_EAST_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_32_21_22 SB_T0_NORTH_SB_IN_B1_enable_value(
		.I(config_reg_2_O),
		.O(SB_T0_NORTH_SB_IN_B1_enable_value_O)
	);
	FanoutHash_47712AAC902ADA2 SB_T0_NORTH_SB_IN_B1_fan_in(
		.E6(const_0_1_out),
		.E3(PE_input_width_1_num_0_enable),
		.I5(PE_input_width_1_num_2_ready),
		.S6(const_0_32_out),
		.E0(SB_T0_WEST_SB_OUT_B1_enable_value_O),
		.S5(PE_input_width_1_num_2_out_sel),
		.I6(const_0_1_out),
		.S3(PE_input_width_1_num_0_out_sel),
		.S4(PE_input_width_1_num_1_out_sel),
		.I3(PE_input_width_1_num_0_ready),
		.I4(PE_input_width_1_num_1_ready),
		.S1(MUX_SB_T1_EAST_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T0_WEST_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel),
		.E2(SB_T0_SOUTH_SB_OUT_B1_enable_value_O),
		.E5(PE_input_width_1_num_2_enable),
		.E4(PE_input_width_1_num_1_enable),
		.I2(MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T1_EAST_SB_OUT_B1_ready_out),
		.O(SB_T0_NORTH_SB_IN_B1_fan_in_O),
		.E1(SB_T1_EAST_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T0_WEST_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T0_NORTH_SB_OUT_B1_FANOUT_I;
	assign SB_T0_NORTH_SB_OUT_B1_FANOUT_I = {REG_T0_NORTH_B1$SplitFifo_1_inst0_ready0[0], RMUX_T0_NORTH_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T0_NORTH_SB_OUT_B1_FANOUT(
		.O(SB_T0_NORTH_SB_OUT_B1_FANOUT_O),
		.I(SB_T0_NORTH_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T0_NORTH_B1_out_sel)
	);
	SliceWrapper_32_22_23 SB_T0_NORTH_SB_OUT_B1_enable_value(
		.I(config_reg_2_O),
		.O(SB_T0_NORTH_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_32_23_26 SB_T0_NORTH_SB_OUT_B1_sel_value(
		.I(config_reg_2_O),
		.O(SB_T0_NORTH_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_32_26_27 SB_T0_SOUTH_SB_IN_B1_enable_value(
		.I(config_reg_2_O),
		.O(SB_T0_SOUTH_SB_IN_B1_enable_value_O)
	);
	FanoutHash_2785CE916183C5C SB_T0_SOUTH_SB_IN_B1_fan_in(
		.E6(const_0_1_out),
		.E3(PE_input_width_1_num_0_enable),
		.I5(PE_input_width_1_num_2_ready),
		.S6(const_0_32_out),
		.E0(SB_T3_EAST_SB_OUT_B1_enable_value_O),
		.S5(PE_input_width_1_num_2_out_sel),
		.I6(const_0_1_out),
		.S3(PE_input_width_1_num_0_out_sel),
		.S4(PE_input_width_1_num_1_out_sel),
		.I3(PE_input_width_1_num_0_ready),
		.I4(PE_input_width_1_num_1_ready),
		.S1(MUX_SB_T0_NORTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T3_EAST_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T1_WEST_SB_OUT_B1_out_sel),
		.E2(SB_T1_WEST_SB_OUT_B1_enable_value_O),
		.E5(PE_input_width_1_num_2_enable),
		.E4(PE_input_width_1_num_1_enable),
		.I2(MUX_SB_T1_WEST_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T0_NORTH_SB_OUT_B1_ready_out),
		.O(SB_T0_SOUTH_SB_IN_B1_fan_in_O),
		.E1(SB_T0_NORTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T3_EAST_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T0_SOUTH_SB_OUT_B1_FANOUT_I;
	assign SB_T0_SOUTH_SB_OUT_B1_FANOUT_I = {REG_T0_SOUTH_B1$SplitFifo_1_inst0_ready0[0], RMUX_T0_SOUTH_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T0_SOUTH_SB_OUT_B1_FANOUT(
		.O(SB_T0_SOUTH_SB_OUT_B1_FANOUT_O),
		.I(SB_T0_SOUTH_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T0_SOUTH_B1_out_sel)
	);
	SliceWrapper_32_27_28 SB_T0_SOUTH_SB_OUT_B1_enable_value(
		.I(config_reg_2_O),
		.O(SB_T0_SOUTH_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_32_28_31 SB_T0_SOUTH_SB_OUT_B1_sel_value(
		.I(config_reg_2_O),
		.O(SB_T0_SOUTH_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_32_31_32 SB_T0_WEST_SB_IN_B1_enable_value(
		.I(config_reg_2_O),
		.O(SB_T0_WEST_SB_IN_B1_enable_value_O)
	);
	FanoutHash_65A468071775C7BB SB_T0_WEST_SB_IN_B1_fan_in(
		.E6(const_0_1_out),
		.E3(PE_input_width_1_num_0_enable),
		.I5(PE_input_width_1_num_2_ready),
		.S6(const_0_32_out),
		.E0(SB_T0_NORTH_SB_OUT_B1_enable_value_O),
		.S5(PE_input_width_1_num_2_out_sel),
		.I6(const_0_1_out),
		.S3(PE_input_width_1_num_0_out_sel),
		.S4(PE_input_width_1_num_1_out_sel),
		.I3(PE_input_width_1_num_0_ready),
		.I4(PE_input_width_1_num_1_ready),
		.S1(MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T0_NORTH_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T0_EAST_SB_OUT_B1_out_sel),
		.E2(SB_T0_EAST_SB_OUT_B1_enable_value_O),
		.E5(PE_input_width_1_num_2_enable),
		.E4(PE_input_width_1_num_1_enable),
		.I2(MUX_SB_T0_EAST_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out),
		.O(SB_T0_WEST_SB_IN_B1_fan_in_O),
		.E1(SB_T4_SOUTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T0_NORTH_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T0_WEST_SB_OUT_B1_FANOUT_I;
	assign SB_T0_WEST_SB_OUT_B1_FANOUT_I = {REG_T0_WEST_B1$SplitFifo_1_inst0_ready0[0], RMUX_T0_WEST_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T0_WEST_SB_OUT_B1_FANOUT(
		.O(SB_T0_WEST_SB_OUT_B1_FANOUT_O),
		.I(SB_T0_WEST_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T0_WEST_B1_out_sel)
	);
	SliceWrapper_31_0_1 SB_T0_WEST_SB_OUT_B1_enable_value(
		.I(config_reg_3_O),
		.O(SB_T0_WEST_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_31_1_4 SB_T0_WEST_SB_OUT_B1_sel_value(
		.I(config_reg_3_O),
		.O(SB_T0_WEST_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_31_4_5 SB_T1_EAST_SB_IN_B1_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_EAST_SB_IN_B1_enable_value_O)
	);
	FanoutHash_4F83851A40824F89 SB_T1_EAST_SB_IN_B1_fan_in(
		.E6(const_0_1_out),
		.E3(PE_input_width_1_num_0_enable),
		.I5(PE_input_width_1_num_2_ready),
		.S6(const_0_32_out),
		.E0(SB_T0_NORTH_SB_OUT_B1_enable_value_O),
		.S5(PE_input_width_1_num_2_out_sel),
		.I6(const_0_1_out),
		.S3(PE_input_width_1_num_0_out_sel),
		.S4(PE_input_width_1_num_1_out_sel),
		.I3(PE_input_width_1_num_0_ready),
		.I4(PE_input_width_1_num_1_ready),
		.S1(MUX_SB_T1_WEST_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T0_NORTH_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel),
		.E2(SB_T2_SOUTH_SB_OUT_B1_enable_value_O),
		.E5(PE_input_width_1_num_2_enable),
		.E4(PE_input_width_1_num_1_enable),
		.I2(MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T1_WEST_SB_OUT_B1_ready_out),
		.O(SB_T1_EAST_SB_IN_B1_fan_in_O),
		.E1(SB_T1_WEST_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T0_NORTH_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T1_EAST_SB_OUT_B1_FANOUT_I;
	assign SB_T1_EAST_SB_OUT_B1_FANOUT_I = {REG_T1_EAST_B1$SplitFifo_1_inst0_ready0[0], RMUX_T1_EAST_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T1_EAST_SB_OUT_B1_FANOUT(
		.O(SB_T1_EAST_SB_OUT_B1_FANOUT_O),
		.I(SB_T1_EAST_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T1_EAST_B1_out_sel)
	);
	SliceWrapper_31_5_6 SB_T1_EAST_SB_OUT_B1_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_EAST_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_31_6_9 SB_T1_EAST_SB_OUT_B1_sel_value(
		.I(config_reg_3_O),
		.O(SB_T1_EAST_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_31_9_10 SB_T1_NORTH_SB_IN_B1_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_NORTH_SB_IN_B1_enable_value_O)
	);
	FanoutHash_4FADDC8F90390680 SB_T1_NORTH_SB_IN_B1_fan_in(
		.E6(const_0_1_out),
		.E3(PE_input_width_1_num_0_enable),
		.I5(PE_input_width_1_num_2_ready),
		.S6(const_0_32_out),
		.E0(SB_T2_EAST_SB_OUT_B1_enable_value_O),
		.S5(PE_input_width_1_num_2_out_sel),
		.I6(const_0_1_out),
		.S3(PE_input_width_1_num_0_out_sel),
		.S4(PE_input_width_1_num_1_out_sel),
		.I3(PE_input_width_1_num_0_ready),
		.I4(PE_input_width_1_num_1_ready),
		.S1(MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T2_EAST_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T4_WEST_SB_OUT_B1_out_sel),
		.E2(SB_T4_WEST_SB_OUT_B1_enable_value_O),
		.E5(PE_input_width_1_num_2_enable),
		.E4(PE_input_width_1_num_1_enable),
		.I2(MUX_SB_T4_WEST_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out),
		.O(SB_T1_NORTH_SB_IN_B1_fan_in_O),
		.E1(SB_T1_SOUTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T2_EAST_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T1_NORTH_SB_OUT_B1_FANOUT_I;
	assign SB_T1_NORTH_SB_OUT_B1_FANOUT_I = {REG_T1_NORTH_B1$SplitFifo_1_inst0_ready0[0], RMUX_T1_NORTH_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T1_NORTH_SB_OUT_B1_FANOUT(
		.O(SB_T1_NORTH_SB_OUT_B1_FANOUT_O),
		.I(SB_T1_NORTH_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T1_NORTH_B1_out_sel)
	);
	SliceWrapper_31_10_11 SB_T1_NORTH_SB_OUT_B1_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_NORTH_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_31_11_14 SB_T1_NORTH_SB_OUT_B1_sel_value(
		.I(config_reg_3_O),
		.O(SB_T1_NORTH_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_31_14_15 SB_T1_SOUTH_SB_IN_B1_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_SOUTH_SB_IN_B1_enable_value_O)
	);
	FanoutHash_466EB88CFD0CAD7B SB_T1_SOUTH_SB_IN_B1_fan_in(
		.E6(const_0_1_out),
		.E3(PE_input_width_1_num_0_enable),
		.I5(PE_input_width_1_num_2_ready),
		.S6(const_0_32_out),
		.E0(SB_T2_EAST_SB_OUT_B1_enable_value_O),
		.S5(PE_input_width_1_num_2_out_sel),
		.I6(const_0_1_out),
		.S3(PE_input_width_1_num_0_out_sel),
		.S4(PE_input_width_1_num_1_out_sel),
		.I3(PE_input_width_1_num_0_ready),
		.I4(PE_input_width_1_num_1_ready),
		.S1(MUX_SB_T1_NORTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T2_EAST_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T2_WEST_SB_OUT_B1_out_sel),
		.E2(SB_T2_WEST_SB_OUT_B1_enable_value_O),
		.E5(PE_input_width_1_num_2_enable),
		.E4(PE_input_width_1_num_1_enable),
		.I2(MUX_SB_T2_WEST_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T1_NORTH_SB_OUT_B1_ready_out),
		.O(SB_T1_SOUTH_SB_IN_B1_fan_in_O),
		.E1(SB_T1_NORTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T2_EAST_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T1_SOUTH_SB_OUT_B1_FANOUT_I;
	assign SB_T1_SOUTH_SB_OUT_B1_FANOUT_I = {REG_T1_SOUTH_B1$SplitFifo_1_inst0_ready0[0], RMUX_T1_SOUTH_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T1_SOUTH_SB_OUT_B1_FANOUT(
		.O(SB_T1_SOUTH_SB_OUT_B1_FANOUT_O),
		.I(SB_T1_SOUTH_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T1_SOUTH_B1_out_sel)
	);
	SliceWrapper_31_15_16 SB_T1_SOUTH_SB_OUT_B1_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_SOUTH_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_31_16_19 SB_T1_SOUTH_SB_OUT_B1_sel_value(
		.I(config_reg_3_O),
		.O(SB_T1_SOUTH_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_31_19_20 SB_T1_WEST_SB_IN_B1_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_WEST_SB_IN_B1_enable_value_O)
	);
	FanoutHash_7ED1C80229B84786 SB_T1_WEST_SB_IN_B1_fan_in(
		.E6(const_0_1_out),
		.E3(PE_input_width_1_num_0_enable),
		.I5(PE_input_width_1_num_2_ready),
		.S6(const_0_32_out),
		.E0(SB_T4_NORTH_SB_OUT_B1_enable_value_O),
		.S5(PE_input_width_1_num_2_out_sel),
		.I6(const_0_1_out),
		.S3(PE_input_width_1_num_0_out_sel),
		.S4(PE_input_width_1_num_1_out_sel),
		.I3(PE_input_width_1_num_0_ready),
		.I4(PE_input_width_1_num_1_ready),
		.S1(MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T4_NORTH_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T1_EAST_SB_OUT_B1_out_sel),
		.E2(SB_T1_EAST_SB_OUT_B1_enable_value_O),
		.E5(PE_input_width_1_num_2_enable),
		.E4(PE_input_width_1_num_1_enable),
		.I2(MUX_SB_T1_EAST_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out),
		.O(SB_T1_WEST_SB_IN_B1_fan_in_O),
		.E1(SB_T0_SOUTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T4_NORTH_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T1_WEST_SB_OUT_B1_FANOUT_I;
	assign SB_T1_WEST_SB_OUT_B1_FANOUT_I = {REG_T1_WEST_B1$SplitFifo_1_inst0_ready0[0], RMUX_T1_WEST_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T1_WEST_SB_OUT_B1_FANOUT(
		.O(SB_T1_WEST_SB_OUT_B1_FANOUT_O),
		.I(SB_T1_WEST_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T1_WEST_B1_out_sel)
	);
	SliceWrapper_31_20_21 SB_T1_WEST_SB_OUT_B1_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_WEST_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_31_21_24 SB_T1_WEST_SB_OUT_B1_sel_value(
		.I(config_reg_3_O),
		.O(SB_T1_WEST_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_31_24_25 SB_T2_EAST_SB_IN_B1_enable_value(
		.I(config_reg_3_O),
		.O(SB_T2_EAST_SB_IN_B1_enable_value_O)
	);
	FanoutHash_7F4660D1463D9234 SB_T2_EAST_SB_IN_B1_fan_in(
		.E6(const_0_1_out),
		.E3(PE_input_width_1_num_0_enable),
		.I5(PE_input_width_1_num_2_ready),
		.S6(const_0_32_out),
		.E0(SB_T1_NORTH_SB_OUT_B1_enable_value_O),
		.S5(PE_input_width_1_num_2_out_sel),
		.I6(const_0_1_out),
		.S3(PE_input_width_1_num_0_out_sel),
		.S4(PE_input_width_1_num_1_out_sel),
		.I3(PE_input_width_1_num_0_ready),
		.I4(PE_input_width_1_num_1_ready),
		.S1(MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T1_NORTH_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T2_WEST_SB_OUT_B1_out_sel),
		.E2(SB_T2_WEST_SB_OUT_B1_enable_value_O),
		.E5(PE_input_width_1_num_2_enable),
		.E4(PE_input_width_1_num_1_enable),
		.I2(MUX_SB_T2_WEST_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out),
		.O(SB_T2_EAST_SB_IN_B1_fan_in_O),
		.E1(SB_T1_SOUTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T1_NORTH_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T2_EAST_SB_OUT_B1_FANOUT_I;
	assign SB_T2_EAST_SB_OUT_B1_FANOUT_I = {REG_T2_EAST_B1$SplitFifo_1_inst0_ready0[0], RMUX_T2_EAST_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T2_EAST_SB_OUT_B1_FANOUT(
		.O(SB_T2_EAST_SB_OUT_B1_FANOUT_O),
		.I(SB_T2_EAST_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T2_EAST_B1_out_sel)
	);
	SliceWrapper_31_25_26 SB_T2_EAST_SB_OUT_B1_enable_value(
		.I(config_reg_3_O),
		.O(SB_T2_EAST_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_31_26_29 SB_T2_EAST_SB_OUT_B1_sel_value(
		.I(config_reg_3_O),
		.O(SB_T2_EAST_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_31_29_30 SB_T2_NORTH_SB_IN_B1_enable_value(
		.I(config_reg_3_O),
		.O(SB_T2_NORTH_SB_IN_B1_enable_value_O)
	);
	FanoutHash_3B67229CB02928BA SB_T2_NORTH_SB_IN_B1_fan_in(
		.E6(const_0_1_out),
		.E3(PE_input_width_1_num_0_enable),
		.I5(PE_input_width_1_num_2_ready),
		.S6(const_0_32_out),
		.E0(SB_T3_EAST_SB_OUT_B1_enable_value_O),
		.S5(PE_input_width_1_num_2_out_sel),
		.I6(const_0_1_out),
		.S3(PE_input_width_1_num_0_out_sel),
		.S4(PE_input_width_1_num_1_out_sel),
		.I3(PE_input_width_1_num_0_ready),
		.I4(PE_input_width_1_num_1_ready),
		.S1(MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T3_EAST_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T3_WEST_SB_OUT_B1_out_sel),
		.E2(SB_T3_WEST_SB_OUT_B1_enable_value_O),
		.E5(PE_input_width_1_num_2_enable),
		.E4(PE_input_width_1_num_1_enable),
		.I2(MUX_SB_T3_WEST_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out),
		.O(SB_T2_NORTH_SB_IN_B1_fan_in_O),
		.E1(SB_T2_SOUTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T3_EAST_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T2_NORTH_SB_OUT_B1_FANOUT_I;
	assign SB_T2_NORTH_SB_OUT_B1_FANOUT_I = {REG_T2_NORTH_B1$SplitFifo_1_inst0_ready0[0], RMUX_T2_NORTH_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T2_NORTH_SB_OUT_B1_FANOUT(
		.O(SB_T2_NORTH_SB_OUT_B1_FANOUT_O),
		.I(SB_T2_NORTH_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T2_NORTH_B1_out_sel)
	);
	SliceWrapper_31_30_31 SB_T2_NORTH_SB_OUT_B1_enable_value(
		.I(config_reg_3_O),
		.O(SB_T2_NORTH_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_30_0_3 SB_T2_NORTH_SB_OUT_B1_sel_value(
		.I(config_reg_4_O),
		.O(SB_T2_NORTH_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_30_3_4 SB_T2_SOUTH_SB_IN_B1_enable_value(
		.I(config_reg_4_O),
		.O(SB_T2_SOUTH_SB_IN_B1_enable_value_O)
	);
	FanoutHash_28125A548B305607 SB_T2_SOUTH_SB_IN_B1_fan_in(
		.E6(const_0_1_out),
		.E3(PE_input_width_1_num_0_enable),
		.I5(PE_input_width_1_num_2_ready),
		.S6(const_0_32_out),
		.E0(SB_T1_EAST_SB_OUT_B1_enable_value_O),
		.S5(PE_input_width_1_num_2_out_sel),
		.I6(const_0_1_out),
		.S3(PE_input_width_1_num_0_out_sel),
		.S4(PE_input_width_1_num_1_out_sel),
		.I3(PE_input_width_1_num_0_ready),
		.I4(PE_input_width_1_num_1_ready),
		.S1(MUX_SB_T2_NORTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T1_EAST_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T3_WEST_SB_OUT_B1_out_sel),
		.E2(SB_T3_WEST_SB_OUT_B1_enable_value_O),
		.E5(PE_input_width_1_num_2_enable),
		.E4(PE_input_width_1_num_1_enable),
		.I2(MUX_SB_T3_WEST_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T2_NORTH_SB_OUT_B1_ready_out),
		.O(SB_T2_SOUTH_SB_IN_B1_fan_in_O),
		.E1(SB_T2_NORTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T1_EAST_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T2_SOUTH_SB_OUT_B1_FANOUT_I;
	assign SB_T2_SOUTH_SB_OUT_B1_FANOUT_I = {REG_T2_SOUTH_B1$SplitFifo_1_inst0_ready0[0], RMUX_T2_SOUTH_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T2_SOUTH_SB_OUT_B1_FANOUT(
		.O(SB_T2_SOUTH_SB_OUT_B1_FANOUT_O),
		.I(SB_T2_SOUTH_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T2_SOUTH_B1_out_sel)
	);
	SliceWrapper_30_4_5 SB_T2_SOUTH_SB_OUT_B1_enable_value(
		.I(config_reg_4_O),
		.O(SB_T2_SOUTH_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_30_5_8 SB_T2_SOUTH_SB_OUT_B1_sel_value(
		.I(config_reg_4_O),
		.O(SB_T2_SOUTH_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_30_8_9 SB_T2_WEST_SB_IN_B1_enable_value(
		.I(config_reg_4_O),
		.O(SB_T2_WEST_SB_IN_B1_enable_value_O)
	);
	FanoutHash_752C11B748DD905C SB_T2_WEST_SB_IN_B1_fan_in(
		.E6(const_0_1_out),
		.E3(PE_input_width_1_num_0_enable),
		.I5(PE_input_width_1_num_2_ready),
		.S6(const_0_32_out),
		.E0(SB_T3_NORTH_SB_OUT_B1_enable_value_O),
		.S5(PE_input_width_1_num_2_out_sel),
		.I6(const_0_1_out),
		.S3(PE_input_width_1_num_0_out_sel),
		.S4(PE_input_width_1_num_1_out_sel),
		.I3(PE_input_width_1_num_0_ready),
		.I4(PE_input_width_1_num_1_ready),
		.S1(MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T3_NORTH_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T2_EAST_SB_OUT_B1_out_sel),
		.E2(SB_T2_EAST_SB_OUT_B1_enable_value_O),
		.E5(PE_input_width_1_num_2_enable),
		.E4(PE_input_width_1_num_1_enable),
		.I2(MUX_SB_T2_EAST_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out),
		.O(SB_T2_WEST_SB_IN_B1_fan_in_O),
		.E1(SB_T1_SOUTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T3_NORTH_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T2_WEST_SB_OUT_B1_FANOUT_I;
	assign SB_T2_WEST_SB_OUT_B1_FANOUT_I = {REG_T2_WEST_B1$SplitFifo_1_inst0_ready0[0], RMUX_T2_WEST_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T2_WEST_SB_OUT_B1_FANOUT(
		.O(SB_T2_WEST_SB_OUT_B1_FANOUT_O),
		.I(SB_T2_WEST_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T2_WEST_B1_out_sel)
	);
	SliceWrapper_30_9_10 SB_T2_WEST_SB_OUT_B1_enable_value(
		.I(config_reg_4_O),
		.O(SB_T2_WEST_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_30_10_13 SB_T2_WEST_SB_OUT_B1_sel_value(
		.I(config_reg_4_O),
		.O(SB_T2_WEST_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_30_13_14 SB_T3_EAST_SB_IN_B1_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_EAST_SB_IN_B1_enable_value_O)
	);
	FanoutHash_43D5C80ABD816837 SB_T3_EAST_SB_IN_B1_fan_in(
		.E6(const_0_1_out),
		.E3(PE_input_width_1_num_0_enable),
		.I5(PE_input_width_1_num_2_ready),
		.S6(const_0_32_out),
		.E0(SB_T0_SOUTH_SB_OUT_B1_enable_value_O),
		.S5(PE_input_width_1_num_2_out_sel),
		.I6(const_0_1_out),
		.S3(PE_input_width_1_num_0_out_sel),
		.S4(PE_input_width_1_num_1_out_sel),
		.I3(PE_input_width_1_num_0_ready),
		.I4(PE_input_width_1_num_1_ready),
		.S1(MUX_SB_T2_NORTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T3_WEST_SB_OUT_B1_out_sel),
		.E2(SB_T3_WEST_SB_OUT_B1_enable_value_O),
		.E5(PE_input_width_1_num_2_enable),
		.E4(PE_input_width_1_num_1_enable),
		.I2(MUX_SB_T3_WEST_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T2_NORTH_SB_OUT_B1_ready_out),
		.O(SB_T3_EAST_SB_IN_B1_fan_in_O),
		.E1(SB_T2_NORTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T3_EAST_SB_OUT_B1_FANOUT_I;
	assign SB_T3_EAST_SB_OUT_B1_FANOUT_I = {REG_T3_EAST_B1$SplitFifo_1_inst0_ready0[0], RMUX_T3_EAST_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T3_EAST_SB_OUT_B1_FANOUT(
		.O(SB_T3_EAST_SB_OUT_B1_FANOUT_O),
		.I(SB_T3_EAST_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T3_EAST_B1_out_sel)
	);
	SliceWrapper_30_14_15 SB_T3_EAST_SB_OUT_B1_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_EAST_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_30_15_18 SB_T3_EAST_SB_OUT_B1_sel_value(
		.I(config_reg_4_O),
		.O(SB_T3_EAST_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_30_18_19 SB_T3_NORTH_SB_IN_B1_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_NORTH_SB_IN_B1_enable_value_O)
	);
	FanoutHash_69376833A2418E2 SB_T3_NORTH_SB_IN_B1_fan_in(
		.E6(const_0_1_out),
		.E3(PE_input_width_1_num_0_enable),
		.I5(PE_input_width_1_num_2_ready),
		.S6(const_0_32_out),
		.E0(SB_T2_WEST_SB_OUT_B1_enable_value_O),
		.S5(PE_input_width_1_num_2_out_sel),
		.I6(const_0_1_out),
		.S3(PE_input_width_1_num_0_out_sel),
		.S4(PE_input_width_1_num_1_out_sel),
		.I3(PE_input_width_1_num_0_ready),
		.I4(PE_input_width_1_num_1_ready),
		.S1(MUX_SB_T4_EAST_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T2_WEST_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel),
		.E2(SB_T3_SOUTH_SB_OUT_B1_enable_value_O),
		.E5(PE_input_width_1_num_2_enable),
		.E4(PE_input_width_1_num_1_enable),
		.I2(MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T4_EAST_SB_OUT_B1_ready_out),
		.O(SB_T3_NORTH_SB_IN_B1_fan_in_O),
		.E1(SB_T4_EAST_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T2_WEST_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T3_NORTH_SB_OUT_B1_FANOUT_I;
	assign SB_T3_NORTH_SB_OUT_B1_FANOUT_I = {REG_T3_NORTH_B1$SplitFifo_1_inst0_ready0[0], RMUX_T3_NORTH_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T3_NORTH_SB_OUT_B1_FANOUT(
		.O(SB_T3_NORTH_SB_OUT_B1_FANOUT_O),
		.I(SB_T3_NORTH_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T3_NORTH_B1_out_sel)
	);
	SliceWrapper_30_19_20 SB_T3_NORTH_SB_OUT_B1_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_NORTH_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_30_20_23 SB_T3_NORTH_SB_OUT_B1_sel_value(
		.I(config_reg_4_O),
		.O(SB_T3_NORTH_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_30_23_24 SB_T3_SOUTH_SB_IN_B1_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_SOUTH_SB_IN_B1_enable_value_O)
	);
	FanoutHash_66A75CC8494A4D6B SB_T3_SOUTH_SB_IN_B1_fan_in(
		.E6(const_0_1_out),
		.E3(PE_input_width_1_num_0_enable),
		.I5(PE_input_width_1_num_2_ready),
		.S6(const_0_32_out),
		.E0(SB_T0_EAST_SB_OUT_B1_enable_value_O),
		.S5(PE_input_width_1_num_2_out_sel),
		.I6(const_0_1_out),
		.S3(PE_input_width_1_num_0_out_sel),
		.S4(PE_input_width_1_num_1_out_sel),
		.I3(PE_input_width_1_num_0_ready),
		.I4(PE_input_width_1_num_1_ready),
		.S1(MUX_SB_T3_NORTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T0_EAST_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T4_WEST_SB_OUT_B1_out_sel),
		.E2(SB_T4_WEST_SB_OUT_B1_enable_value_O),
		.E5(PE_input_width_1_num_2_enable),
		.E4(PE_input_width_1_num_1_enable),
		.I2(MUX_SB_T4_WEST_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T3_NORTH_SB_OUT_B1_ready_out),
		.O(SB_T3_SOUTH_SB_IN_B1_fan_in_O),
		.E1(SB_T3_NORTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T0_EAST_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T3_SOUTH_SB_OUT_B1_FANOUT_I;
	assign SB_T3_SOUTH_SB_OUT_B1_FANOUT_I = {REG_T3_SOUTH_B1$SplitFifo_1_inst0_ready0[0], RMUX_T3_SOUTH_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T3_SOUTH_SB_OUT_B1_FANOUT(
		.O(SB_T3_SOUTH_SB_OUT_B1_FANOUT_O),
		.I(SB_T3_SOUTH_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T3_SOUTH_B1_out_sel)
	);
	SliceWrapper_30_24_25 SB_T3_SOUTH_SB_OUT_B1_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_SOUTH_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_30_25_28 SB_T3_SOUTH_SB_OUT_B1_sel_value(
		.I(config_reg_4_O),
		.O(SB_T3_SOUTH_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_30_28_29 SB_T3_WEST_SB_IN_B1_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_WEST_SB_IN_B1_enable_value_O)
	);
	FanoutHash_31AE65CCDD94603 SB_T3_WEST_SB_IN_B1_fan_in(
		.E6(const_0_1_out),
		.E3(PE_input_width_1_num_0_enable),
		.I5(PE_input_width_1_num_2_ready),
		.S6(const_0_32_out),
		.E0(SB_T2_NORTH_SB_OUT_B1_enable_value_O),
		.S5(PE_input_width_1_num_2_out_sel),
		.I6(const_0_1_out),
		.S3(PE_input_width_1_num_0_out_sel),
		.S4(PE_input_width_1_num_1_out_sel),
		.I3(PE_input_width_1_num_0_ready),
		.I4(PE_input_width_1_num_1_ready),
		.S1(MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T2_NORTH_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T3_EAST_SB_OUT_B1_out_sel),
		.E2(SB_T3_EAST_SB_OUT_B1_enable_value_O),
		.E5(PE_input_width_1_num_2_enable),
		.E4(PE_input_width_1_num_1_enable),
		.I2(MUX_SB_T3_EAST_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out),
		.O(SB_T3_WEST_SB_IN_B1_fan_in_O),
		.E1(SB_T2_SOUTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T2_NORTH_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T3_WEST_SB_OUT_B1_FANOUT_I;
	assign SB_T3_WEST_SB_OUT_B1_FANOUT_I = {REG_T3_WEST_B1$SplitFifo_1_inst0_ready0[0], RMUX_T3_WEST_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T3_WEST_SB_OUT_B1_FANOUT(
		.O(SB_T3_WEST_SB_OUT_B1_FANOUT_O),
		.I(SB_T3_WEST_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T3_WEST_B1_out_sel)
	);
	SliceWrapper_30_29_30 SB_T3_WEST_SB_OUT_B1_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_WEST_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_23_0_3 SB_T3_WEST_SB_OUT_B1_sel_value(
		.I(config_reg_5_O),
		.O(SB_T3_WEST_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_23_3_4 SB_T4_EAST_SB_IN_B1_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_EAST_SB_IN_B1_enable_value_O)
	);
	FanoutHash_5D7AEC1255CDC1CC SB_T4_EAST_SB_IN_B1_fan_in(
		.E6(const_0_1_out),
		.E3(PE_input_width_1_num_0_enable),
		.I5(PE_input_width_1_num_2_ready),
		.S6(const_0_32_out),
		.E0(SB_T3_NORTH_SB_OUT_B1_enable_value_O),
		.S5(PE_input_width_1_num_2_out_sel),
		.I6(const_0_1_out),
		.S3(PE_input_width_1_num_0_out_sel),
		.S4(PE_input_width_1_num_1_out_sel),
		.I3(PE_input_width_1_num_0_ready),
		.I4(PE_input_width_1_num_1_ready),
		.S1(MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T3_NORTH_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T4_WEST_SB_OUT_B1_out_sel),
		.E2(SB_T4_WEST_SB_OUT_B1_enable_value_O),
		.E5(PE_input_width_1_num_2_enable),
		.E4(PE_input_width_1_num_1_enable),
		.I2(MUX_SB_T4_WEST_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out),
		.O(SB_T4_EAST_SB_IN_B1_fan_in_O),
		.E1(SB_T4_SOUTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T3_NORTH_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T4_EAST_SB_OUT_B1_FANOUT_I;
	assign SB_T4_EAST_SB_OUT_B1_FANOUT_I = {REG_T4_EAST_B1$SplitFifo_1_inst0_ready0[0], RMUX_T4_EAST_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T4_EAST_SB_OUT_B1_FANOUT(
		.O(SB_T4_EAST_SB_OUT_B1_FANOUT_O),
		.I(SB_T4_EAST_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T4_EAST_B1_out_sel)
	);
	SliceWrapper_23_4_5 SB_T4_EAST_SB_OUT_B1_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_EAST_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_23_5_8 SB_T4_EAST_SB_OUT_B1_sel_value(
		.I(config_reg_5_O),
		.O(SB_T4_EAST_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_23_8_9 SB_T4_NORTH_SB_IN_B1_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_NORTH_SB_IN_B1_enable_value_O)
	);
	FanoutHash_184DFC10DAF19BE9 SB_T4_NORTH_SB_IN_B1_fan_in(
		.E6(const_0_1_out),
		.E3(PE_input_width_1_num_0_enable),
		.I5(PE_input_width_1_num_2_ready),
		.S6(const_0_32_out),
		.E0(SB_T1_WEST_SB_OUT_B1_enable_value_O),
		.S5(PE_input_width_1_num_2_out_sel),
		.I6(const_0_1_out),
		.S3(PE_input_width_1_num_0_out_sel),
		.S4(PE_input_width_1_num_1_out_sel),
		.I3(PE_input_width_1_num_0_ready),
		.I4(PE_input_width_1_num_1_ready),
		.S1(MUX_SB_T0_EAST_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T1_WEST_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel),
		.E2(SB_T4_SOUTH_SB_OUT_B1_enable_value_O),
		.E5(PE_input_width_1_num_2_enable),
		.E4(PE_input_width_1_num_1_enable),
		.I2(MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T0_EAST_SB_OUT_B1_ready_out),
		.O(SB_T4_NORTH_SB_IN_B1_fan_in_O),
		.E1(SB_T0_EAST_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T1_WEST_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T4_NORTH_SB_OUT_B1_FANOUT_I;
	assign SB_T4_NORTH_SB_OUT_B1_FANOUT_I = {REG_T4_NORTH_B1$SplitFifo_1_inst0_ready0[0], RMUX_T4_NORTH_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T4_NORTH_SB_OUT_B1_FANOUT(
		.O(SB_T4_NORTH_SB_OUT_B1_FANOUT_O),
		.I(SB_T4_NORTH_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T4_NORTH_B1_out_sel)
	);
	SliceWrapper_23_9_10 SB_T4_NORTH_SB_OUT_B1_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_NORTH_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_23_10_13 SB_T4_NORTH_SB_OUT_B1_sel_value(
		.I(config_reg_5_O),
		.O(SB_T4_NORTH_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_23_13_14 SB_T4_SOUTH_SB_IN_B1_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_SOUTH_SB_IN_B1_enable_value_O)
	);
	FanoutHash_26B6474864379B6A SB_T4_SOUTH_SB_IN_B1_fan_in(
		.E6(const_0_1_out),
		.E3(PE_input_width_1_num_0_enable),
		.I5(PE_input_width_1_num_2_ready),
		.S6(const_0_32_out),
		.E0(SB_T0_WEST_SB_OUT_B1_enable_value_O),
		.S5(PE_input_width_1_num_2_out_sel),
		.I6(const_0_1_out),
		.S3(PE_input_width_1_num_0_out_sel),
		.S4(PE_input_width_1_num_1_out_sel),
		.I3(PE_input_width_1_num_0_ready),
		.I4(PE_input_width_1_num_1_ready),
		.S1(MUX_SB_T4_EAST_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T0_WEST_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T4_NORTH_SB_OUT_B1_out_sel),
		.E2(SB_T4_NORTH_SB_OUT_B1_enable_value_O),
		.E5(PE_input_width_1_num_2_enable),
		.E4(PE_input_width_1_num_1_enable),
		.I2(MUX_SB_T4_NORTH_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T4_EAST_SB_OUT_B1_ready_out),
		.O(SB_T4_SOUTH_SB_IN_B1_fan_in_O),
		.E1(SB_T4_EAST_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T0_WEST_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T4_SOUTH_SB_OUT_B1_FANOUT_I;
	assign SB_T4_SOUTH_SB_OUT_B1_FANOUT_I = {REG_T4_SOUTH_B1$SplitFifo_1_inst0_ready0[0], RMUX_T4_SOUTH_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T4_SOUTH_SB_OUT_B1_FANOUT(
		.O(SB_T4_SOUTH_SB_OUT_B1_FANOUT_O),
		.I(SB_T4_SOUTH_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T4_SOUTH_B1_out_sel)
	);
	SliceWrapper_23_14_15 SB_T4_SOUTH_SB_OUT_B1_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_SOUTH_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_23_15_18 SB_T4_SOUTH_SB_OUT_B1_sel_value(
		.I(config_reg_5_O),
		.O(SB_T4_SOUTH_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_23_18_19 SB_T4_WEST_SB_IN_B1_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_WEST_SB_IN_B1_enable_value_O)
	);
	FanoutHash_1816466D6957000 SB_T4_WEST_SB_IN_B1_fan_in(
		.E6(const_0_1_out),
		.E3(PE_input_width_1_num_0_enable),
		.I5(PE_input_width_1_num_2_ready),
		.S6(const_0_32_out),
		.E0(SB_T1_NORTH_SB_OUT_B1_enable_value_O),
		.S5(PE_input_width_1_num_2_out_sel),
		.I6(const_0_1_out),
		.S3(PE_input_width_1_num_0_out_sel),
		.S4(PE_input_width_1_num_1_out_sel),
		.I3(PE_input_width_1_num_0_ready),
		.I4(PE_input_width_1_num_1_ready),
		.S1(MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T1_NORTH_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T4_EAST_SB_OUT_B1_out_sel),
		.E2(SB_T4_EAST_SB_OUT_B1_enable_value_O),
		.E5(PE_input_width_1_num_2_enable),
		.E4(PE_input_width_1_num_1_enable),
		.I2(MUX_SB_T4_EAST_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out),
		.O(SB_T4_WEST_SB_IN_B1_fan_in_O),
		.E1(SB_T3_SOUTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T1_NORTH_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T4_WEST_SB_OUT_B1_FANOUT_I;
	assign SB_T4_WEST_SB_OUT_B1_FANOUT_I = {REG_T4_WEST_B1$SplitFifo_1_inst0_ready0[0], RMUX_T4_WEST_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T4_WEST_SB_OUT_B1_FANOUT(
		.O(SB_T4_WEST_SB_OUT_B1_FANOUT_O),
		.I(SB_T4_WEST_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T4_WEST_B1_out_sel)
	);
	SliceWrapper_23_19_20 SB_T4_WEST_SB_OUT_B1_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_WEST_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_23_20_23 SB_T4_WEST_SB_OUT_B1_sel_value(
		.I(config_reg_5_O),
		.O(SB_T4_WEST_SB_OUT_B1_sel_value_O)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T0_EAST_SB_IN_B1(
		.I(SB_T0_EAST_SB_IN_B1),
		.O(WIRE_SB_T0_EAST_SB_IN_B1_O),
		.ready_in(SB_T0_EAST_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T0_EAST_SB_IN_B1_ready_out),
		.valid_in(SB_T0_EAST_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T0_EAST_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T0_NORTH_SB_IN_B1(
		.I(SB_T0_NORTH_SB_IN_B1),
		.O(WIRE_SB_T0_NORTH_SB_IN_B1_O),
		.ready_in(SB_T0_NORTH_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T0_NORTH_SB_IN_B1_ready_out),
		.valid_in(SB_T0_NORTH_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T0_NORTH_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T0_SOUTH_SB_IN_B1(
		.I(SB_T0_SOUTH_SB_IN_B1),
		.O(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
		.ready_in(SB_T0_SOUTH_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T0_SOUTH_SB_IN_B1_ready_out),
		.valid_in(SB_T0_SOUTH_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T0_SOUTH_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T0_WEST_SB_IN_B1(
		.I(SB_T0_WEST_SB_IN_B1),
		.O(WIRE_SB_T0_WEST_SB_IN_B1_O),
		.ready_in(SB_T0_WEST_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T0_WEST_SB_IN_B1_ready_out),
		.valid_in(SB_T0_WEST_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T0_WEST_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T1_EAST_SB_IN_B1(
		.I(SB_T1_EAST_SB_IN_B1),
		.O(WIRE_SB_T1_EAST_SB_IN_B1_O),
		.ready_in(SB_T1_EAST_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T1_EAST_SB_IN_B1_ready_out),
		.valid_in(SB_T1_EAST_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T1_EAST_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T1_NORTH_SB_IN_B1(
		.I(SB_T1_NORTH_SB_IN_B1),
		.O(WIRE_SB_T1_NORTH_SB_IN_B1_O),
		.ready_in(SB_T1_NORTH_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T1_NORTH_SB_IN_B1_ready_out),
		.valid_in(SB_T1_NORTH_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T1_NORTH_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T1_SOUTH_SB_IN_B1(
		.I(SB_T1_SOUTH_SB_IN_B1),
		.O(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
		.ready_in(SB_T1_SOUTH_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T1_SOUTH_SB_IN_B1_ready_out),
		.valid_in(SB_T1_SOUTH_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T1_SOUTH_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T1_WEST_SB_IN_B1(
		.I(SB_T1_WEST_SB_IN_B1),
		.O(WIRE_SB_T1_WEST_SB_IN_B1_O),
		.ready_in(SB_T1_WEST_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T1_WEST_SB_IN_B1_ready_out),
		.valid_in(SB_T1_WEST_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T1_WEST_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T2_EAST_SB_IN_B1(
		.I(SB_T2_EAST_SB_IN_B1),
		.O(WIRE_SB_T2_EAST_SB_IN_B1_O),
		.ready_in(SB_T2_EAST_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T2_EAST_SB_IN_B1_ready_out),
		.valid_in(SB_T2_EAST_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T2_EAST_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T2_NORTH_SB_IN_B1(
		.I(SB_T2_NORTH_SB_IN_B1),
		.O(WIRE_SB_T2_NORTH_SB_IN_B1_O),
		.ready_in(SB_T2_NORTH_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T2_NORTH_SB_IN_B1_ready_out),
		.valid_in(SB_T2_NORTH_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T2_NORTH_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T2_SOUTH_SB_IN_B1(
		.I(SB_T2_SOUTH_SB_IN_B1),
		.O(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
		.ready_in(SB_T2_SOUTH_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T2_SOUTH_SB_IN_B1_ready_out),
		.valid_in(SB_T2_SOUTH_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T2_SOUTH_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T2_WEST_SB_IN_B1(
		.I(SB_T2_WEST_SB_IN_B1),
		.O(WIRE_SB_T2_WEST_SB_IN_B1_O),
		.ready_in(SB_T2_WEST_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T2_WEST_SB_IN_B1_ready_out),
		.valid_in(SB_T2_WEST_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T2_WEST_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T3_EAST_SB_IN_B1(
		.I(SB_T3_EAST_SB_IN_B1),
		.O(WIRE_SB_T3_EAST_SB_IN_B1_O),
		.ready_in(SB_T3_EAST_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T3_EAST_SB_IN_B1_ready_out),
		.valid_in(SB_T3_EAST_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T3_EAST_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T3_NORTH_SB_IN_B1(
		.I(SB_T3_NORTH_SB_IN_B1),
		.O(WIRE_SB_T3_NORTH_SB_IN_B1_O),
		.ready_in(SB_T3_NORTH_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T3_NORTH_SB_IN_B1_ready_out),
		.valid_in(SB_T3_NORTH_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T3_NORTH_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T3_SOUTH_SB_IN_B1(
		.I(SB_T3_SOUTH_SB_IN_B1),
		.O(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
		.ready_in(SB_T3_SOUTH_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T3_SOUTH_SB_IN_B1_ready_out),
		.valid_in(SB_T3_SOUTH_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T3_SOUTH_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T3_WEST_SB_IN_B1(
		.I(SB_T3_WEST_SB_IN_B1),
		.O(WIRE_SB_T3_WEST_SB_IN_B1_O),
		.ready_in(SB_T3_WEST_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T3_WEST_SB_IN_B1_ready_out),
		.valid_in(SB_T3_WEST_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T3_WEST_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T4_EAST_SB_IN_B1(
		.I(SB_T4_EAST_SB_IN_B1),
		.O(WIRE_SB_T4_EAST_SB_IN_B1_O),
		.ready_in(SB_T4_EAST_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T4_EAST_SB_IN_B1_ready_out),
		.valid_in(SB_T4_EAST_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T4_EAST_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T4_NORTH_SB_IN_B1(
		.I(SB_T4_NORTH_SB_IN_B1),
		.O(WIRE_SB_T4_NORTH_SB_IN_B1_O),
		.ready_in(SB_T4_NORTH_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T4_NORTH_SB_IN_B1_ready_out),
		.valid_in(SB_T4_NORTH_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T4_NORTH_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T4_SOUTH_SB_IN_B1(
		.I(SB_T4_SOUTH_SB_IN_B1),
		.O(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
		.ready_in(SB_T4_SOUTH_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T4_SOUTH_SB_IN_B1_ready_out),
		.valid_in(SB_T4_SOUTH_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T4_SOUTH_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T4_WEST_SB_IN_B1(
		.I(SB_T4_WEST_SB_IN_B1),
		.O(WIRE_SB_T4_WEST_SB_IN_B1_O),
		.ready_in(SB_T4_WEST_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T4_WEST_SB_IN_B1_ready_out),
		.valid_in(SB_T4_WEST_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T4_WEST_SB_IN_B1_valid_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_23_32_inst0$bit_const_0_None(.out(ZextWrapper_23_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_23_32_inst0$self_O_out;
	assign ZextWrapper_23_32_inst0$self_O_out = {ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, config_reg_5_O};
	mantle_wire__typeBitIn32 ZextWrapper_23_32_inst0$self_O(
		.in(ZextWrapper_23_32_inst0$self_O_in),
		.out(ZextWrapper_23_32_inst0$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_30_32_inst0$bit_const_0_None(.out(ZextWrapper_30_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_30_32_inst0$self_O_out;
	assign ZextWrapper_30_32_inst0$self_O_out = {ZextWrapper_30_32_inst0$bit_const_0_None_out, ZextWrapper_30_32_inst0$bit_const_0_None_out, config_reg_4_O};
	mantle_wire__typeBitIn32 ZextWrapper_30_32_inst0$self_O(
		.in(ZextWrapper_30_32_inst0$self_O_in),
		.out(ZextWrapper_30_32_inst0$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_31_32_inst0$bit_const_0_None(.out(ZextWrapper_31_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_31_32_inst0$self_O_out;
	assign ZextWrapper_31_32_inst0$self_O_out = {ZextWrapper_31_32_inst0$bit_const_0_None_out, config_reg_3_O};
	mantle_wire__typeBitIn32 ZextWrapper_31_32_inst0$self_O(
		.in(ZextWrapper_31_32_inst0$self_O_in),
		.out(ZextWrapper_31_32_inst0$self_O_out)
	);
	coreir_and #(.width(1)) and1_inst0(
		.in0(coreir_eq_1_inst0_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst0_out)
	);
	coreir_and #(.width(1)) and1_inst1(
		.in0(coreir_eq_1_inst1_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst1_out)
	);
	coreir_and #(.width(1)) and1_inst10(
		.in0(coreir_eq_1_inst10_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst10_out)
	);
	coreir_and #(.width(1)) and1_inst11(
		.in0(coreir_eq_1_inst11_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst11_out)
	);
	coreir_and #(.width(1)) and1_inst12(
		.in0(coreir_eq_1_inst12_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst12_out)
	);
	coreir_and #(.width(1)) and1_inst13(
		.in0(coreir_eq_1_inst13_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst13_out)
	);
	coreir_and #(.width(1)) and1_inst14(
		.in0(coreir_eq_1_inst14_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst14_out)
	);
	coreir_and #(.width(1)) and1_inst15(
		.in0(coreir_eq_1_inst15_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst15_out)
	);
	coreir_and #(.width(1)) and1_inst16(
		.in0(coreir_eq_1_inst16_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst16_out)
	);
	coreir_and #(.width(1)) and1_inst17(
		.in0(coreir_eq_1_inst17_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst17_out)
	);
	coreir_and #(.width(1)) and1_inst18(
		.in0(coreir_eq_1_inst18_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst18_out)
	);
	coreir_and #(.width(1)) and1_inst19(
		.in0(coreir_eq_1_inst19_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst19_out)
	);
	coreir_and #(.width(1)) and1_inst2(
		.in0(coreir_eq_1_inst2_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst2_out)
	);
	coreir_and #(.width(1)) and1_inst3(
		.in0(coreir_eq_1_inst3_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst3_out)
	);
	coreir_and #(.width(1)) and1_inst4(
		.in0(coreir_eq_1_inst4_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst4_out)
	);
	coreir_and #(.width(1)) and1_inst5(
		.in0(coreir_eq_1_inst5_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst5_out)
	);
	coreir_and #(.width(1)) and1_inst6(
		.in0(coreir_eq_1_inst6_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst6_out)
	);
	coreir_and #(.width(1)) and1_inst7(
		.in0(coreir_eq_1_inst7_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst7_out)
	);
	coreir_and #(.width(1)) and1_inst8(
		.in0(coreir_eq_1_inst8_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst8_out)
	);
	coreir_and #(.width(1)) and1_inst9(
		.in0(coreir_eq_1_inst9_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst9_out)
	);
	wire [7:0] config_reg_0_config_addr;
	assign config_reg_0_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4], self_config_config_addr_out[3], self_config_config_addr_out[2:0]};
	ConfigRegister_32_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_reg_0_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_1_config_addr;
	assign config_reg_1_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4], self_config_config_addr_out[3], self_config_config_addr_out[2:0]};
	ConfigRegister_32_8_32_1 config_reg_1(
		.clk(clk),
		.reset(reset),
		.O(config_reg_1_O),
		.config_addr(config_reg_1_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_2_config_addr;
	assign config_reg_2_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4], self_config_config_addr_out[3], self_config_config_addr_out[2:0]};
	ConfigRegister_32_8_32_2 config_reg_2(
		.clk(clk),
		.reset(reset),
		.O(config_reg_2_O),
		.config_addr(config_reg_2_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_3_config_addr;
	assign config_reg_3_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4], self_config_config_addr_out[3], self_config_config_addr_out[2:0]};
	ConfigRegister_31_8_32_3 config_reg_3(
		.clk(clk),
		.reset(reset),
		.O(config_reg_3_O),
		.config_addr(config_reg_3_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_4_config_addr;
	assign config_reg_4_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4], self_config_config_addr_out[3], self_config_config_addr_out[2:0]};
	ConfigRegister_30_8_32_4 config_reg_4(
		.clk(clk),
		.reset(reset),
		.O(config_reg_4_O),
		.config_addr(config_reg_4_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_5_config_addr;
	assign config_reg_5_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4], self_config_config_addr_out[3], self_config_config_addr_out[2:0]};
	ConfigRegister_23_8_32_5 config_reg_5(
		.clk(clk),
		.reset(reset),
		.O(config_reg_5_O),
		.config_addr(config_reg_5_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	coreir_const #(
		.value(1'h0),
		.width(1)
	) const_0_1(.out(const_0_1_out));
	coreir_const #(
		.value(32'h00000000),
		.width(32)
	) const_0_32(.out(const_0_32_out));
	coreir_const #(
		.value(1'h1),
		.width(1)
	) const_1_1(.out(const_1_1_out));
	coreir_eq #(.width(1)) coreir_eq_1_inst0(
		.in0(const_1_1_out),
		.in1(RMUX_T0_NORTH_B1_sel_value_O),
		.out(coreir_eq_1_inst0_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst1(
		.in0(const_1_1_out),
		.in1(RMUX_T0_SOUTH_B1_sel_value_O),
		.out(coreir_eq_1_inst1_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst10(
		.in0(const_1_1_out),
		.in1(RMUX_T2_EAST_B1_sel_value_O),
		.out(coreir_eq_1_inst10_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst11(
		.in0(const_1_1_out),
		.in1(RMUX_T2_WEST_B1_sel_value_O),
		.out(coreir_eq_1_inst11_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst12(
		.in0(const_1_1_out),
		.in1(RMUX_T3_NORTH_B1_sel_value_O),
		.out(coreir_eq_1_inst12_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst13(
		.in0(const_1_1_out),
		.in1(RMUX_T3_SOUTH_B1_sel_value_O),
		.out(coreir_eq_1_inst13_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst14(
		.in0(const_1_1_out),
		.in1(RMUX_T3_EAST_B1_sel_value_O),
		.out(coreir_eq_1_inst14_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst15(
		.in0(const_1_1_out),
		.in1(RMUX_T3_WEST_B1_sel_value_O),
		.out(coreir_eq_1_inst15_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst16(
		.in0(const_1_1_out),
		.in1(RMUX_T4_NORTH_B1_sel_value_O),
		.out(coreir_eq_1_inst16_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst17(
		.in0(const_1_1_out),
		.in1(RMUX_T4_SOUTH_B1_sel_value_O),
		.out(coreir_eq_1_inst17_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst18(
		.in0(const_1_1_out),
		.in1(RMUX_T4_EAST_B1_sel_value_O),
		.out(coreir_eq_1_inst18_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst19(
		.in0(const_1_1_out),
		.in1(RMUX_T4_WEST_B1_sel_value_O),
		.out(coreir_eq_1_inst19_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst2(
		.in0(const_1_1_out),
		.in1(RMUX_T0_EAST_B1_sel_value_O),
		.out(coreir_eq_1_inst2_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst3(
		.in0(const_1_1_out),
		.in1(RMUX_T0_WEST_B1_sel_value_O),
		.out(coreir_eq_1_inst3_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst4(
		.in0(const_1_1_out),
		.in1(RMUX_T1_NORTH_B1_sel_value_O),
		.out(coreir_eq_1_inst4_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst5(
		.in0(const_1_1_out),
		.in1(RMUX_T1_SOUTH_B1_sel_value_O),
		.out(coreir_eq_1_inst5_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst6(
		.in0(const_1_1_out),
		.in1(RMUX_T1_EAST_B1_sel_value_O),
		.out(coreir_eq_1_inst6_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst7(
		.in0(const_1_1_out),
		.in1(RMUX_T1_WEST_B1_sel_value_O),
		.out(coreir_eq_1_inst7_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst8(
		.in0(const_1_1_out),
		.in1(RMUX_T2_NORTH_B1_sel_value_O),
		.out(coreir_eq_1_inst8_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst9(
		.in0(const_1_1_out),
		.in1(RMUX_T2_SOUTH_B1_sel_value_O),
		.out(coreir_eq_1_inst9_out)
	);
	wire [191:0] mux_aoi_6_32_inst0_I;
	assign mux_aoi_6_32_inst0_I[160+:32] = ZextWrapper_23_32_inst0$self_O_in;
	assign mux_aoi_6_32_inst0_I[128+:32] = ZextWrapper_30_32_inst0$self_O_in;
	assign mux_aoi_6_32_inst0_I[96+:32] = ZextWrapper_31_32_inst0$self_O_in;
	assign mux_aoi_6_32_inst0_I[64+:32] = config_reg_2_O;
	assign mux_aoi_6_32_inst0_I[32+:32] = config_reg_1_O;
	assign mux_aoi_6_32_inst0_I[0+:32] = config_reg_0_O;
	mux_aoi_6_32 mux_aoi_6_32_inst0(
		.I(mux_aoi_6_32_inst0_I),
		.O(mux_aoi_6_32_inst0_O),
		.S(self_config_config_addr_out[2:0]),
		.out_sel(mux_aoi_6_32_inst0_out_sel)
	);
	mantle_wire__typeBit8 self_config_config_addr(
		.in(config_config_addr),
		.out(self_config_config_addr_out)
	);
	assign PE_output_width_1_num_0_ready_out = CB_PE_output_width_1_num_0_fan_in_O[0];
	assign PondTop_output_width_1_num_0_ready_out = CB_PondTop_output_width_1_num_0_fan_in_O[0];
	assign PondTop_output_width_1_num_1_ready_out = CB_PondTop_output_width_1_num_1_fan_in_O[0];
	assign SB_T0_EAST_SB_IN_B1_enable = SB_T0_EAST_SB_IN_B1_enable_value_O[0];
	assign SB_T0_EAST_SB_IN_B1_ready_out = WIRE_SB_T0_EAST_SB_IN_B1_ready_out;
	assign SB_T0_EAST_SB_OUT_B1 = RMUX_T0_EAST_B1_O;
	assign SB_T0_EAST_SB_OUT_B1_enable = SB_T0_EAST_SB_OUT_B1_enable_value_O[0];
	assign SB_T0_EAST_SB_OUT_B1_valid_out = RMUX_T0_EAST_B1_valid_out;
	assign SB_T0_NORTH_SB_IN_B1_enable = SB_T0_NORTH_SB_IN_B1_enable_value_O[0];
	assign SB_T0_NORTH_SB_IN_B1_ready_out = WIRE_SB_T0_NORTH_SB_IN_B1_ready_out;
	assign SB_T0_NORTH_SB_OUT_B1 = RMUX_T0_NORTH_B1_O;
	assign SB_T0_NORTH_SB_OUT_B1_enable = SB_T0_NORTH_SB_OUT_B1_enable_value_O[0];
	assign SB_T0_NORTH_SB_OUT_B1_valid_out = RMUX_T0_NORTH_B1_valid_out;
	assign SB_T0_SOUTH_SB_IN_B1_enable = SB_T0_SOUTH_SB_IN_B1_enable_value_O[0];
	assign SB_T0_SOUTH_SB_IN_B1_ready_out = WIRE_SB_T0_SOUTH_SB_IN_B1_ready_out;
	assign SB_T0_SOUTH_SB_OUT_B1 = RMUX_T0_SOUTH_B1_O;
	assign SB_T0_SOUTH_SB_OUT_B1_enable = SB_T0_SOUTH_SB_OUT_B1_enable_value_O[0];
	assign SB_T0_SOUTH_SB_OUT_B1_valid_out = RMUX_T0_SOUTH_B1_valid_out;
	assign SB_T0_WEST_SB_IN_B1_enable = SB_T0_WEST_SB_IN_B1_enable_value_O[0];
	assign SB_T0_WEST_SB_IN_B1_ready_out = WIRE_SB_T0_WEST_SB_IN_B1_ready_out;
	assign SB_T0_WEST_SB_OUT_B1 = RMUX_T0_WEST_B1_O;
	assign SB_T0_WEST_SB_OUT_B1_enable = SB_T0_WEST_SB_OUT_B1_enable_value_O[0];
	assign SB_T0_WEST_SB_OUT_B1_valid_out = RMUX_T0_WEST_B1_valid_out;
	assign SB_T1_EAST_SB_IN_B1_enable = SB_T1_EAST_SB_IN_B1_enable_value_O[0];
	assign SB_T1_EAST_SB_IN_B1_ready_out = WIRE_SB_T1_EAST_SB_IN_B1_ready_out;
	assign SB_T1_EAST_SB_OUT_B1 = RMUX_T1_EAST_B1_O;
	assign SB_T1_EAST_SB_OUT_B1_enable = SB_T1_EAST_SB_OUT_B1_enable_value_O[0];
	assign SB_T1_EAST_SB_OUT_B1_valid_out = RMUX_T1_EAST_B1_valid_out;
	assign SB_T1_NORTH_SB_IN_B1_enable = SB_T1_NORTH_SB_IN_B1_enable_value_O[0];
	assign SB_T1_NORTH_SB_IN_B1_ready_out = WIRE_SB_T1_NORTH_SB_IN_B1_ready_out;
	assign SB_T1_NORTH_SB_OUT_B1 = RMUX_T1_NORTH_B1_O;
	assign SB_T1_NORTH_SB_OUT_B1_enable = SB_T1_NORTH_SB_OUT_B1_enable_value_O[0];
	assign SB_T1_NORTH_SB_OUT_B1_valid_out = RMUX_T1_NORTH_B1_valid_out;
	assign SB_T1_SOUTH_SB_IN_B1_enable = SB_T1_SOUTH_SB_IN_B1_enable_value_O[0];
	assign SB_T1_SOUTH_SB_IN_B1_ready_out = WIRE_SB_T1_SOUTH_SB_IN_B1_ready_out;
	assign SB_T1_SOUTH_SB_OUT_B1 = RMUX_T1_SOUTH_B1_O;
	assign SB_T1_SOUTH_SB_OUT_B1_enable = SB_T1_SOUTH_SB_OUT_B1_enable_value_O[0];
	assign SB_T1_SOUTH_SB_OUT_B1_valid_out = RMUX_T1_SOUTH_B1_valid_out;
	assign SB_T1_WEST_SB_IN_B1_enable = SB_T1_WEST_SB_IN_B1_enable_value_O[0];
	assign SB_T1_WEST_SB_IN_B1_ready_out = WIRE_SB_T1_WEST_SB_IN_B1_ready_out;
	assign SB_T1_WEST_SB_OUT_B1 = RMUX_T1_WEST_B1_O;
	assign SB_T1_WEST_SB_OUT_B1_enable = SB_T1_WEST_SB_OUT_B1_enable_value_O[0];
	assign SB_T1_WEST_SB_OUT_B1_valid_out = RMUX_T1_WEST_B1_valid_out;
	assign SB_T2_EAST_SB_IN_B1_enable = SB_T2_EAST_SB_IN_B1_enable_value_O[0];
	assign SB_T2_EAST_SB_IN_B1_ready_out = WIRE_SB_T2_EAST_SB_IN_B1_ready_out;
	assign SB_T2_EAST_SB_OUT_B1 = RMUX_T2_EAST_B1_O;
	assign SB_T2_EAST_SB_OUT_B1_enable = SB_T2_EAST_SB_OUT_B1_enable_value_O[0];
	assign SB_T2_EAST_SB_OUT_B1_valid_out = RMUX_T2_EAST_B1_valid_out;
	assign SB_T2_NORTH_SB_IN_B1_enable = SB_T2_NORTH_SB_IN_B1_enable_value_O[0];
	assign SB_T2_NORTH_SB_IN_B1_ready_out = WIRE_SB_T2_NORTH_SB_IN_B1_ready_out;
	assign SB_T2_NORTH_SB_OUT_B1 = RMUX_T2_NORTH_B1_O;
	assign SB_T2_NORTH_SB_OUT_B1_enable = SB_T2_NORTH_SB_OUT_B1_enable_value_O[0];
	assign SB_T2_NORTH_SB_OUT_B1_valid_out = RMUX_T2_NORTH_B1_valid_out;
	assign SB_T2_SOUTH_SB_IN_B1_enable = SB_T2_SOUTH_SB_IN_B1_enable_value_O[0];
	assign SB_T2_SOUTH_SB_IN_B1_ready_out = WIRE_SB_T2_SOUTH_SB_IN_B1_ready_out;
	assign SB_T2_SOUTH_SB_OUT_B1 = RMUX_T2_SOUTH_B1_O;
	assign SB_T2_SOUTH_SB_OUT_B1_enable = SB_T2_SOUTH_SB_OUT_B1_enable_value_O[0];
	assign SB_T2_SOUTH_SB_OUT_B1_valid_out = RMUX_T2_SOUTH_B1_valid_out;
	assign SB_T2_WEST_SB_IN_B1_enable = SB_T2_WEST_SB_IN_B1_enable_value_O[0];
	assign SB_T2_WEST_SB_IN_B1_ready_out = WIRE_SB_T2_WEST_SB_IN_B1_ready_out;
	assign SB_T2_WEST_SB_OUT_B1 = RMUX_T2_WEST_B1_O;
	assign SB_T2_WEST_SB_OUT_B1_enable = SB_T2_WEST_SB_OUT_B1_enable_value_O[0];
	assign SB_T2_WEST_SB_OUT_B1_valid_out = RMUX_T2_WEST_B1_valid_out;
	assign SB_T3_EAST_SB_IN_B1_enable = SB_T3_EAST_SB_IN_B1_enable_value_O[0];
	assign SB_T3_EAST_SB_IN_B1_ready_out = WIRE_SB_T3_EAST_SB_IN_B1_ready_out;
	assign SB_T3_EAST_SB_OUT_B1 = RMUX_T3_EAST_B1_O;
	assign SB_T3_EAST_SB_OUT_B1_enable = SB_T3_EAST_SB_OUT_B1_enable_value_O[0];
	assign SB_T3_EAST_SB_OUT_B1_valid_out = RMUX_T3_EAST_B1_valid_out;
	assign SB_T3_NORTH_SB_IN_B1_enable = SB_T3_NORTH_SB_IN_B1_enable_value_O[0];
	assign SB_T3_NORTH_SB_IN_B1_ready_out = WIRE_SB_T3_NORTH_SB_IN_B1_ready_out;
	assign SB_T3_NORTH_SB_OUT_B1 = RMUX_T3_NORTH_B1_O;
	assign SB_T3_NORTH_SB_OUT_B1_enable = SB_T3_NORTH_SB_OUT_B1_enable_value_O[0];
	assign SB_T3_NORTH_SB_OUT_B1_valid_out = RMUX_T3_NORTH_B1_valid_out;
	assign SB_T3_SOUTH_SB_IN_B1_enable = SB_T3_SOUTH_SB_IN_B1_enable_value_O[0];
	assign SB_T3_SOUTH_SB_IN_B1_ready_out = WIRE_SB_T3_SOUTH_SB_IN_B1_ready_out;
	assign SB_T3_SOUTH_SB_OUT_B1 = RMUX_T3_SOUTH_B1_O;
	assign SB_T3_SOUTH_SB_OUT_B1_enable = SB_T3_SOUTH_SB_OUT_B1_enable_value_O[0];
	assign SB_T3_SOUTH_SB_OUT_B1_valid_out = RMUX_T3_SOUTH_B1_valid_out;
	assign SB_T3_WEST_SB_IN_B1_enable = SB_T3_WEST_SB_IN_B1_enable_value_O[0];
	assign SB_T3_WEST_SB_IN_B1_ready_out = WIRE_SB_T3_WEST_SB_IN_B1_ready_out;
	assign SB_T3_WEST_SB_OUT_B1 = RMUX_T3_WEST_B1_O;
	assign SB_T3_WEST_SB_OUT_B1_enable = SB_T3_WEST_SB_OUT_B1_enable_value_O[0];
	assign SB_T3_WEST_SB_OUT_B1_valid_out = RMUX_T3_WEST_B1_valid_out;
	assign SB_T4_EAST_SB_IN_B1_enable = SB_T4_EAST_SB_IN_B1_enable_value_O[0];
	assign SB_T4_EAST_SB_IN_B1_ready_out = WIRE_SB_T4_EAST_SB_IN_B1_ready_out;
	assign SB_T4_EAST_SB_OUT_B1 = RMUX_T4_EAST_B1_O;
	assign SB_T4_EAST_SB_OUT_B1_enable = SB_T4_EAST_SB_OUT_B1_enable_value_O[0];
	assign SB_T4_EAST_SB_OUT_B1_valid_out = RMUX_T4_EAST_B1_valid_out;
	assign SB_T4_NORTH_SB_IN_B1_enable = SB_T4_NORTH_SB_IN_B1_enable_value_O[0];
	assign SB_T4_NORTH_SB_IN_B1_ready_out = WIRE_SB_T4_NORTH_SB_IN_B1_ready_out;
	assign SB_T4_NORTH_SB_OUT_B1 = RMUX_T4_NORTH_B1_O;
	assign SB_T4_NORTH_SB_OUT_B1_enable = SB_T4_NORTH_SB_OUT_B1_enable_value_O[0];
	assign SB_T4_NORTH_SB_OUT_B1_valid_out = RMUX_T4_NORTH_B1_valid_out;
	assign SB_T4_SOUTH_SB_IN_B1_enable = SB_T4_SOUTH_SB_IN_B1_enable_value_O[0];
	assign SB_T4_SOUTH_SB_IN_B1_ready_out = WIRE_SB_T4_SOUTH_SB_IN_B1_ready_out;
	assign SB_T4_SOUTH_SB_OUT_B1 = RMUX_T4_SOUTH_B1_O;
	assign SB_T4_SOUTH_SB_OUT_B1_enable = SB_T4_SOUTH_SB_OUT_B1_enable_value_O[0];
	assign SB_T4_SOUTH_SB_OUT_B1_valid_out = RMUX_T4_SOUTH_B1_valid_out;
	assign SB_T4_WEST_SB_IN_B1_enable = SB_T4_WEST_SB_IN_B1_enable_value_O[0];
	assign SB_T4_WEST_SB_IN_B1_ready_out = WIRE_SB_T4_WEST_SB_IN_B1_ready_out;
	assign SB_T4_WEST_SB_OUT_B1 = RMUX_T4_WEST_B1_O;
	assign SB_T4_WEST_SB_OUT_B1_enable = SB_T4_WEST_SB_OUT_B1_enable_value_O[0];
	assign SB_T4_WEST_SB_OUT_B1_valid_out = RMUX_T4_WEST_B1_valid_out;
	assign read_config_data = mux_aoi_6_32_inst0_O;
endmodule
module SB_ID0_5TRACKS_B1_MemCore (
	MEM_input_width_1_num_0_enable,
	MEM_input_width_1_num_0_out_sel,
	MEM_input_width_1_num_0_ready,
	MEM_input_width_1_num_1_enable,
	MEM_input_width_1_num_1_out_sel,
	MEM_input_width_1_num_1_ready,
	MEM_output_width_1_num_0,
	MEM_output_width_1_num_0_ready_out,
	MEM_output_width_1_num_0_valid,
	MEM_output_width_1_num_1,
	MEM_output_width_1_num_1_ready_out,
	MEM_output_width_1_num_1_valid,
	MEM_output_width_1_num_2,
	MEM_output_width_1_num_2_ready_out,
	MEM_output_width_1_num_2_valid,
	SB_T0_EAST_SB_IN_B1,
	SB_T0_EAST_SB_IN_B1_enable,
	SB_T0_EAST_SB_IN_B1_ready_out,
	SB_T0_EAST_SB_IN_B1_valid_in,
	SB_T0_EAST_SB_OUT_B1,
	SB_T0_EAST_SB_OUT_B1_enable,
	SB_T0_EAST_SB_OUT_B1_ready_in,
	SB_T0_EAST_SB_OUT_B1_valid_out,
	SB_T0_NORTH_SB_IN_B1,
	SB_T0_NORTH_SB_IN_B1_enable,
	SB_T0_NORTH_SB_IN_B1_ready_out,
	SB_T0_NORTH_SB_IN_B1_valid_in,
	SB_T0_NORTH_SB_OUT_B1,
	SB_T0_NORTH_SB_OUT_B1_enable,
	SB_T0_NORTH_SB_OUT_B1_ready_in,
	SB_T0_NORTH_SB_OUT_B1_valid_out,
	SB_T0_SOUTH_SB_IN_B1,
	SB_T0_SOUTH_SB_IN_B1_enable,
	SB_T0_SOUTH_SB_IN_B1_ready_out,
	SB_T0_SOUTH_SB_IN_B1_valid_in,
	SB_T0_SOUTH_SB_OUT_B1,
	SB_T0_SOUTH_SB_OUT_B1_enable,
	SB_T0_SOUTH_SB_OUT_B1_ready_in,
	SB_T0_SOUTH_SB_OUT_B1_valid_out,
	SB_T0_WEST_SB_IN_B1,
	SB_T0_WEST_SB_IN_B1_enable,
	SB_T0_WEST_SB_IN_B1_ready_out,
	SB_T0_WEST_SB_IN_B1_valid_in,
	SB_T0_WEST_SB_OUT_B1,
	SB_T0_WEST_SB_OUT_B1_enable,
	SB_T0_WEST_SB_OUT_B1_ready_in,
	SB_T0_WEST_SB_OUT_B1_valid_out,
	SB_T1_EAST_SB_IN_B1,
	SB_T1_EAST_SB_IN_B1_enable,
	SB_T1_EAST_SB_IN_B1_ready_out,
	SB_T1_EAST_SB_IN_B1_valid_in,
	SB_T1_EAST_SB_OUT_B1,
	SB_T1_EAST_SB_OUT_B1_enable,
	SB_T1_EAST_SB_OUT_B1_ready_in,
	SB_T1_EAST_SB_OUT_B1_valid_out,
	SB_T1_NORTH_SB_IN_B1,
	SB_T1_NORTH_SB_IN_B1_enable,
	SB_T1_NORTH_SB_IN_B1_ready_out,
	SB_T1_NORTH_SB_IN_B1_valid_in,
	SB_T1_NORTH_SB_OUT_B1,
	SB_T1_NORTH_SB_OUT_B1_enable,
	SB_T1_NORTH_SB_OUT_B1_ready_in,
	SB_T1_NORTH_SB_OUT_B1_valid_out,
	SB_T1_SOUTH_SB_IN_B1,
	SB_T1_SOUTH_SB_IN_B1_enable,
	SB_T1_SOUTH_SB_IN_B1_ready_out,
	SB_T1_SOUTH_SB_IN_B1_valid_in,
	SB_T1_SOUTH_SB_OUT_B1,
	SB_T1_SOUTH_SB_OUT_B1_enable,
	SB_T1_SOUTH_SB_OUT_B1_ready_in,
	SB_T1_SOUTH_SB_OUT_B1_valid_out,
	SB_T1_WEST_SB_IN_B1,
	SB_T1_WEST_SB_IN_B1_enable,
	SB_T1_WEST_SB_IN_B1_ready_out,
	SB_T1_WEST_SB_IN_B1_valid_in,
	SB_T1_WEST_SB_OUT_B1,
	SB_T1_WEST_SB_OUT_B1_enable,
	SB_T1_WEST_SB_OUT_B1_ready_in,
	SB_T1_WEST_SB_OUT_B1_valid_out,
	SB_T2_EAST_SB_IN_B1,
	SB_T2_EAST_SB_IN_B1_enable,
	SB_T2_EAST_SB_IN_B1_ready_out,
	SB_T2_EAST_SB_IN_B1_valid_in,
	SB_T2_EAST_SB_OUT_B1,
	SB_T2_EAST_SB_OUT_B1_enable,
	SB_T2_EAST_SB_OUT_B1_ready_in,
	SB_T2_EAST_SB_OUT_B1_valid_out,
	SB_T2_NORTH_SB_IN_B1,
	SB_T2_NORTH_SB_IN_B1_enable,
	SB_T2_NORTH_SB_IN_B1_ready_out,
	SB_T2_NORTH_SB_IN_B1_valid_in,
	SB_T2_NORTH_SB_OUT_B1,
	SB_T2_NORTH_SB_OUT_B1_enable,
	SB_T2_NORTH_SB_OUT_B1_ready_in,
	SB_T2_NORTH_SB_OUT_B1_valid_out,
	SB_T2_SOUTH_SB_IN_B1,
	SB_T2_SOUTH_SB_IN_B1_enable,
	SB_T2_SOUTH_SB_IN_B1_ready_out,
	SB_T2_SOUTH_SB_IN_B1_valid_in,
	SB_T2_SOUTH_SB_OUT_B1,
	SB_T2_SOUTH_SB_OUT_B1_enable,
	SB_T2_SOUTH_SB_OUT_B1_ready_in,
	SB_T2_SOUTH_SB_OUT_B1_valid_out,
	SB_T2_WEST_SB_IN_B1,
	SB_T2_WEST_SB_IN_B1_enable,
	SB_T2_WEST_SB_IN_B1_ready_out,
	SB_T2_WEST_SB_IN_B1_valid_in,
	SB_T2_WEST_SB_OUT_B1,
	SB_T2_WEST_SB_OUT_B1_enable,
	SB_T2_WEST_SB_OUT_B1_ready_in,
	SB_T2_WEST_SB_OUT_B1_valid_out,
	SB_T3_EAST_SB_IN_B1,
	SB_T3_EAST_SB_IN_B1_enable,
	SB_T3_EAST_SB_IN_B1_ready_out,
	SB_T3_EAST_SB_IN_B1_valid_in,
	SB_T3_EAST_SB_OUT_B1,
	SB_T3_EAST_SB_OUT_B1_enable,
	SB_T3_EAST_SB_OUT_B1_ready_in,
	SB_T3_EAST_SB_OUT_B1_valid_out,
	SB_T3_NORTH_SB_IN_B1,
	SB_T3_NORTH_SB_IN_B1_enable,
	SB_T3_NORTH_SB_IN_B1_ready_out,
	SB_T3_NORTH_SB_IN_B1_valid_in,
	SB_T3_NORTH_SB_OUT_B1,
	SB_T3_NORTH_SB_OUT_B1_enable,
	SB_T3_NORTH_SB_OUT_B1_ready_in,
	SB_T3_NORTH_SB_OUT_B1_valid_out,
	SB_T3_SOUTH_SB_IN_B1,
	SB_T3_SOUTH_SB_IN_B1_enable,
	SB_T3_SOUTH_SB_IN_B1_ready_out,
	SB_T3_SOUTH_SB_IN_B1_valid_in,
	SB_T3_SOUTH_SB_OUT_B1,
	SB_T3_SOUTH_SB_OUT_B1_enable,
	SB_T3_SOUTH_SB_OUT_B1_ready_in,
	SB_T3_SOUTH_SB_OUT_B1_valid_out,
	SB_T3_WEST_SB_IN_B1,
	SB_T3_WEST_SB_IN_B1_enable,
	SB_T3_WEST_SB_IN_B1_ready_out,
	SB_T3_WEST_SB_IN_B1_valid_in,
	SB_T3_WEST_SB_OUT_B1,
	SB_T3_WEST_SB_OUT_B1_enable,
	SB_T3_WEST_SB_OUT_B1_ready_in,
	SB_T3_WEST_SB_OUT_B1_valid_out,
	SB_T4_EAST_SB_IN_B1,
	SB_T4_EAST_SB_IN_B1_enable,
	SB_T4_EAST_SB_IN_B1_ready_out,
	SB_T4_EAST_SB_IN_B1_valid_in,
	SB_T4_EAST_SB_OUT_B1,
	SB_T4_EAST_SB_OUT_B1_enable,
	SB_T4_EAST_SB_OUT_B1_ready_in,
	SB_T4_EAST_SB_OUT_B1_valid_out,
	SB_T4_NORTH_SB_IN_B1,
	SB_T4_NORTH_SB_IN_B1_enable,
	SB_T4_NORTH_SB_IN_B1_ready_out,
	SB_T4_NORTH_SB_IN_B1_valid_in,
	SB_T4_NORTH_SB_OUT_B1,
	SB_T4_NORTH_SB_OUT_B1_enable,
	SB_T4_NORTH_SB_OUT_B1_ready_in,
	SB_T4_NORTH_SB_OUT_B1_valid_out,
	SB_T4_SOUTH_SB_IN_B1,
	SB_T4_SOUTH_SB_IN_B1_enable,
	SB_T4_SOUTH_SB_IN_B1_ready_out,
	SB_T4_SOUTH_SB_IN_B1_valid_in,
	SB_T4_SOUTH_SB_OUT_B1,
	SB_T4_SOUTH_SB_OUT_B1_enable,
	SB_T4_SOUTH_SB_OUT_B1_ready_in,
	SB_T4_SOUTH_SB_OUT_B1_valid_out,
	SB_T4_WEST_SB_IN_B1,
	SB_T4_WEST_SB_IN_B1_enable,
	SB_T4_WEST_SB_IN_B1_ready_out,
	SB_T4_WEST_SB_IN_B1_valid_in,
	SB_T4_WEST_SB_OUT_B1,
	SB_T4_WEST_SB_OUT_B1_enable,
	SB_T4_WEST_SB_OUT_B1_ready_in,
	SB_T4_WEST_SB_OUT_B1_valid_out,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	read_config_data,
	reset,
	stall
);
	input [0:0] MEM_input_width_1_num_0_enable;
	input [31:0] MEM_input_width_1_num_0_out_sel;
	input MEM_input_width_1_num_0_ready;
	input [0:0] MEM_input_width_1_num_1_enable;
	input [31:0] MEM_input_width_1_num_1_out_sel;
	input MEM_input_width_1_num_1_ready;
	input [0:0] MEM_output_width_1_num_0;
	output wire MEM_output_width_1_num_0_ready_out;
	input MEM_output_width_1_num_0_valid;
	input [0:0] MEM_output_width_1_num_1;
	output wire MEM_output_width_1_num_1_ready_out;
	input MEM_output_width_1_num_1_valid;
	input [0:0] MEM_output_width_1_num_2;
	output wire MEM_output_width_1_num_2_ready_out;
	input MEM_output_width_1_num_2_valid;
	input [0:0] SB_T0_EAST_SB_IN_B1;
	output wire SB_T0_EAST_SB_IN_B1_enable;
	output wire SB_T0_EAST_SB_IN_B1_ready_out;
	input SB_T0_EAST_SB_IN_B1_valid_in;
	output wire [0:0] SB_T0_EAST_SB_OUT_B1;
	output wire SB_T0_EAST_SB_OUT_B1_enable;
	input SB_T0_EAST_SB_OUT_B1_ready_in;
	output wire SB_T0_EAST_SB_OUT_B1_valid_out;
	input [0:0] SB_T0_NORTH_SB_IN_B1;
	output wire SB_T0_NORTH_SB_IN_B1_enable;
	output wire SB_T0_NORTH_SB_IN_B1_ready_out;
	input SB_T0_NORTH_SB_IN_B1_valid_in;
	output wire [0:0] SB_T0_NORTH_SB_OUT_B1;
	output wire SB_T0_NORTH_SB_OUT_B1_enable;
	input SB_T0_NORTH_SB_OUT_B1_ready_in;
	output wire SB_T0_NORTH_SB_OUT_B1_valid_out;
	input [0:0] SB_T0_SOUTH_SB_IN_B1;
	output wire SB_T0_SOUTH_SB_IN_B1_enable;
	output wire SB_T0_SOUTH_SB_IN_B1_ready_out;
	input SB_T0_SOUTH_SB_IN_B1_valid_in;
	output wire [0:0] SB_T0_SOUTH_SB_OUT_B1;
	output wire SB_T0_SOUTH_SB_OUT_B1_enable;
	input SB_T0_SOUTH_SB_OUT_B1_ready_in;
	output wire SB_T0_SOUTH_SB_OUT_B1_valid_out;
	input [0:0] SB_T0_WEST_SB_IN_B1;
	output wire SB_T0_WEST_SB_IN_B1_enable;
	output wire SB_T0_WEST_SB_IN_B1_ready_out;
	input SB_T0_WEST_SB_IN_B1_valid_in;
	output wire [0:0] SB_T0_WEST_SB_OUT_B1;
	output wire SB_T0_WEST_SB_OUT_B1_enable;
	input SB_T0_WEST_SB_OUT_B1_ready_in;
	output wire SB_T0_WEST_SB_OUT_B1_valid_out;
	input [0:0] SB_T1_EAST_SB_IN_B1;
	output wire SB_T1_EAST_SB_IN_B1_enable;
	output wire SB_T1_EAST_SB_IN_B1_ready_out;
	input SB_T1_EAST_SB_IN_B1_valid_in;
	output wire [0:0] SB_T1_EAST_SB_OUT_B1;
	output wire SB_T1_EAST_SB_OUT_B1_enable;
	input SB_T1_EAST_SB_OUT_B1_ready_in;
	output wire SB_T1_EAST_SB_OUT_B1_valid_out;
	input [0:0] SB_T1_NORTH_SB_IN_B1;
	output wire SB_T1_NORTH_SB_IN_B1_enable;
	output wire SB_T1_NORTH_SB_IN_B1_ready_out;
	input SB_T1_NORTH_SB_IN_B1_valid_in;
	output wire [0:0] SB_T1_NORTH_SB_OUT_B1;
	output wire SB_T1_NORTH_SB_OUT_B1_enable;
	input SB_T1_NORTH_SB_OUT_B1_ready_in;
	output wire SB_T1_NORTH_SB_OUT_B1_valid_out;
	input [0:0] SB_T1_SOUTH_SB_IN_B1;
	output wire SB_T1_SOUTH_SB_IN_B1_enable;
	output wire SB_T1_SOUTH_SB_IN_B1_ready_out;
	input SB_T1_SOUTH_SB_IN_B1_valid_in;
	output wire [0:0] SB_T1_SOUTH_SB_OUT_B1;
	output wire SB_T1_SOUTH_SB_OUT_B1_enable;
	input SB_T1_SOUTH_SB_OUT_B1_ready_in;
	output wire SB_T1_SOUTH_SB_OUT_B1_valid_out;
	input [0:0] SB_T1_WEST_SB_IN_B1;
	output wire SB_T1_WEST_SB_IN_B1_enable;
	output wire SB_T1_WEST_SB_IN_B1_ready_out;
	input SB_T1_WEST_SB_IN_B1_valid_in;
	output wire [0:0] SB_T1_WEST_SB_OUT_B1;
	output wire SB_T1_WEST_SB_OUT_B1_enable;
	input SB_T1_WEST_SB_OUT_B1_ready_in;
	output wire SB_T1_WEST_SB_OUT_B1_valid_out;
	input [0:0] SB_T2_EAST_SB_IN_B1;
	output wire SB_T2_EAST_SB_IN_B1_enable;
	output wire SB_T2_EAST_SB_IN_B1_ready_out;
	input SB_T2_EAST_SB_IN_B1_valid_in;
	output wire [0:0] SB_T2_EAST_SB_OUT_B1;
	output wire SB_T2_EAST_SB_OUT_B1_enable;
	input SB_T2_EAST_SB_OUT_B1_ready_in;
	output wire SB_T2_EAST_SB_OUT_B1_valid_out;
	input [0:0] SB_T2_NORTH_SB_IN_B1;
	output wire SB_T2_NORTH_SB_IN_B1_enable;
	output wire SB_T2_NORTH_SB_IN_B1_ready_out;
	input SB_T2_NORTH_SB_IN_B1_valid_in;
	output wire [0:0] SB_T2_NORTH_SB_OUT_B1;
	output wire SB_T2_NORTH_SB_OUT_B1_enable;
	input SB_T2_NORTH_SB_OUT_B1_ready_in;
	output wire SB_T2_NORTH_SB_OUT_B1_valid_out;
	input [0:0] SB_T2_SOUTH_SB_IN_B1;
	output wire SB_T2_SOUTH_SB_IN_B1_enable;
	output wire SB_T2_SOUTH_SB_IN_B1_ready_out;
	input SB_T2_SOUTH_SB_IN_B1_valid_in;
	output wire [0:0] SB_T2_SOUTH_SB_OUT_B1;
	output wire SB_T2_SOUTH_SB_OUT_B1_enable;
	input SB_T2_SOUTH_SB_OUT_B1_ready_in;
	output wire SB_T2_SOUTH_SB_OUT_B1_valid_out;
	input [0:0] SB_T2_WEST_SB_IN_B1;
	output wire SB_T2_WEST_SB_IN_B1_enable;
	output wire SB_T2_WEST_SB_IN_B1_ready_out;
	input SB_T2_WEST_SB_IN_B1_valid_in;
	output wire [0:0] SB_T2_WEST_SB_OUT_B1;
	output wire SB_T2_WEST_SB_OUT_B1_enable;
	input SB_T2_WEST_SB_OUT_B1_ready_in;
	output wire SB_T2_WEST_SB_OUT_B1_valid_out;
	input [0:0] SB_T3_EAST_SB_IN_B1;
	output wire SB_T3_EAST_SB_IN_B1_enable;
	output wire SB_T3_EAST_SB_IN_B1_ready_out;
	input SB_T3_EAST_SB_IN_B1_valid_in;
	output wire [0:0] SB_T3_EAST_SB_OUT_B1;
	output wire SB_T3_EAST_SB_OUT_B1_enable;
	input SB_T3_EAST_SB_OUT_B1_ready_in;
	output wire SB_T3_EAST_SB_OUT_B1_valid_out;
	input [0:0] SB_T3_NORTH_SB_IN_B1;
	output wire SB_T3_NORTH_SB_IN_B1_enable;
	output wire SB_T3_NORTH_SB_IN_B1_ready_out;
	input SB_T3_NORTH_SB_IN_B1_valid_in;
	output wire [0:0] SB_T3_NORTH_SB_OUT_B1;
	output wire SB_T3_NORTH_SB_OUT_B1_enable;
	input SB_T3_NORTH_SB_OUT_B1_ready_in;
	output wire SB_T3_NORTH_SB_OUT_B1_valid_out;
	input [0:0] SB_T3_SOUTH_SB_IN_B1;
	output wire SB_T3_SOUTH_SB_IN_B1_enable;
	output wire SB_T3_SOUTH_SB_IN_B1_ready_out;
	input SB_T3_SOUTH_SB_IN_B1_valid_in;
	output wire [0:0] SB_T3_SOUTH_SB_OUT_B1;
	output wire SB_T3_SOUTH_SB_OUT_B1_enable;
	input SB_T3_SOUTH_SB_OUT_B1_ready_in;
	output wire SB_T3_SOUTH_SB_OUT_B1_valid_out;
	input [0:0] SB_T3_WEST_SB_IN_B1;
	output wire SB_T3_WEST_SB_IN_B1_enable;
	output wire SB_T3_WEST_SB_IN_B1_ready_out;
	input SB_T3_WEST_SB_IN_B1_valid_in;
	output wire [0:0] SB_T3_WEST_SB_OUT_B1;
	output wire SB_T3_WEST_SB_OUT_B1_enable;
	input SB_T3_WEST_SB_OUT_B1_ready_in;
	output wire SB_T3_WEST_SB_OUT_B1_valid_out;
	input [0:0] SB_T4_EAST_SB_IN_B1;
	output wire SB_T4_EAST_SB_IN_B1_enable;
	output wire SB_T4_EAST_SB_IN_B1_ready_out;
	input SB_T4_EAST_SB_IN_B1_valid_in;
	output wire [0:0] SB_T4_EAST_SB_OUT_B1;
	output wire SB_T4_EAST_SB_OUT_B1_enable;
	input SB_T4_EAST_SB_OUT_B1_ready_in;
	output wire SB_T4_EAST_SB_OUT_B1_valid_out;
	input [0:0] SB_T4_NORTH_SB_IN_B1;
	output wire SB_T4_NORTH_SB_IN_B1_enable;
	output wire SB_T4_NORTH_SB_IN_B1_ready_out;
	input SB_T4_NORTH_SB_IN_B1_valid_in;
	output wire [0:0] SB_T4_NORTH_SB_OUT_B1;
	output wire SB_T4_NORTH_SB_OUT_B1_enable;
	input SB_T4_NORTH_SB_OUT_B1_ready_in;
	output wire SB_T4_NORTH_SB_OUT_B1_valid_out;
	input [0:0] SB_T4_SOUTH_SB_IN_B1;
	output wire SB_T4_SOUTH_SB_IN_B1_enable;
	output wire SB_T4_SOUTH_SB_IN_B1_ready_out;
	input SB_T4_SOUTH_SB_IN_B1_valid_in;
	output wire [0:0] SB_T4_SOUTH_SB_OUT_B1;
	output wire SB_T4_SOUTH_SB_OUT_B1_enable;
	input SB_T4_SOUTH_SB_OUT_B1_ready_in;
	output wire SB_T4_SOUTH_SB_OUT_B1_valid_out;
	input [0:0] SB_T4_WEST_SB_IN_B1;
	output wire SB_T4_WEST_SB_IN_B1_enable;
	output wire SB_T4_WEST_SB_IN_B1_ready_out;
	input SB_T4_WEST_SB_IN_B1_valid_in;
	output wire [0:0] SB_T4_WEST_SB_OUT_B1;
	output wire SB_T4_WEST_SB_OUT_B1_enable;
	input SB_T4_WEST_SB_OUT_B1_ready_in;
	output wire SB_T4_WEST_SB_OUT_B1_valid_out;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output wire [31:0] read_config_data;
	input reset;
	input [0:0] stall;
	wire [0:0] CB_MEM_output_width_1_num_0_fan_in_O;
	wire [0:0] CB_MEM_output_width_1_num_1_fan_in_O;
	wire [0:0] CB_MEM_output_width_1_num_2_fan_in_O;
	wire [0:0] Invert1_inst0_out;
	wire [0:0] MUX_SB_T0_EAST_SB_OUT_B1_O;
	wire MUX_SB_T0_EAST_SB_OUT_B1_ready_out;
	wire MUX_SB_T0_EAST_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T0_EAST_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T0_NORTH_SB_OUT_B1_O;
	wire MUX_SB_T0_NORTH_SB_OUT_B1_ready_out;
	wire MUX_SB_T0_NORTH_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T0_NORTH_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T0_SOUTH_SB_OUT_B1_O;
	wire MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out;
	wire MUX_SB_T0_SOUTH_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T0_WEST_SB_OUT_B1_O;
	wire MUX_SB_T0_WEST_SB_OUT_B1_ready_out;
	wire MUX_SB_T0_WEST_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T0_WEST_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T1_EAST_SB_OUT_B1_O;
	wire MUX_SB_T1_EAST_SB_OUT_B1_ready_out;
	wire MUX_SB_T1_EAST_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T1_EAST_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T1_NORTH_SB_OUT_B1_O;
	wire MUX_SB_T1_NORTH_SB_OUT_B1_ready_out;
	wire MUX_SB_T1_NORTH_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T1_NORTH_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T1_SOUTH_SB_OUT_B1_O;
	wire MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out;
	wire MUX_SB_T1_SOUTH_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T1_WEST_SB_OUT_B1_O;
	wire MUX_SB_T1_WEST_SB_OUT_B1_ready_out;
	wire MUX_SB_T1_WEST_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T1_WEST_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T2_EAST_SB_OUT_B1_O;
	wire MUX_SB_T2_EAST_SB_OUT_B1_ready_out;
	wire MUX_SB_T2_EAST_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T2_EAST_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T2_NORTH_SB_OUT_B1_O;
	wire MUX_SB_T2_NORTH_SB_OUT_B1_ready_out;
	wire MUX_SB_T2_NORTH_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T2_NORTH_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T2_SOUTH_SB_OUT_B1_O;
	wire MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out;
	wire MUX_SB_T2_SOUTH_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T2_WEST_SB_OUT_B1_O;
	wire MUX_SB_T2_WEST_SB_OUT_B1_ready_out;
	wire MUX_SB_T2_WEST_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T2_WEST_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T3_EAST_SB_OUT_B1_O;
	wire MUX_SB_T3_EAST_SB_OUT_B1_ready_out;
	wire MUX_SB_T3_EAST_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T3_EAST_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T3_NORTH_SB_OUT_B1_O;
	wire MUX_SB_T3_NORTH_SB_OUT_B1_ready_out;
	wire MUX_SB_T3_NORTH_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T3_NORTH_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T3_SOUTH_SB_OUT_B1_O;
	wire MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out;
	wire MUX_SB_T3_SOUTH_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T3_WEST_SB_OUT_B1_O;
	wire MUX_SB_T3_WEST_SB_OUT_B1_ready_out;
	wire MUX_SB_T3_WEST_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T3_WEST_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T4_EAST_SB_OUT_B1_O;
	wire MUX_SB_T4_EAST_SB_OUT_B1_ready_out;
	wire MUX_SB_T4_EAST_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T4_EAST_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T4_NORTH_SB_OUT_B1_O;
	wire MUX_SB_T4_NORTH_SB_OUT_B1_ready_out;
	wire MUX_SB_T4_NORTH_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T4_NORTH_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T4_SOUTH_SB_OUT_B1_O;
	wire MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out;
	wire MUX_SB_T4_SOUTH_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel;
	wire [0:0] MUX_SB_T4_WEST_SB_OUT_B1_O;
	wire MUX_SB_T4_WEST_SB_OUT_B1_ready_out;
	wire MUX_SB_T4_WEST_SB_OUT_B1_valid_out;
	wire [7:0] MUX_SB_T4_WEST_SB_OUT_B1_out_sel;
	wire [0:0] REG_T0_EAST_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T0_EAST_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T0_EAST_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T0_EAST_B1_end_value_O;
	wire [0:0] REG_T0_EAST_B1_fifo_value_O;
	wire [0:0] REG_T0_EAST_B1_start_value_O;
	wire [0:0] REG_T0_NORTH_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T0_NORTH_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T0_NORTH_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T0_NORTH_B1_end_value_O;
	wire [0:0] REG_T0_NORTH_B1_fifo_value_O;
	wire [0:0] REG_T0_NORTH_B1_start_value_O;
	wire [0:0] REG_T0_SOUTH_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T0_SOUTH_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T0_SOUTH_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T0_SOUTH_B1_end_value_O;
	wire [0:0] REG_T0_SOUTH_B1_fifo_value_O;
	wire [0:0] REG_T0_SOUTH_B1_start_value_O;
	wire [0:0] REG_T0_WEST_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T0_WEST_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T0_WEST_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T0_WEST_B1_end_value_O;
	wire [0:0] REG_T0_WEST_B1_fifo_value_O;
	wire [0:0] REG_T0_WEST_B1_start_value_O;
	wire [0:0] REG_T1_EAST_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T1_EAST_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T1_EAST_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T1_EAST_B1_end_value_O;
	wire [0:0] REG_T1_EAST_B1_fifo_value_O;
	wire [0:0] REG_T1_EAST_B1_start_value_O;
	wire [0:0] REG_T1_NORTH_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T1_NORTH_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T1_NORTH_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T1_NORTH_B1_end_value_O;
	wire [0:0] REG_T1_NORTH_B1_fifo_value_O;
	wire [0:0] REG_T1_NORTH_B1_start_value_O;
	wire [0:0] REG_T1_SOUTH_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T1_SOUTH_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T1_SOUTH_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T1_SOUTH_B1_end_value_O;
	wire [0:0] REG_T1_SOUTH_B1_fifo_value_O;
	wire [0:0] REG_T1_SOUTH_B1_start_value_O;
	wire [0:0] REG_T1_WEST_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T1_WEST_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T1_WEST_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T1_WEST_B1_end_value_O;
	wire [0:0] REG_T1_WEST_B1_fifo_value_O;
	wire [0:0] REG_T1_WEST_B1_start_value_O;
	wire [0:0] REG_T2_EAST_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T2_EAST_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T2_EAST_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T2_EAST_B1_end_value_O;
	wire [0:0] REG_T2_EAST_B1_fifo_value_O;
	wire [0:0] REG_T2_EAST_B1_start_value_O;
	wire [0:0] REG_T2_NORTH_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T2_NORTH_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T2_NORTH_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T2_NORTH_B1_end_value_O;
	wire [0:0] REG_T2_NORTH_B1_fifo_value_O;
	wire [0:0] REG_T2_NORTH_B1_start_value_O;
	wire [0:0] REG_T2_SOUTH_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T2_SOUTH_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T2_SOUTH_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T2_SOUTH_B1_end_value_O;
	wire [0:0] REG_T2_SOUTH_B1_fifo_value_O;
	wire [0:0] REG_T2_SOUTH_B1_start_value_O;
	wire [0:0] REG_T2_WEST_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T2_WEST_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T2_WEST_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T2_WEST_B1_end_value_O;
	wire [0:0] REG_T2_WEST_B1_fifo_value_O;
	wire [0:0] REG_T2_WEST_B1_start_value_O;
	wire [0:0] REG_T3_EAST_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T3_EAST_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T3_EAST_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T3_EAST_B1_end_value_O;
	wire [0:0] REG_T3_EAST_B1_fifo_value_O;
	wire [0:0] REG_T3_EAST_B1_start_value_O;
	wire [0:0] REG_T3_NORTH_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T3_NORTH_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T3_NORTH_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T3_NORTH_B1_end_value_O;
	wire [0:0] REG_T3_NORTH_B1_fifo_value_O;
	wire [0:0] REG_T3_NORTH_B1_start_value_O;
	wire [0:0] REG_T3_SOUTH_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T3_SOUTH_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T3_SOUTH_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T3_SOUTH_B1_end_value_O;
	wire [0:0] REG_T3_SOUTH_B1_fifo_value_O;
	wire [0:0] REG_T3_SOUTH_B1_start_value_O;
	wire [0:0] REG_T3_WEST_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T3_WEST_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T3_WEST_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T3_WEST_B1_end_value_O;
	wire [0:0] REG_T3_WEST_B1_fifo_value_O;
	wire [0:0] REG_T3_WEST_B1_start_value_O;
	wire [0:0] REG_T4_EAST_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T4_EAST_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T4_EAST_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T4_EAST_B1_end_value_O;
	wire [0:0] REG_T4_EAST_B1_fifo_value_O;
	wire [0:0] REG_T4_EAST_B1_start_value_O;
	wire [0:0] REG_T4_NORTH_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T4_NORTH_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T4_NORTH_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T4_NORTH_B1_end_value_O;
	wire [0:0] REG_T4_NORTH_B1_fifo_value_O;
	wire [0:0] REG_T4_NORTH_B1_start_value_O;
	wire [0:0] REG_T4_SOUTH_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T4_SOUTH_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T4_SOUTH_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T4_SOUTH_B1_end_value_O;
	wire [0:0] REG_T4_SOUTH_B1_fifo_value_O;
	wire [0:0] REG_T4_SOUTH_B1_start_value_O;
	wire [0:0] REG_T4_WEST_B1$SplitFifo_1_inst0_ready0;
	wire [0:0] REG_T4_WEST_B1$SplitFifo_1_inst0_data_out;
	wire [0:0] REG_T4_WEST_B1$SplitFifo_1_inst0_valid1;
	wire [0:0] REG_T4_WEST_B1_end_value_O;
	wire [0:0] REG_T4_WEST_B1_fifo_value_O;
	wire [0:0] REG_T4_WEST_B1_start_value_O;
	wire [0:0] RMUX_T0_EAST_B1_O;
	wire RMUX_T0_EAST_B1_ready_out;
	wire RMUX_T0_EAST_B1_valid_out;
	wire [1:0] RMUX_T0_EAST_B1_out_sel;
	wire [0:0] RMUX_T0_EAST_B1_sel_value_O;
	wire [0:0] RMUX_T0_NORTH_B1_O;
	wire RMUX_T0_NORTH_B1_ready_out;
	wire RMUX_T0_NORTH_B1_valid_out;
	wire [1:0] RMUX_T0_NORTH_B1_out_sel;
	wire [0:0] RMUX_T0_NORTH_B1_sel_value_O;
	wire [0:0] RMUX_T0_SOUTH_B1_O;
	wire RMUX_T0_SOUTH_B1_ready_out;
	wire RMUX_T0_SOUTH_B1_valid_out;
	wire [1:0] RMUX_T0_SOUTH_B1_out_sel;
	wire [0:0] RMUX_T0_SOUTH_B1_sel_value_O;
	wire [0:0] RMUX_T0_WEST_B1_O;
	wire RMUX_T0_WEST_B1_ready_out;
	wire RMUX_T0_WEST_B1_valid_out;
	wire [1:0] RMUX_T0_WEST_B1_out_sel;
	wire [0:0] RMUX_T0_WEST_B1_sel_value_O;
	wire [0:0] RMUX_T1_EAST_B1_O;
	wire RMUX_T1_EAST_B1_ready_out;
	wire RMUX_T1_EAST_B1_valid_out;
	wire [1:0] RMUX_T1_EAST_B1_out_sel;
	wire [0:0] RMUX_T1_EAST_B1_sel_value_O;
	wire [0:0] RMUX_T1_NORTH_B1_O;
	wire RMUX_T1_NORTH_B1_ready_out;
	wire RMUX_T1_NORTH_B1_valid_out;
	wire [1:0] RMUX_T1_NORTH_B1_out_sel;
	wire [0:0] RMUX_T1_NORTH_B1_sel_value_O;
	wire [0:0] RMUX_T1_SOUTH_B1_O;
	wire RMUX_T1_SOUTH_B1_ready_out;
	wire RMUX_T1_SOUTH_B1_valid_out;
	wire [1:0] RMUX_T1_SOUTH_B1_out_sel;
	wire [0:0] RMUX_T1_SOUTH_B1_sel_value_O;
	wire [0:0] RMUX_T1_WEST_B1_O;
	wire RMUX_T1_WEST_B1_ready_out;
	wire RMUX_T1_WEST_B1_valid_out;
	wire [1:0] RMUX_T1_WEST_B1_out_sel;
	wire [0:0] RMUX_T1_WEST_B1_sel_value_O;
	wire [0:0] RMUX_T2_EAST_B1_O;
	wire RMUX_T2_EAST_B1_ready_out;
	wire RMUX_T2_EAST_B1_valid_out;
	wire [1:0] RMUX_T2_EAST_B1_out_sel;
	wire [0:0] RMUX_T2_EAST_B1_sel_value_O;
	wire [0:0] RMUX_T2_NORTH_B1_O;
	wire RMUX_T2_NORTH_B1_ready_out;
	wire RMUX_T2_NORTH_B1_valid_out;
	wire [1:0] RMUX_T2_NORTH_B1_out_sel;
	wire [0:0] RMUX_T2_NORTH_B1_sel_value_O;
	wire [0:0] RMUX_T2_SOUTH_B1_O;
	wire RMUX_T2_SOUTH_B1_ready_out;
	wire RMUX_T2_SOUTH_B1_valid_out;
	wire [1:0] RMUX_T2_SOUTH_B1_out_sel;
	wire [0:0] RMUX_T2_SOUTH_B1_sel_value_O;
	wire [0:0] RMUX_T2_WEST_B1_O;
	wire RMUX_T2_WEST_B1_ready_out;
	wire RMUX_T2_WEST_B1_valid_out;
	wire [1:0] RMUX_T2_WEST_B1_out_sel;
	wire [0:0] RMUX_T2_WEST_B1_sel_value_O;
	wire [0:0] RMUX_T3_EAST_B1_O;
	wire RMUX_T3_EAST_B1_ready_out;
	wire RMUX_T3_EAST_B1_valid_out;
	wire [1:0] RMUX_T3_EAST_B1_out_sel;
	wire [0:0] RMUX_T3_EAST_B1_sel_value_O;
	wire [0:0] RMUX_T3_NORTH_B1_O;
	wire RMUX_T3_NORTH_B1_ready_out;
	wire RMUX_T3_NORTH_B1_valid_out;
	wire [1:0] RMUX_T3_NORTH_B1_out_sel;
	wire [0:0] RMUX_T3_NORTH_B1_sel_value_O;
	wire [0:0] RMUX_T3_SOUTH_B1_O;
	wire RMUX_T3_SOUTH_B1_ready_out;
	wire RMUX_T3_SOUTH_B1_valid_out;
	wire [1:0] RMUX_T3_SOUTH_B1_out_sel;
	wire [0:0] RMUX_T3_SOUTH_B1_sel_value_O;
	wire [0:0] RMUX_T3_WEST_B1_O;
	wire RMUX_T3_WEST_B1_ready_out;
	wire RMUX_T3_WEST_B1_valid_out;
	wire [1:0] RMUX_T3_WEST_B1_out_sel;
	wire [0:0] RMUX_T3_WEST_B1_sel_value_O;
	wire [0:0] RMUX_T4_EAST_B1_O;
	wire RMUX_T4_EAST_B1_ready_out;
	wire RMUX_T4_EAST_B1_valid_out;
	wire [1:0] RMUX_T4_EAST_B1_out_sel;
	wire [0:0] RMUX_T4_EAST_B1_sel_value_O;
	wire [0:0] RMUX_T4_NORTH_B1_O;
	wire RMUX_T4_NORTH_B1_ready_out;
	wire RMUX_T4_NORTH_B1_valid_out;
	wire [1:0] RMUX_T4_NORTH_B1_out_sel;
	wire [0:0] RMUX_T4_NORTH_B1_sel_value_O;
	wire [0:0] RMUX_T4_SOUTH_B1_O;
	wire RMUX_T4_SOUTH_B1_ready_out;
	wire RMUX_T4_SOUTH_B1_valid_out;
	wire [1:0] RMUX_T4_SOUTH_B1_out_sel;
	wire [0:0] RMUX_T4_SOUTH_B1_sel_value_O;
	wire [0:0] RMUX_T4_WEST_B1_O;
	wire RMUX_T4_WEST_B1_ready_out;
	wire RMUX_T4_WEST_B1_valid_out;
	wire [1:0] RMUX_T4_WEST_B1_out_sel;
	wire [0:0] RMUX_T4_WEST_B1_sel_value_O;
	wire [0:0] SB_T0_EAST_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T0_EAST_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T0_EAST_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T0_EAST_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T0_EAST_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T0_NORTH_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T0_NORTH_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T0_NORTH_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T0_NORTH_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T0_NORTH_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T0_SOUTH_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T0_SOUTH_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T0_SOUTH_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T0_SOUTH_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T0_SOUTH_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T0_WEST_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T0_WEST_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T0_WEST_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T0_WEST_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T0_WEST_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T1_EAST_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T1_EAST_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T1_EAST_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T1_EAST_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T1_EAST_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T1_NORTH_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T1_NORTH_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T1_NORTH_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T1_NORTH_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T1_NORTH_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T1_SOUTH_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T1_SOUTH_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T1_SOUTH_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T1_SOUTH_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T1_SOUTH_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T1_WEST_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T1_WEST_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T1_WEST_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T1_WEST_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T1_WEST_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T2_EAST_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T2_EAST_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T2_EAST_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T2_EAST_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T2_EAST_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T2_NORTH_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T2_NORTH_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T2_NORTH_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T2_NORTH_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T2_NORTH_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T2_SOUTH_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T2_SOUTH_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T2_SOUTH_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T2_SOUTH_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T2_SOUTH_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T2_WEST_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T2_WEST_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T2_WEST_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T2_WEST_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T2_WEST_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T3_EAST_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T3_EAST_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T3_EAST_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T3_EAST_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T3_EAST_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T3_NORTH_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T3_NORTH_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T3_NORTH_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T3_NORTH_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T3_NORTH_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T3_SOUTH_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T3_SOUTH_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T3_SOUTH_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T3_SOUTH_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T3_SOUTH_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T3_WEST_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T3_WEST_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T3_WEST_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T3_WEST_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T3_WEST_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T4_EAST_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T4_EAST_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T4_EAST_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T4_EAST_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T4_EAST_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T4_NORTH_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T4_NORTH_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T4_NORTH_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T4_NORTH_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T4_NORTH_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T4_SOUTH_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T4_SOUTH_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T4_SOUTH_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T4_SOUTH_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T4_SOUTH_SB_OUT_B1_sel_value_O;
	wire [0:0] SB_T4_WEST_SB_IN_B1_enable_value_O;
	wire [0:0] SB_T4_WEST_SB_IN_B1_fan_in_O;
	wire [0:0] SB_T4_WEST_SB_OUT_B1_FANOUT_O;
	wire [0:0] SB_T4_WEST_SB_OUT_B1_enable_value_O;
	wire [2:0] SB_T4_WEST_SB_OUT_B1_sel_value_O;
	wire [0:0] WIRE_SB_T0_EAST_SB_IN_B1_O;
	wire WIRE_SB_T0_EAST_SB_IN_B1_ready_out;
	wire WIRE_SB_T0_EAST_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T0_NORTH_SB_IN_B1_O;
	wire WIRE_SB_T0_NORTH_SB_IN_B1_ready_out;
	wire WIRE_SB_T0_NORTH_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T0_SOUTH_SB_IN_B1_O;
	wire WIRE_SB_T0_SOUTH_SB_IN_B1_ready_out;
	wire WIRE_SB_T0_SOUTH_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T0_WEST_SB_IN_B1_O;
	wire WIRE_SB_T0_WEST_SB_IN_B1_ready_out;
	wire WIRE_SB_T0_WEST_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T1_EAST_SB_IN_B1_O;
	wire WIRE_SB_T1_EAST_SB_IN_B1_ready_out;
	wire WIRE_SB_T1_EAST_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T1_NORTH_SB_IN_B1_O;
	wire WIRE_SB_T1_NORTH_SB_IN_B1_ready_out;
	wire WIRE_SB_T1_NORTH_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T1_SOUTH_SB_IN_B1_O;
	wire WIRE_SB_T1_SOUTH_SB_IN_B1_ready_out;
	wire WIRE_SB_T1_SOUTH_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T1_WEST_SB_IN_B1_O;
	wire WIRE_SB_T1_WEST_SB_IN_B1_ready_out;
	wire WIRE_SB_T1_WEST_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T2_EAST_SB_IN_B1_O;
	wire WIRE_SB_T2_EAST_SB_IN_B1_ready_out;
	wire WIRE_SB_T2_EAST_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T2_NORTH_SB_IN_B1_O;
	wire WIRE_SB_T2_NORTH_SB_IN_B1_ready_out;
	wire WIRE_SB_T2_NORTH_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T2_SOUTH_SB_IN_B1_O;
	wire WIRE_SB_T2_SOUTH_SB_IN_B1_ready_out;
	wire WIRE_SB_T2_SOUTH_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T2_WEST_SB_IN_B1_O;
	wire WIRE_SB_T2_WEST_SB_IN_B1_ready_out;
	wire WIRE_SB_T2_WEST_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T3_EAST_SB_IN_B1_O;
	wire WIRE_SB_T3_EAST_SB_IN_B1_ready_out;
	wire WIRE_SB_T3_EAST_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T3_NORTH_SB_IN_B1_O;
	wire WIRE_SB_T3_NORTH_SB_IN_B1_ready_out;
	wire WIRE_SB_T3_NORTH_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T3_SOUTH_SB_IN_B1_O;
	wire WIRE_SB_T3_SOUTH_SB_IN_B1_ready_out;
	wire WIRE_SB_T3_SOUTH_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T3_WEST_SB_IN_B1_O;
	wire WIRE_SB_T3_WEST_SB_IN_B1_ready_out;
	wire WIRE_SB_T3_WEST_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T4_EAST_SB_IN_B1_O;
	wire WIRE_SB_T4_EAST_SB_IN_B1_ready_out;
	wire WIRE_SB_T4_EAST_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T4_NORTH_SB_IN_B1_O;
	wire WIRE_SB_T4_NORTH_SB_IN_B1_ready_out;
	wire WIRE_SB_T4_NORTH_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T4_SOUTH_SB_IN_B1_O;
	wire WIRE_SB_T4_SOUTH_SB_IN_B1_ready_out;
	wire WIRE_SB_T4_SOUTH_SB_IN_B1_valid_out;
	wire [0:0] WIRE_SB_T4_WEST_SB_IN_B1_O;
	wire WIRE_SB_T4_WEST_SB_IN_B1_ready_out;
	wire WIRE_SB_T4_WEST_SB_IN_B1_valid_out;
	wire ZextWrapper_23_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_23_32_inst0$self_O_in;
	wire ZextWrapper_30_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_30_32_inst0$self_O_in;
	wire ZextWrapper_31_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_31_32_inst0$self_O_in;
	wire [0:0] and1_inst0_out;
	wire [0:0] and1_inst1_out;
	wire [0:0] and1_inst10_out;
	wire [0:0] and1_inst11_out;
	wire [0:0] and1_inst12_out;
	wire [0:0] and1_inst13_out;
	wire [0:0] and1_inst14_out;
	wire [0:0] and1_inst15_out;
	wire [0:0] and1_inst16_out;
	wire [0:0] and1_inst17_out;
	wire [0:0] and1_inst18_out;
	wire [0:0] and1_inst19_out;
	wire [0:0] and1_inst2_out;
	wire [0:0] and1_inst3_out;
	wire [0:0] and1_inst4_out;
	wire [0:0] and1_inst5_out;
	wire [0:0] and1_inst6_out;
	wire [0:0] and1_inst7_out;
	wire [0:0] and1_inst8_out;
	wire [0:0] and1_inst9_out;
	wire [31:0] config_reg_0_O;
	wire [31:0] config_reg_1_O;
	wire [31:0] config_reg_2_O;
	wire [30:0] config_reg_3_O;
	wire [29:0] config_reg_4_O;
	wire [22:0] config_reg_5_O;
	wire [0:0] const_0_1_out;
	wire [31:0] const_0_32_out;
	wire [0:0] const_1_1_out;
	wire coreir_eq_1_inst0_out;
	wire coreir_eq_1_inst1_out;
	wire coreir_eq_1_inst10_out;
	wire coreir_eq_1_inst11_out;
	wire coreir_eq_1_inst12_out;
	wire coreir_eq_1_inst13_out;
	wire coreir_eq_1_inst14_out;
	wire coreir_eq_1_inst15_out;
	wire coreir_eq_1_inst16_out;
	wire coreir_eq_1_inst17_out;
	wire coreir_eq_1_inst18_out;
	wire coreir_eq_1_inst19_out;
	wire coreir_eq_1_inst2_out;
	wire coreir_eq_1_inst3_out;
	wire coreir_eq_1_inst4_out;
	wire coreir_eq_1_inst5_out;
	wire coreir_eq_1_inst6_out;
	wire coreir_eq_1_inst7_out;
	wire coreir_eq_1_inst8_out;
	wire coreir_eq_1_inst9_out;
	wire [31:0] mux_aoi_6_32_inst0_O;
	wire [7:0] mux_aoi_6_32_inst0_out_sel;
	wire [7:0] self_config_config_addr_out;
	FanoutHash_E70AF988E4250F5 CB_MEM_output_width_1_num_0_fan_in(
		.I13(MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out),
		.E8(SB_T2_NORTH_SB_OUT_B1_enable_value_O),
		.E17(SB_T4_SOUTH_SB_OUT_B1_enable_value_O),
		.I15(MUX_SB_T3_WEST_SB_OUT_B1_ready_out),
		.I12(MUX_SB_T3_NORTH_SB_OUT_B1_ready_out),
		.E6(SB_T1_EAST_SB_OUT_B1_enable_value_O),
		.I9(MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out),
		.I16(MUX_SB_T4_NORTH_SB_OUT_B1_ready_out),
		.E3(SB_T0_WEST_SB_OUT_B1_enable_value_O),
		.S14(MUX_SB_T3_EAST_SB_OUT_B1_out_sel),
		.E10(SB_T2_EAST_SB_OUT_B1_enable_value_O),
		.I5(MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out),
		.S6(MUX_SB_T1_EAST_SB_OUT_B1_out_sel),
		.E0(SB_T0_NORTH_SB_OUT_B1_enable_value_O),
		.E18(SB_T4_EAST_SB_OUT_B1_enable_value_O),
		.I19(MUX_SB_T4_WEST_SB_OUT_B1_ready_out),
		.I10(MUX_SB_T2_EAST_SB_OUT_B1_ready_out),
		.S5(MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel),
		.I6(MUX_SB_T1_EAST_SB_OUT_B1_ready_out),
		.I8(MUX_SB_T2_NORTH_SB_OUT_B1_ready_out),
		.S3(MUX_SB_T0_WEST_SB_OUT_B1_out_sel),
		.S10(MUX_SB_T2_EAST_SB_OUT_B1_out_sel),
		.E16(SB_T4_NORTH_SB_OUT_B1_enable_value_O),
		.S4(MUX_SB_T1_NORTH_SB_OUT_B1_out_sel),
		.E11(SB_T2_WEST_SB_OUT_B1_enable_value_O),
		.S19(MUX_SB_T4_WEST_SB_OUT_B1_out_sel),
		.E15(SB_T3_WEST_SB_OUT_B1_enable_value_O),
		.E19(SB_T4_WEST_SB_OUT_B1_enable_value_O),
		.I3(MUX_SB_T0_WEST_SB_OUT_B1_ready_out),
		.I4(MUX_SB_T1_NORTH_SB_OUT_B1_ready_out),
		.S1(MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel),
		.E13(SB_T3_SOUTH_SB_OUT_B1_enable_value_O),
		.S0(MUX_SB_T0_NORTH_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T0_EAST_SB_OUT_B1_out_sel),
		.I11(MUX_SB_T2_WEST_SB_OUT_B1_ready_out),
		.S8(MUX_SB_T2_NORTH_SB_OUT_B1_out_sel),
		.E2(SB_T0_EAST_SB_OUT_B1_enable_value_O),
		.E14(SB_T3_EAST_SB_OUT_B1_enable_value_O),
		.S17(MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel),
		.E5(SB_T1_SOUTH_SB_OUT_B1_enable_value_O),
		.E4(SB_T1_NORTH_SB_OUT_B1_enable_value_O),
		.I1(MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out),
		.I2(MUX_SB_T0_EAST_SB_OUT_B1_ready_out),
		.I17(MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out),
		.O(CB_MEM_output_width_1_num_0_fan_in_O),
		.E9(SB_T2_SOUTH_SB_OUT_B1_enable_value_O),
		.S13(MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel),
		.S11(MUX_SB_T2_WEST_SB_OUT_B1_out_sel),
		.S7(MUX_SB_T1_WEST_SB_OUT_B1_out_sel),
		.E1(SB_T0_SOUTH_SB_OUT_B1_enable_value_O),
		.S15(MUX_SB_T3_WEST_SB_OUT_B1_out_sel),
		.S9(MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel),
		.S18(MUX_SB_T4_EAST_SB_OUT_B1_out_sel),
		.S12(MUX_SB_T3_NORTH_SB_OUT_B1_out_sel),
		.I14(MUX_SB_T3_EAST_SB_OUT_B1_ready_out),
		.I7(MUX_SB_T1_WEST_SB_OUT_B1_ready_out),
		.S16(MUX_SB_T4_NORTH_SB_OUT_B1_out_sel),
		.E12(SB_T3_NORTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T0_NORTH_SB_OUT_B1_ready_out),
		.E7(SB_T1_WEST_SB_OUT_B1_enable_value_O),
		.I18(MUX_SB_T4_EAST_SB_OUT_B1_ready_out)
	);
	FanoutHash_82899D6851EDC11 CB_MEM_output_width_1_num_1_fan_in(
		.I13(MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out),
		.E8(SB_T2_NORTH_SB_OUT_B1_enable_value_O),
		.E17(SB_T4_SOUTH_SB_OUT_B1_enable_value_O),
		.I15(MUX_SB_T3_WEST_SB_OUT_B1_ready_out),
		.I12(MUX_SB_T3_NORTH_SB_OUT_B1_ready_out),
		.E6(SB_T1_EAST_SB_OUT_B1_enable_value_O),
		.I9(MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out),
		.I16(MUX_SB_T4_NORTH_SB_OUT_B1_ready_out),
		.E3(SB_T0_WEST_SB_OUT_B1_enable_value_O),
		.S14(MUX_SB_T3_EAST_SB_OUT_B1_out_sel),
		.E10(SB_T2_EAST_SB_OUT_B1_enable_value_O),
		.I5(MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out),
		.S6(MUX_SB_T1_EAST_SB_OUT_B1_out_sel),
		.E0(SB_T0_NORTH_SB_OUT_B1_enable_value_O),
		.E18(SB_T4_EAST_SB_OUT_B1_enable_value_O),
		.I19(MUX_SB_T4_WEST_SB_OUT_B1_ready_out),
		.I10(MUX_SB_T2_EAST_SB_OUT_B1_ready_out),
		.S5(MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel),
		.I6(MUX_SB_T1_EAST_SB_OUT_B1_ready_out),
		.I8(MUX_SB_T2_NORTH_SB_OUT_B1_ready_out),
		.S3(MUX_SB_T0_WEST_SB_OUT_B1_out_sel),
		.S10(MUX_SB_T2_EAST_SB_OUT_B1_out_sel),
		.E16(SB_T4_NORTH_SB_OUT_B1_enable_value_O),
		.S4(MUX_SB_T1_NORTH_SB_OUT_B1_out_sel),
		.E11(SB_T2_WEST_SB_OUT_B1_enable_value_O),
		.S19(MUX_SB_T4_WEST_SB_OUT_B1_out_sel),
		.E15(SB_T3_WEST_SB_OUT_B1_enable_value_O),
		.E19(SB_T4_WEST_SB_OUT_B1_enable_value_O),
		.I3(MUX_SB_T0_WEST_SB_OUT_B1_ready_out),
		.I4(MUX_SB_T1_NORTH_SB_OUT_B1_ready_out),
		.S1(MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel),
		.E13(SB_T3_SOUTH_SB_OUT_B1_enable_value_O),
		.S0(MUX_SB_T0_NORTH_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T0_EAST_SB_OUT_B1_out_sel),
		.I11(MUX_SB_T2_WEST_SB_OUT_B1_ready_out),
		.S8(MUX_SB_T2_NORTH_SB_OUT_B1_out_sel),
		.E2(SB_T0_EAST_SB_OUT_B1_enable_value_O),
		.E14(SB_T3_EAST_SB_OUT_B1_enable_value_O),
		.S17(MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel),
		.E5(SB_T1_SOUTH_SB_OUT_B1_enable_value_O),
		.E4(SB_T1_NORTH_SB_OUT_B1_enable_value_O),
		.I1(MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out),
		.I2(MUX_SB_T0_EAST_SB_OUT_B1_ready_out),
		.I17(MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out),
		.O(CB_MEM_output_width_1_num_1_fan_in_O),
		.E9(SB_T2_SOUTH_SB_OUT_B1_enable_value_O),
		.S13(MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel),
		.S11(MUX_SB_T2_WEST_SB_OUT_B1_out_sel),
		.S7(MUX_SB_T1_WEST_SB_OUT_B1_out_sel),
		.E1(SB_T0_SOUTH_SB_OUT_B1_enable_value_O),
		.S15(MUX_SB_T3_WEST_SB_OUT_B1_out_sel),
		.S9(MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel),
		.S18(MUX_SB_T4_EAST_SB_OUT_B1_out_sel),
		.S12(MUX_SB_T3_NORTH_SB_OUT_B1_out_sel),
		.I14(MUX_SB_T3_EAST_SB_OUT_B1_ready_out),
		.I7(MUX_SB_T1_WEST_SB_OUT_B1_ready_out),
		.S16(MUX_SB_T4_NORTH_SB_OUT_B1_out_sel),
		.E12(SB_T3_NORTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T0_NORTH_SB_OUT_B1_ready_out),
		.E7(SB_T1_WEST_SB_OUT_B1_enable_value_O),
		.I18(MUX_SB_T4_EAST_SB_OUT_B1_ready_out)
	);
	FanoutHash_CE1AA874B742213 CB_MEM_output_width_1_num_2_fan_in(
		.I13(MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out),
		.E8(SB_T2_NORTH_SB_OUT_B1_enable_value_O),
		.E17(SB_T4_SOUTH_SB_OUT_B1_enable_value_O),
		.I15(MUX_SB_T3_WEST_SB_OUT_B1_ready_out),
		.I12(MUX_SB_T3_NORTH_SB_OUT_B1_ready_out),
		.E6(SB_T1_EAST_SB_OUT_B1_enable_value_O),
		.I9(MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out),
		.I16(MUX_SB_T4_NORTH_SB_OUT_B1_ready_out),
		.E3(SB_T0_WEST_SB_OUT_B1_enable_value_O),
		.S14(MUX_SB_T3_EAST_SB_OUT_B1_out_sel),
		.E10(SB_T2_EAST_SB_OUT_B1_enable_value_O),
		.I5(MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out),
		.S6(MUX_SB_T1_EAST_SB_OUT_B1_out_sel),
		.E0(SB_T0_NORTH_SB_OUT_B1_enable_value_O),
		.E18(SB_T4_EAST_SB_OUT_B1_enable_value_O),
		.I19(MUX_SB_T4_WEST_SB_OUT_B1_ready_out),
		.I10(MUX_SB_T2_EAST_SB_OUT_B1_ready_out),
		.S5(MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel),
		.I6(MUX_SB_T1_EAST_SB_OUT_B1_ready_out),
		.I8(MUX_SB_T2_NORTH_SB_OUT_B1_ready_out),
		.S3(MUX_SB_T0_WEST_SB_OUT_B1_out_sel),
		.S10(MUX_SB_T2_EAST_SB_OUT_B1_out_sel),
		.E16(SB_T4_NORTH_SB_OUT_B1_enable_value_O),
		.S4(MUX_SB_T1_NORTH_SB_OUT_B1_out_sel),
		.E11(SB_T2_WEST_SB_OUT_B1_enable_value_O),
		.S19(MUX_SB_T4_WEST_SB_OUT_B1_out_sel),
		.E15(SB_T3_WEST_SB_OUT_B1_enable_value_O),
		.E19(SB_T4_WEST_SB_OUT_B1_enable_value_O),
		.I3(MUX_SB_T0_WEST_SB_OUT_B1_ready_out),
		.I4(MUX_SB_T1_NORTH_SB_OUT_B1_ready_out),
		.S1(MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel),
		.E13(SB_T3_SOUTH_SB_OUT_B1_enable_value_O),
		.S0(MUX_SB_T0_NORTH_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T0_EAST_SB_OUT_B1_out_sel),
		.I11(MUX_SB_T2_WEST_SB_OUT_B1_ready_out),
		.S8(MUX_SB_T2_NORTH_SB_OUT_B1_out_sel),
		.E2(SB_T0_EAST_SB_OUT_B1_enable_value_O),
		.E14(SB_T3_EAST_SB_OUT_B1_enable_value_O),
		.S17(MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel),
		.E5(SB_T1_SOUTH_SB_OUT_B1_enable_value_O),
		.E4(SB_T1_NORTH_SB_OUT_B1_enable_value_O),
		.I1(MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out),
		.I2(MUX_SB_T0_EAST_SB_OUT_B1_ready_out),
		.I17(MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out),
		.O(CB_MEM_output_width_1_num_2_fan_in_O),
		.E9(SB_T2_SOUTH_SB_OUT_B1_enable_value_O),
		.S13(MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel),
		.S11(MUX_SB_T2_WEST_SB_OUT_B1_out_sel),
		.S7(MUX_SB_T1_WEST_SB_OUT_B1_out_sel),
		.E1(SB_T0_SOUTH_SB_OUT_B1_enable_value_O),
		.S15(MUX_SB_T3_WEST_SB_OUT_B1_out_sel),
		.S9(MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel),
		.S18(MUX_SB_T4_EAST_SB_OUT_B1_out_sel),
		.S12(MUX_SB_T3_NORTH_SB_OUT_B1_out_sel),
		.I14(MUX_SB_T3_EAST_SB_OUT_B1_ready_out),
		.I7(MUX_SB_T1_WEST_SB_OUT_B1_ready_out),
		.S16(MUX_SB_T4_NORTH_SB_OUT_B1_out_sel),
		.E12(SB_T3_NORTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T0_NORTH_SB_OUT_B1_ready_out),
		.E7(SB_T1_WEST_SB_OUT_B1_enable_value_O),
		.I18(MUX_SB_T4_EAST_SB_OUT_B1_ready_out)
	);
	coreir_not #(.width(1)) Invert1_inst0(
		.in(stall),
		.out(Invert1_inst0_out)
	);
	wire [5:0] MUX_SB_T0_EAST_SB_OUT_B1_I;
	assign MUX_SB_T0_EAST_SB_OUT_B1_I[5+:1] = MEM_output_width_1_num_2;
	assign MUX_SB_T0_EAST_SB_OUT_B1_I[4+:1] = MEM_output_width_1_num_1;
	assign MUX_SB_T0_EAST_SB_OUT_B1_I[3+:1] = MEM_output_width_1_num_0;
	assign MUX_SB_T0_EAST_SB_OUT_B1_I[2+:1] = WIRE_SB_T4_NORTH_SB_IN_B1_O;
	assign MUX_SB_T0_EAST_SB_OUT_B1_I[1+:1] = WIRE_SB_T3_SOUTH_SB_IN_B1_O;
	assign MUX_SB_T0_EAST_SB_OUT_B1_I[0+:1] = WIRE_SB_T0_WEST_SB_IN_B1_O;
	wire [5:0] MUX_SB_T0_EAST_SB_OUT_B1_valid_in;
	assign MUX_SB_T0_EAST_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid, MEM_output_width_1_num_1_valid, MEM_output_width_1_num_0_valid, WIRE_SB_T4_NORTH_SB_IN_B1_valid_out, WIRE_SB_T3_SOUTH_SB_IN_B1_valid_out, WIRE_SB_T0_WEST_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T0_EAST_SB_OUT_B1(
		.I(MUX_SB_T0_EAST_SB_OUT_B1_I),
		.O(MUX_SB_T0_EAST_SB_OUT_B1_O),
		.ready_in(SB_T0_EAST_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T0_EAST_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T0_EAST_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T0_EAST_SB_OUT_B1_valid_out),
		.S(SB_T0_EAST_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T0_EAST_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T0_NORTH_SB_OUT_B1_I;
	assign MUX_SB_T0_NORTH_SB_OUT_B1_I[5+:1] = MEM_output_width_1_num_2;
	assign MUX_SB_T0_NORTH_SB_OUT_B1_I[4+:1] = MEM_output_width_1_num_1;
	assign MUX_SB_T0_NORTH_SB_OUT_B1_I[3+:1] = MEM_output_width_1_num_0;
	assign MUX_SB_T0_NORTH_SB_OUT_B1_I[2+:1] = WIRE_SB_T0_SOUTH_SB_IN_B1_O;
	assign MUX_SB_T0_NORTH_SB_OUT_B1_I[1+:1] = WIRE_SB_T1_EAST_SB_IN_B1_O;
	assign MUX_SB_T0_NORTH_SB_OUT_B1_I[0+:1] = WIRE_SB_T0_WEST_SB_IN_B1_O;
	wire [5:0] MUX_SB_T0_NORTH_SB_OUT_B1_valid_in;
	assign MUX_SB_T0_NORTH_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid, MEM_output_width_1_num_1_valid, MEM_output_width_1_num_0_valid, WIRE_SB_T0_SOUTH_SB_IN_B1_valid_out, WIRE_SB_T1_EAST_SB_IN_B1_valid_out, WIRE_SB_T0_WEST_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T0_NORTH_SB_OUT_B1(
		.I(MUX_SB_T0_NORTH_SB_OUT_B1_I),
		.O(MUX_SB_T0_NORTH_SB_OUT_B1_O),
		.ready_in(SB_T0_NORTH_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T0_NORTH_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T0_NORTH_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T0_NORTH_SB_OUT_B1_valid_out),
		.S(SB_T0_NORTH_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T0_NORTH_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T0_SOUTH_SB_OUT_B1_I;
	assign MUX_SB_T0_SOUTH_SB_OUT_B1_I[5+:1] = MEM_output_width_1_num_2;
	assign MUX_SB_T0_SOUTH_SB_OUT_B1_I[4+:1] = MEM_output_width_1_num_1;
	assign MUX_SB_T0_SOUTH_SB_OUT_B1_I[3+:1] = MEM_output_width_1_num_0;
	assign MUX_SB_T0_SOUTH_SB_OUT_B1_I[2+:1] = WIRE_SB_T1_WEST_SB_IN_B1_O;
	assign MUX_SB_T0_SOUTH_SB_OUT_B1_I[1+:1] = WIRE_SB_T0_NORTH_SB_IN_B1_O;
	assign MUX_SB_T0_SOUTH_SB_OUT_B1_I[0+:1] = WIRE_SB_T3_EAST_SB_IN_B1_O;
	wire [5:0] MUX_SB_T0_SOUTH_SB_OUT_B1_valid_in;
	assign MUX_SB_T0_SOUTH_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid, MEM_output_width_1_num_1_valid, MEM_output_width_1_num_0_valid, WIRE_SB_T1_WEST_SB_IN_B1_valid_out, WIRE_SB_T0_NORTH_SB_IN_B1_valid_out, WIRE_SB_T3_EAST_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T0_SOUTH_SB_OUT_B1(
		.I(MUX_SB_T0_SOUTH_SB_OUT_B1_I),
		.O(MUX_SB_T0_SOUTH_SB_OUT_B1_O),
		.ready_in(SB_T0_SOUTH_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T0_SOUTH_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T0_SOUTH_SB_OUT_B1_valid_out),
		.S(SB_T0_SOUTH_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T0_WEST_SB_OUT_B1_I;
	assign MUX_SB_T0_WEST_SB_OUT_B1_I[5+:1] = MEM_output_width_1_num_2;
	assign MUX_SB_T0_WEST_SB_OUT_B1_I[4+:1] = MEM_output_width_1_num_1;
	assign MUX_SB_T0_WEST_SB_OUT_B1_I[3+:1] = MEM_output_width_1_num_0;
	assign MUX_SB_T0_WEST_SB_OUT_B1_I[2+:1] = WIRE_SB_T0_EAST_SB_IN_B1_O;
	assign MUX_SB_T0_WEST_SB_OUT_B1_I[1+:1] = WIRE_SB_T4_SOUTH_SB_IN_B1_O;
	assign MUX_SB_T0_WEST_SB_OUT_B1_I[0+:1] = WIRE_SB_T0_NORTH_SB_IN_B1_O;
	wire [5:0] MUX_SB_T0_WEST_SB_OUT_B1_valid_in;
	assign MUX_SB_T0_WEST_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid, MEM_output_width_1_num_1_valid, MEM_output_width_1_num_0_valid, WIRE_SB_T0_EAST_SB_IN_B1_valid_out, WIRE_SB_T4_SOUTH_SB_IN_B1_valid_out, WIRE_SB_T0_NORTH_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T0_WEST_SB_OUT_B1(
		.I(MUX_SB_T0_WEST_SB_OUT_B1_I),
		.O(MUX_SB_T0_WEST_SB_OUT_B1_O),
		.ready_in(SB_T0_WEST_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T0_WEST_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T0_WEST_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T0_WEST_SB_OUT_B1_valid_out),
		.S(SB_T0_WEST_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T0_WEST_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T1_EAST_SB_OUT_B1_I;
	assign MUX_SB_T1_EAST_SB_OUT_B1_I[5+:1] = MEM_output_width_1_num_2;
	assign MUX_SB_T1_EAST_SB_OUT_B1_I[4+:1] = MEM_output_width_1_num_1;
	assign MUX_SB_T1_EAST_SB_OUT_B1_I[3+:1] = MEM_output_width_1_num_0;
	assign MUX_SB_T1_EAST_SB_OUT_B1_I[2+:1] = WIRE_SB_T2_SOUTH_SB_IN_B1_O;
	assign MUX_SB_T1_EAST_SB_OUT_B1_I[1+:1] = WIRE_SB_T1_WEST_SB_IN_B1_O;
	assign MUX_SB_T1_EAST_SB_OUT_B1_I[0+:1] = WIRE_SB_T0_NORTH_SB_IN_B1_O;
	wire [5:0] MUX_SB_T1_EAST_SB_OUT_B1_valid_in;
	assign MUX_SB_T1_EAST_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid, MEM_output_width_1_num_1_valid, MEM_output_width_1_num_0_valid, WIRE_SB_T2_SOUTH_SB_IN_B1_valid_out, WIRE_SB_T1_WEST_SB_IN_B1_valid_out, WIRE_SB_T0_NORTH_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T1_EAST_SB_OUT_B1(
		.I(MUX_SB_T1_EAST_SB_OUT_B1_I),
		.O(MUX_SB_T1_EAST_SB_OUT_B1_O),
		.ready_in(SB_T1_EAST_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T1_EAST_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T1_EAST_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T1_EAST_SB_OUT_B1_valid_out),
		.S(SB_T1_EAST_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T1_EAST_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T1_NORTH_SB_OUT_B1_I;
	assign MUX_SB_T1_NORTH_SB_OUT_B1_I[5+:1] = MEM_output_width_1_num_2;
	assign MUX_SB_T1_NORTH_SB_OUT_B1_I[4+:1] = MEM_output_width_1_num_1;
	assign MUX_SB_T1_NORTH_SB_OUT_B1_I[3+:1] = MEM_output_width_1_num_0;
	assign MUX_SB_T1_NORTH_SB_OUT_B1_I[2+:1] = WIRE_SB_T4_WEST_SB_IN_B1_O;
	assign MUX_SB_T1_NORTH_SB_OUT_B1_I[1+:1] = WIRE_SB_T1_SOUTH_SB_IN_B1_O;
	assign MUX_SB_T1_NORTH_SB_OUT_B1_I[0+:1] = WIRE_SB_T2_EAST_SB_IN_B1_O;
	wire [5:0] MUX_SB_T1_NORTH_SB_OUT_B1_valid_in;
	assign MUX_SB_T1_NORTH_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid, MEM_output_width_1_num_1_valid, MEM_output_width_1_num_0_valid, WIRE_SB_T4_WEST_SB_IN_B1_valid_out, WIRE_SB_T1_SOUTH_SB_IN_B1_valid_out, WIRE_SB_T2_EAST_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T1_NORTH_SB_OUT_B1(
		.I(MUX_SB_T1_NORTH_SB_OUT_B1_I),
		.O(MUX_SB_T1_NORTH_SB_OUT_B1_O),
		.ready_in(SB_T1_NORTH_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T1_NORTH_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T1_NORTH_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T1_NORTH_SB_OUT_B1_valid_out),
		.S(SB_T1_NORTH_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T1_NORTH_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T1_SOUTH_SB_OUT_B1_I;
	assign MUX_SB_T1_SOUTH_SB_OUT_B1_I[5+:1] = MEM_output_width_1_num_2;
	assign MUX_SB_T1_SOUTH_SB_OUT_B1_I[4+:1] = MEM_output_width_1_num_1;
	assign MUX_SB_T1_SOUTH_SB_OUT_B1_I[3+:1] = MEM_output_width_1_num_0;
	assign MUX_SB_T1_SOUTH_SB_OUT_B1_I[2+:1] = WIRE_SB_T2_WEST_SB_IN_B1_O;
	assign MUX_SB_T1_SOUTH_SB_OUT_B1_I[1+:1] = WIRE_SB_T1_NORTH_SB_IN_B1_O;
	assign MUX_SB_T1_SOUTH_SB_OUT_B1_I[0+:1] = WIRE_SB_T2_EAST_SB_IN_B1_O;
	wire [5:0] MUX_SB_T1_SOUTH_SB_OUT_B1_valid_in;
	assign MUX_SB_T1_SOUTH_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid, MEM_output_width_1_num_1_valid, MEM_output_width_1_num_0_valid, WIRE_SB_T2_WEST_SB_IN_B1_valid_out, WIRE_SB_T1_NORTH_SB_IN_B1_valid_out, WIRE_SB_T2_EAST_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T1_SOUTH_SB_OUT_B1(
		.I(MUX_SB_T1_SOUTH_SB_OUT_B1_I),
		.O(MUX_SB_T1_SOUTH_SB_OUT_B1_O),
		.ready_in(SB_T1_SOUTH_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T1_SOUTH_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T1_SOUTH_SB_OUT_B1_valid_out),
		.S(SB_T1_SOUTH_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T1_WEST_SB_OUT_B1_I;
	assign MUX_SB_T1_WEST_SB_OUT_B1_I[5+:1] = MEM_output_width_1_num_2;
	assign MUX_SB_T1_WEST_SB_OUT_B1_I[4+:1] = MEM_output_width_1_num_1;
	assign MUX_SB_T1_WEST_SB_OUT_B1_I[3+:1] = MEM_output_width_1_num_0;
	assign MUX_SB_T1_WEST_SB_OUT_B1_I[2+:1] = WIRE_SB_T1_EAST_SB_IN_B1_O;
	assign MUX_SB_T1_WEST_SB_OUT_B1_I[1+:1] = WIRE_SB_T0_SOUTH_SB_IN_B1_O;
	assign MUX_SB_T1_WEST_SB_OUT_B1_I[0+:1] = WIRE_SB_T4_NORTH_SB_IN_B1_O;
	wire [5:0] MUX_SB_T1_WEST_SB_OUT_B1_valid_in;
	assign MUX_SB_T1_WEST_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid, MEM_output_width_1_num_1_valid, MEM_output_width_1_num_0_valid, WIRE_SB_T1_EAST_SB_IN_B1_valid_out, WIRE_SB_T0_SOUTH_SB_IN_B1_valid_out, WIRE_SB_T4_NORTH_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T1_WEST_SB_OUT_B1(
		.I(MUX_SB_T1_WEST_SB_OUT_B1_I),
		.O(MUX_SB_T1_WEST_SB_OUT_B1_O),
		.ready_in(SB_T1_WEST_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T1_WEST_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T1_WEST_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T1_WEST_SB_OUT_B1_valid_out),
		.S(SB_T1_WEST_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T1_WEST_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T2_EAST_SB_OUT_B1_I;
	assign MUX_SB_T2_EAST_SB_OUT_B1_I[5+:1] = MEM_output_width_1_num_2;
	assign MUX_SB_T2_EAST_SB_OUT_B1_I[4+:1] = MEM_output_width_1_num_1;
	assign MUX_SB_T2_EAST_SB_OUT_B1_I[3+:1] = MEM_output_width_1_num_0;
	assign MUX_SB_T2_EAST_SB_OUT_B1_I[2+:1] = WIRE_SB_T2_WEST_SB_IN_B1_O;
	assign MUX_SB_T2_EAST_SB_OUT_B1_I[1+:1] = WIRE_SB_T1_SOUTH_SB_IN_B1_O;
	assign MUX_SB_T2_EAST_SB_OUT_B1_I[0+:1] = WIRE_SB_T1_NORTH_SB_IN_B1_O;
	wire [5:0] MUX_SB_T2_EAST_SB_OUT_B1_valid_in;
	assign MUX_SB_T2_EAST_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid, MEM_output_width_1_num_1_valid, MEM_output_width_1_num_0_valid, WIRE_SB_T2_WEST_SB_IN_B1_valid_out, WIRE_SB_T1_SOUTH_SB_IN_B1_valid_out, WIRE_SB_T1_NORTH_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T2_EAST_SB_OUT_B1(
		.I(MUX_SB_T2_EAST_SB_OUT_B1_I),
		.O(MUX_SB_T2_EAST_SB_OUT_B1_O),
		.ready_in(SB_T2_EAST_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T2_EAST_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T2_EAST_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T2_EAST_SB_OUT_B1_valid_out),
		.S(SB_T2_EAST_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T2_EAST_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T2_NORTH_SB_OUT_B1_I;
	assign MUX_SB_T2_NORTH_SB_OUT_B1_I[5+:1] = MEM_output_width_1_num_2;
	assign MUX_SB_T2_NORTH_SB_OUT_B1_I[4+:1] = MEM_output_width_1_num_1;
	assign MUX_SB_T2_NORTH_SB_OUT_B1_I[3+:1] = MEM_output_width_1_num_0;
	assign MUX_SB_T2_NORTH_SB_OUT_B1_I[2+:1] = WIRE_SB_T3_WEST_SB_IN_B1_O;
	assign MUX_SB_T2_NORTH_SB_OUT_B1_I[1+:1] = WIRE_SB_T2_SOUTH_SB_IN_B1_O;
	assign MUX_SB_T2_NORTH_SB_OUT_B1_I[0+:1] = WIRE_SB_T3_EAST_SB_IN_B1_O;
	wire [5:0] MUX_SB_T2_NORTH_SB_OUT_B1_valid_in;
	assign MUX_SB_T2_NORTH_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid, MEM_output_width_1_num_1_valid, MEM_output_width_1_num_0_valid, WIRE_SB_T3_WEST_SB_IN_B1_valid_out, WIRE_SB_T2_SOUTH_SB_IN_B1_valid_out, WIRE_SB_T3_EAST_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T2_NORTH_SB_OUT_B1(
		.I(MUX_SB_T2_NORTH_SB_OUT_B1_I),
		.O(MUX_SB_T2_NORTH_SB_OUT_B1_O),
		.ready_in(SB_T2_NORTH_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T2_NORTH_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T2_NORTH_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T2_NORTH_SB_OUT_B1_valid_out),
		.S(SB_T2_NORTH_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T2_NORTH_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T2_SOUTH_SB_OUT_B1_I;
	assign MUX_SB_T2_SOUTH_SB_OUT_B1_I[5+:1] = MEM_output_width_1_num_2;
	assign MUX_SB_T2_SOUTH_SB_OUT_B1_I[4+:1] = MEM_output_width_1_num_1;
	assign MUX_SB_T2_SOUTH_SB_OUT_B1_I[3+:1] = MEM_output_width_1_num_0;
	assign MUX_SB_T2_SOUTH_SB_OUT_B1_I[2+:1] = WIRE_SB_T3_WEST_SB_IN_B1_O;
	assign MUX_SB_T2_SOUTH_SB_OUT_B1_I[1+:1] = WIRE_SB_T2_NORTH_SB_IN_B1_O;
	assign MUX_SB_T2_SOUTH_SB_OUT_B1_I[0+:1] = WIRE_SB_T1_EAST_SB_IN_B1_O;
	wire [5:0] MUX_SB_T2_SOUTH_SB_OUT_B1_valid_in;
	assign MUX_SB_T2_SOUTH_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid, MEM_output_width_1_num_1_valid, MEM_output_width_1_num_0_valid, WIRE_SB_T3_WEST_SB_IN_B1_valid_out, WIRE_SB_T2_NORTH_SB_IN_B1_valid_out, WIRE_SB_T1_EAST_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T2_SOUTH_SB_OUT_B1(
		.I(MUX_SB_T2_SOUTH_SB_OUT_B1_I),
		.O(MUX_SB_T2_SOUTH_SB_OUT_B1_O),
		.ready_in(SB_T2_SOUTH_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T2_SOUTH_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T2_SOUTH_SB_OUT_B1_valid_out),
		.S(SB_T2_SOUTH_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T2_WEST_SB_OUT_B1_I;
	assign MUX_SB_T2_WEST_SB_OUT_B1_I[5+:1] = MEM_output_width_1_num_2;
	assign MUX_SB_T2_WEST_SB_OUT_B1_I[4+:1] = MEM_output_width_1_num_1;
	assign MUX_SB_T2_WEST_SB_OUT_B1_I[3+:1] = MEM_output_width_1_num_0;
	assign MUX_SB_T2_WEST_SB_OUT_B1_I[2+:1] = WIRE_SB_T2_EAST_SB_IN_B1_O;
	assign MUX_SB_T2_WEST_SB_OUT_B1_I[1+:1] = WIRE_SB_T1_SOUTH_SB_IN_B1_O;
	assign MUX_SB_T2_WEST_SB_OUT_B1_I[0+:1] = WIRE_SB_T3_NORTH_SB_IN_B1_O;
	wire [5:0] MUX_SB_T2_WEST_SB_OUT_B1_valid_in;
	assign MUX_SB_T2_WEST_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid, MEM_output_width_1_num_1_valid, MEM_output_width_1_num_0_valid, WIRE_SB_T2_EAST_SB_IN_B1_valid_out, WIRE_SB_T1_SOUTH_SB_IN_B1_valid_out, WIRE_SB_T3_NORTH_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T2_WEST_SB_OUT_B1(
		.I(MUX_SB_T2_WEST_SB_OUT_B1_I),
		.O(MUX_SB_T2_WEST_SB_OUT_B1_O),
		.ready_in(SB_T2_WEST_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T2_WEST_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T2_WEST_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T2_WEST_SB_OUT_B1_valid_out),
		.S(SB_T2_WEST_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T2_WEST_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T3_EAST_SB_OUT_B1_I;
	assign MUX_SB_T3_EAST_SB_OUT_B1_I[5+:1] = MEM_output_width_1_num_2;
	assign MUX_SB_T3_EAST_SB_OUT_B1_I[4+:1] = MEM_output_width_1_num_1;
	assign MUX_SB_T3_EAST_SB_OUT_B1_I[3+:1] = MEM_output_width_1_num_0;
	assign MUX_SB_T3_EAST_SB_OUT_B1_I[2+:1] = WIRE_SB_T3_WEST_SB_IN_B1_O;
	assign MUX_SB_T3_EAST_SB_OUT_B1_I[1+:1] = WIRE_SB_T2_NORTH_SB_IN_B1_O;
	assign MUX_SB_T3_EAST_SB_OUT_B1_I[0+:1] = WIRE_SB_T0_SOUTH_SB_IN_B1_O;
	wire [5:0] MUX_SB_T3_EAST_SB_OUT_B1_valid_in;
	assign MUX_SB_T3_EAST_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid, MEM_output_width_1_num_1_valid, MEM_output_width_1_num_0_valid, WIRE_SB_T3_WEST_SB_IN_B1_valid_out, WIRE_SB_T2_NORTH_SB_IN_B1_valid_out, WIRE_SB_T0_SOUTH_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T3_EAST_SB_OUT_B1(
		.I(MUX_SB_T3_EAST_SB_OUT_B1_I),
		.O(MUX_SB_T3_EAST_SB_OUT_B1_O),
		.ready_in(SB_T3_EAST_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T3_EAST_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T3_EAST_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T3_EAST_SB_OUT_B1_valid_out),
		.S(SB_T3_EAST_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T3_EAST_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T3_NORTH_SB_OUT_B1_I;
	assign MUX_SB_T3_NORTH_SB_OUT_B1_I[5+:1] = MEM_output_width_1_num_2;
	assign MUX_SB_T3_NORTH_SB_OUT_B1_I[4+:1] = MEM_output_width_1_num_1;
	assign MUX_SB_T3_NORTH_SB_OUT_B1_I[3+:1] = MEM_output_width_1_num_0;
	assign MUX_SB_T3_NORTH_SB_OUT_B1_I[2+:1] = WIRE_SB_T3_SOUTH_SB_IN_B1_O;
	assign MUX_SB_T3_NORTH_SB_OUT_B1_I[1+:1] = WIRE_SB_T4_EAST_SB_IN_B1_O;
	assign MUX_SB_T3_NORTH_SB_OUT_B1_I[0+:1] = WIRE_SB_T2_WEST_SB_IN_B1_O;
	wire [5:0] MUX_SB_T3_NORTH_SB_OUT_B1_valid_in;
	assign MUX_SB_T3_NORTH_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid, MEM_output_width_1_num_1_valid, MEM_output_width_1_num_0_valid, WIRE_SB_T3_SOUTH_SB_IN_B1_valid_out, WIRE_SB_T4_EAST_SB_IN_B1_valid_out, WIRE_SB_T2_WEST_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T3_NORTH_SB_OUT_B1(
		.I(MUX_SB_T3_NORTH_SB_OUT_B1_I),
		.O(MUX_SB_T3_NORTH_SB_OUT_B1_O),
		.ready_in(SB_T3_NORTH_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T3_NORTH_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T3_NORTH_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T3_NORTH_SB_OUT_B1_valid_out),
		.S(SB_T3_NORTH_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T3_NORTH_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T3_SOUTH_SB_OUT_B1_I;
	assign MUX_SB_T3_SOUTH_SB_OUT_B1_I[5+:1] = MEM_output_width_1_num_2;
	assign MUX_SB_T3_SOUTH_SB_OUT_B1_I[4+:1] = MEM_output_width_1_num_1;
	assign MUX_SB_T3_SOUTH_SB_OUT_B1_I[3+:1] = MEM_output_width_1_num_0;
	assign MUX_SB_T3_SOUTH_SB_OUT_B1_I[2+:1] = WIRE_SB_T4_WEST_SB_IN_B1_O;
	assign MUX_SB_T3_SOUTH_SB_OUT_B1_I[1+:1] = WIRE_SB_T3_NORTH_SB_IN_B1_O;
	assign MUX_SB_T3_SOUTH_SB_OUT_B1_I[0+:1] = WIRE_SB_T0_EAST_SB_IN_B1_O;
	wire [5:0] MUX_SB_T3_SOUTH_SB_OUT_B1_valid_in;
	assign MUX_SB_T3_SOUTH_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid, MEM_output_width_1_num_1_valid, MEM_output_width_1_num_0_valid, WIRE_SB_T4_WEST_SB_IN_B1_valid_out, WIRE_SB_T3_NORTH_SB_IN_B1_valid_out, WIRE_SB_T0_EAST_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T3_SOUTH_SB_OUT_B1(
		.I(MUX_SB_T3_SOUTH_SB_OUT_B1_I),
		.O(MUX_SB_T3_SOUTH_SB_OUT_B1_O),
		.ready_in(SB_T3_SOUTH_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T3_SOUTH_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T3_SOUTH_SB_OUT_B1_valid_out),
		.S(SB_T3_SOUTH_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T3_WEST_SB_OUT_B1_I;
	assign MUX_SB_T3_WEST_SB_OUT_B1_I[5+:1] = MEM_output_width_1_num_2;
	assign MUX_SB_T3_WEST_SB_OUT_B1_I[4+:1] = MEM_output_width_1_num_1;
	assign MUX_SB_T3_WEST_SB_OUT_B1_I[3+:1] = MEM_output_width_1_num_0;
	assign MUX_SB_T3_WEST_SB_OUT_B1_I[2+:1] = WIRE_SB_T3_EAST_SB_IN_B1_O;
	assign MUX_SB_T3_WEST_SB_OUT_B1_I[1+:1] = WIRE_SB_T2_SOUTH_SB_IN_B1_O;
	assign MUX_SB_T3_WEST_SB_OUT_B1_I[0+:1] = WIRE_SB_T2_NORTH_SB_IN_B1_O;
	wire [5:0] MUX_SB_T3_WEST_SB_OUT_B1_valid_in;
	assign MUX_SB_T3_WEST_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid, MEM_output_width_1_num_1_valid, MEM_output_width_1_num_0_valid, WIRE_SB_T3_EAST_SB_IN_B1_valid_out, WIRE_SB_T2_SOUTH_SB_IN_B1_valid_out, WIRE_SB_T2_NORTH_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T3_WEST_SB_OUT_B1(
		.I(MUX_SB_T3_WEST_SB_OUT_B1_I),
		.O(MUX_SB_T3_WEST_SB_OUT_B1_O),
		.ready_in(SB_T3_WEST_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T3_WEST_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T3_WEST_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T3_WEST_SB_OUT_B1_valid_out),
		.S(SB_T3_WEST_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T3_WEST_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T4_EAST_SB_OUT_B1_I;
	assign MUX_SB_T4_EAST_SB_OUT_B1_I[5+:1] = MEM_output_width_1_num_2;
	assign MUX_SB_T4_EAST_SB_OUT_B1_I[4+:1] = MEM_output_width_1_num_1;
	assign MUX_SB_T4_EAST_SB_OUT_B1_I[3+:1] = MEM_output_width_1_num_0;
	assign MUX_SB_T4_EAST_SB_OUT_B1_I[2+:1] = WIRE_SB_T4_WEST_SB_IN_B1_O;
	assign MUX_SB_T4_EAST_SB_OUT_B1_I[1+:1] = WIRE_SB_T4_SOUTH_SB_IN_B1_O;
	assign MUX_SB_T4_EAST_SB_OUT_B1_I[0+:1] = WIRE_SB_T3_NORTH_SB_IN_B1_O;
	wire [5:0] MUX_SB_T4_EAST_SB_OUT_B1_valid_in;
	assign MUX_SB_T4_EAST_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid, MEM_output_width_1_num_1_valid, MEM_output_width_1_num_0_valid, WIRE_SB_T4_WEST_SB_IN_B1_valid_out, WIRE_SB_T4_SOUTH_SB_IN_B1_valid_out, WIRE_SB_T3_NORTH_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T4_EAST_SB_OUT_B1(
		.I(MUX_SB_T4_EAST_SB_OUT_B1_I),
		.O(MUX_SB_T4_EAST_SB_OUT_B1_O),
		.ready_in(SB_T4_EAST_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T4_EAST_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T4_EAST_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T4_EAST_SB_OUT_B1_valid_out),
		.S(SB_T4_EAST_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T4_EAST_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T4_NORTH_SB_OUT_B1_I;
	assign MUX_SB_T4_NORTH_SB_OUT_B1_I[5+:1] = MEM_output_width_1_num_2;
	assign MUX_SB_T4_NORTH_SB_OUT_B1_I[4+:1] = MEM_output_width_1_num_1;
	assign MUX_SB_T4_NORTH_SB_OUT_B1_I[3+:1] = MEM_output_width_1_num_0;
	assign MUX_SB_T4_NORTH_SB_OUT_B1_I[2+:1] = WIRE_SB_T4_SOUTH_SB_IN_B1_O;
	assign MUX_SB_T4_NORTH_SB_OUT_B1_I[1+:1] = WIRE_SB_T0_EAST_SB_IN_B1_O;
	assign MUX_SB_T4_NORTH_SB_OUT_B1_I[0+:1] = WIRE_SB_T1_WEST_SB_IN_B1_O;
	wire [5:0] MUX_SB_T4_NORTH_SB_OUT_B1_valid_in;
	assign MUX_SB_T4_NORTH_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid, MEM_output_width_1_num_1_valid, MEM_output_width_1_num_0_valid, WIRE_SB_T4_SOUTH_SB_IN_B1_valid_out, WIRE_SB_T0_EAST_SB_IN_B1_valid_out, WIRE_SB_T1_WEST_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T4_NORTH_SB_OUT_B1(
		.I(MUX_SB_T4_NORTH_SB_OUT_B1_I),
		.O(MUX_SB_T4_NORTH_SB_OUT_B1_O),
		.ready_in(SB_T4_NORTH_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T4_NORTH_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T4_NORTH_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T4_NORTH_SB_OUT_B1_valid_out),
		.S(SB_T4_NORTH_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T4_NORTH_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T4_SOUTH_SB_OUT_B1_I;
	assign MUX_SB_T4_SOUTH_SB_OUT_B1_I[5+:1] = MEM_output_width_1_num_2;
	assign MUX_SB_T4_SOUTH_SB_OUT_B1_I[4+:1] = MEM_output_width_1_num_1;
	assign MUX_SB_T4_SOUTH_SB_OUT_B1_I[3+:1] = MEM_output_width_1_num_0;
	assign MUX_SB_T4_SOUTH_SB_OUT_B1_I[2+:1] = WIRE_SB_T4_NORTH_SB_IN_B1_O;
	assign MUX_SB_T4_SOUTH_SB_OUT_B1_I[1+:1] = WIRE_SB_T4_EAST_SB_IN_B1_O;
	assign MUX_SB_T4_SOUTH_SB_OUT_B1_I[0+:1] = WIRE_SB_T0_WEST_SB_IN_B1_O;
	wire [5:0] MUX_SB_T4_SOUTH_SB_OUT_B1_valid_in;
	assign MUX_SB_T4_SOUTH_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid, MEM_output_width_1_num_1_valid, MEM_output_width_1_num_0_valid, WIRE_SB_T4_NORTH_SB_IN_B1_valid_out, WIRE_SB_T4_EAST_SB_IN_B1_valid_out, WIRE_SB_T0_WEST_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T4_SOUTH_SB_OUT_B1(
		.I(MUX_SB_T4_SOUTH_SB_OUT_B1_I),
		.O(MUX_SB_T4_SOUTH_SB_OUT_B1_O),
		.ready_in(SB_T4_SOUTH_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T4_SOUTH_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T4_SOUTH_SB_OUT_B1_valid_out),
		.S(SB_T4_SOUTH_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel)
	);
	wire [5:0] MUX_SB_T4_WEST_SB_OUT_B1_I;
	assign MUX_SB_T4_WEST_SB_OUT_B1_I[5+:1] = MEM_output_width_1_num_2;
	assign MUX_SB_T4_WEST_SB_OUT_B1_I[4+:1] = MEM_output_width_1_num_1;
	assign MUX_SB_T4_WEST_SB_OUT_B1_I[3+:1] = MEM_output_width_1_num_0;
	assign MUX_SB_T4_WEST_SB_OUT_B1_I[2+:1] = WIRE_SB_T4_EAST_SB_IN_B1_O;
	assign MUX_SB_T4_WEST_SB_OUT_B1_I[1+:1] = WIRE_SB_T3_SOUTH_SB_IN_B1_O;
	assign MUX_SB_T4_WEST_SB_OUT_B1_I[0+:1] = WIRE_SB_T1_NORTH_SB_IN_B1_O;
	wire [5:0] MUX_SB_T4_WEST_SB_OUT_B1_valid_in;
	assign MUX_SB_T4_WEST_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid, MEM_output_width_1_num_1_valid, MEM_output_width_1_num_0_valid, WIRE_SB_T4_EAST_SB_IN_B1_valid_out, WIRE_SB_T3_SOUTH_SB_IN_B1_valid_out, WIRE_SB_T1_NORTH_SB_IN_B1_valid_out};
	mux_aoi_ready_valid_6_1 MUX_SB_T4_WEST_SB_OUT_B1(
		.I(MUX_SB_T4_WEST_SB_OUT_B1_I),
		.O(MUX_SB_T4_WEST_SB_OUT_B1_O),
		.ready_in(SB_T4_WEST_SB_OUT_B1_FANOUT_O[0]),
		.ready_out(MUX_SB_T4_WEST_SB_OUT_B1_ready_out),
		.valid_in(MUX_SB_T4_WEST_SB_OUT_B1_valid_in),
		.valid_out(MUX_SB_T4_WEST_SB_OUT_B1_valid_out),
		.S(SB_T4_WEST_SB_OUT_B1_sel_value_O),
		.out_sel(MUX_SB_T4_WEST_SB_OUT_B1_out_sel)
	);
	SplitFifo_1 REG_T0_EAST_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T0_EAST_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T0_EAST_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T0_EAST_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T0_EAST_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst2_out[0]),
		.end_fifo(REG_T0_EAST_B1_end_value_O[0]),
		.valid0(MUX_SB_T0_EAST_SB_OUT_B1_valid_out),
		.valid1(REG_T0_EAST_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T0_EAST_B1_ready_out),
		.fifo_en(REG_T0_EAST_B1_fifo_value_O[0])
	);
	SliceWrapper_32_0_1 REG_T0_EAST_B1_end_value(
		.I(config_reg_0_O),
		.O(REG_T0_EAST_B1_end_value_O)
	);
	SliceWrapper_32_1_2 REG_T0_EAST_B1_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T0_EAST_B1_fifo_value_O)
	);
	SliceWrapper_32_2_3 REG_T0_EAST_B1_start_value(
		.I(config_reg_0_O),
		.O(REG_T0_EAST_B1_start_value_O)
	);
	SplitFifo_1 REG_T0_NORTH_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T0_NORTH_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T0_NORTH_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T0_NORTH_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T0_NORTH_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst0_out[0]),
		.end_fifo(REG_T0_NORTH_B1_end_value_O[0]),
		.valid0(MUX_SB_T0_NORTH_SB_OUT_B1_valid_out),
		.valid1(REG_T0_NORTH_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T0_NORTH_B1_ready_out),
		.fifo_en(REG_T0_NORTH_B1_fifo_value_O[0])
	);
	SliceWrapper_32_3_4 REG_T0_NORTH_B1_end_value(
		.I(config_reg_0_O),
		.O(REG_T0_NORTH_B1_end_value_O)
	);
	SliceWrapper_32_4_5 REG_T0_NORTH_B1_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T0_NORTH_B1_fifo_value_O)
	);
	SliceWrapper_32_5_6 REG_T0_NORTH_B1_start_value(
		.I(config_reg_0_O),
		.O(REG_T0_NORTH_B1_start_value_O)
	);
	SplitFifo_1 REG_T0_SOUTH_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T0_SOUTH_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T0_SOUTH_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T0_SOUTH_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T0_SOUTH_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst1_out[0]),
		.end_fifo(REG_T0_SOUTH_B1_end_value_O[0]),
		.valid0(MUX_SB_T0_SOUTH_SB_OUT_B1_valid_out),
		.valid1(REG_T0_SOUTH_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T0_SOUTH_B1_ready_out),
		.fifo_en(REG_T0_SOUTH_B1_fifo_value_O[0])
	);
	SliceWrapper_32_6_7 REG_T0_SOUTH_B1_end_value(
		.I(config_reg_0_O),
		.O(REG_T0_SOUTH_B1_end_value_O)
	);
	SliceWrapper_32_7_8 REG_T0_SOUTH_B1_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T0_SOUTH_B1_fifo_value_O)
	);
	SliceWrapper_32_8_9 REG_T0_SOUTH_B1_start_value(
		.I(config_reg_0_O),
		.O(REG_T0_SOUTH_B1_start_value_O)
	);
	SplitFifo_1 REG_T0_WEST_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T0_WEST_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T0_WEST_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T0_WEST_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T0_WEST_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst3_out[0]),
		.end_fifo(REG_T0_WEST_B1_end_value_O[0]),
		.valid0(MUX_SB_T0_WEST_SB_OUT_B1_valid_out),
		.valid1(REG_T0_WEST_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T0_WEST_B1_ready_out),
		.fifo_en(REG_T0_WEST_B1_fifo_value_O[0])
	);
	SliceWrapper_32_9_10 REG_T0_WEST_B1_end_value(
		.I(config_reg_0_O),
		.O(REG_T0_WEST_B1_end_value_O)
	);
	SliceWrapper_32_10_11 REG_T0_WEST_B1_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T0_WEST_B1_fifo_value_O)
	);
	SliceWrapper_32_11_12 REG_T0_WEST_B1_start_value(
		.I(config_reg_0_O),
		.O(REG_T0_WEST_B1_start_value_O)
	);
	SplitFifo_1 REG_T1_EAST_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T1_EAST_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T1_EAST_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T1_EAST_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T1_EAST_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst6_out[0]),
		.end_fifo(REG_T1_EAST_B1_end_value_O[0]),
		.valid0(MUX_SB_T1_EAST_SB_OUT_B1_valid_out),
		.valid1(REG_T1_EAST_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T1_EAST_B1_ready_out),
		.fifo_en(REG_T1_EAST_B1_fifo_value_O[0])
	);
	SliceWrapper_32_12_13 REG_T1_EAST_B1_end_value(
		.I(config_reg_0_O),
		.O(REG_T1_EAST_B1_end_value_O)
	);
	SliceWrapper_32_13_14 REG_T1_EAST_B1_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T1_EAST_B1_fifo_value_O)
	);
	SliceWrapper_32_14_15 REG_T1_EAST_B1_start_value(
		.I(config_reg_0_O),
		.O(REG_T1_EAST_B1_start_value_O)
	);
	SplitFifo_1 REG_T1_NORTH_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T1_NORTH_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T1_NORTH_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T1_NORTH_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T1_NORTH_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst4_out[0]),
		.end_fifo(REG_T1_NORTH_B1_end_value_O[0]),
		.valid0(MUX_SB_T1_NORTH_SB_OUT_B1_valid_out),
		.valid1(REG_T1_NORTH_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T1_NORTH_B1_ready_out),
		.fifo_en(REG_T1_NORTH_B1_fifo_value_O[0])
	);
	SliceWrapper_32_15_16 REG_T1_NORTH_B1_end_value(
		.I(config_reg_0_O),
		.O(REG_T1_NORTH_B1_end_value_O)
	);
	SliceWrapper_32_16_17 REG_T1_NORTH_B1_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T1_NORTH_B1_fifo_value_O)
	);
	SliceWrapper_32_17_18 REG_T1_NORTH_B1_start_value(
		.I(config_reg_0_O),
		.O(REG_T1_NORTH_B1_start_value_O)
	);
	SplitFifo_1 REG_T1_SOUTH_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T1_SOUTH_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T1_SOUTH_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T1_SOUTH_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T1_SOUTH_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst5_out[0]),
		.end_fifo(REG_T1_SOUTH_B1_end_value_O[0]),
		.valid0(MUX_SB_T1_SOUTH_SB_OUT_B1_valid_out),
		.valid1(REG_T1_SOUTH_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T1_SOUTH_B1_ready_out),
		.fifo_en(REG_T1_SOUTH_B1_fifo_value_O[0])
	);
	SliceWrapper_32_18_19 REG_T1_SOUTH_B1_end_value(
		.I(config_reg_0_O),
		.O(REG_T1_SOUTH_B1_end_value_O)
	);
	SliceWrapper_32_19_20 REG_T1_SOUTH_B1_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T1_SOUTH_B1_fifo_value_O)
	);
	SliceWrapper_32_20_21 REG_T1_SOUTH_B1_start_value(
		.I(config_reg_0_O),
		.O(REG_T1_SOUTH_B1_start_value_O)
	);
	SplitFifo_1 REG_T1_WEST_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T1_WEST_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T1_WEST_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T1_WEST_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T1_WEST_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst7_out[0]),
		.end_fifo(REG_T1_WEST_B1_end_value_O[0]),
		.valid0(MUX_SB_T1_WEST_SB_OUT_B1_valid_out),
		.valid1(REG_T1_WEST_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T1_WEST_B1_ready_out),
		.fifo_en(REG_T1_WEST_B1_fifo_value_O[0])
	);
	SliceWrapper_32_21_22 REG_T1_WEST_B1_end_value(
		.I(config_reg_0_O),
		.O(REG_T1_WEST_B1_end_value_O)
	);
	SliceWrapper_32_22_23 REG_T1_WEST_B1_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T1_WEST_B1_fifo_value_O)
	);
	SliceWrapper_32_23_24 REG_T1_WEST_B1_start_value(
		.I(config_reg_0_O),
		.O(REG_T1_WEST_B1_start_value_O)
	);
	SplitFifo_1 REG_T2_EAST_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T2_EAST_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T2_EAST_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T2_EAST_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T2_EAST_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst10_out[0]),
		.end_fifo(REG_T2_EAST_B1_end_value_O[0]),
		.valid0(MUX_SB_T2_EAST_SB_OUT_B1_valid_out),
		.valid1(REG_T2_EAST_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T2_EAST_B1_ready_out),
		.fifo_en(REG_T2_EAST_B1_fifo_value_O[0])
	);
	SliceWrapper_32_24_25 REG_T2_EAST_B1_end_value(
		.I(config_reg_0_O),
		.O(REG_T2_EAST_B1_end_value_O)
	);
	SliceWrapper_32_25_26 REG_T2_EAST_B1_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T2_EAST_B1_fifo_value_O)
	);
	SliceWrapper_32_26_27 REG_T2_EAST_B1_start_value(
		.I(config_reg_0_O),
		.O(REG_T2_EAST_B1_start_value_O)
	);
	SplitFifo_1 REG_T2_NORTH_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T2_NORTH_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T2_NORTH_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T2_NORTH_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T2_NORTH_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst8_out[0]),
		.end_fifo(REG_T2_NORTH_B1_end_value_O[0]),
		.valid0(MUX_SB_T2_NORTH_SB_OUT_B1_valid_out),
		.valid1(REG_T2_NORTH_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T2_NORTH_B1_ready_out),
		.fifo_en(REG_T2_NORTH_B1_fifo_value_O[0])
	);
	SliceWrapper_32_27_28 REG_T2_NORTH_B1_end_value(
		.I(config_reg_0_O),
		.O(REG_T2_NORTH_B1_end_value_O)
	);
	SliceWrapper_32_28_29 REG_T2_NORTH_B1_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T2_NORTH_B1_fifo_value_O)
	);
	SliceWrapper_32_29_30 REG_T2_NORTH_B1_start_value(
		.I(config_reg_0_O),
		.O(REG_T2_NORTH_B1_start_value_O)
	);
	SplitFifo_1 REG_T2_SOUTH_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T2_SOUTH_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T2_SOUTH_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T2_SOUTH_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T2_SOUTH_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst9_out[0]),
		.end_fifo(REG_T2_SOUTH_B1_end_value_O[0]),
		.valid0(MUX_SB_T2_SOUTH_SB_OUT_B1_valid_out),
		.valid1(REG_T2_SOUTH_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T2_SOUTH_B1_ready_out),
		.fifo_en(REG_T2_SOUTH_B1_fifo_value_O[0])
	);
	SliceWrapper_32_30_31 REG_T2_SOUTH_B1_end_value(
		.I(config_reg_0_O),
		.O(REG_T2_SOUTH_B1_end_value_O)
	);
	SliceWrapper_32_31_32 REG_T2_SOUTH_B1_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T2_SOUTH_B1_fifo_value_O)
	);
	SliceWrapper_32_0_1 REG_T2_SOUTH_B1_start_value(
		.I(config_reg_1_O),
		.O(REG_T2_SOUTH_B1_start_value_O)
	);
	SplitFifo_1 REG_T2_WEST_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T2_WEST_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T2_WEST_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T2_WEST_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T2_WEST_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst11_out[0]),
		.end_fifo(REG_T2_WEST_B1_end_value_O[0]),
		.valid0(MUX_SB_T2_WEST_SB_OUT_B1_valid_out),
		.valid1(REG_T2_WEST_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T2_WEST_B1_ready_out),
		.fifo_en(REG_T2_WEST_B1_fifo_value_O[0])
	);
	SliceWrapper_32_1_2 REG_T2_WEST_B1_end_value(
		.I(config_reg_1_O),
		.O(REG_T2_WEST_B1_end_value_O)
	);
	SliceWrapper_32_2_3 REG_T2_WEST_B1_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T2_WEST_B1_fifo_value_O)
	);
	SliceWrapper_32_3_4 REG_T2_WEST_B1_start_value(
		.I(config_reg_1_O),
		.O(REG_T2_WEST_B1_start_value_O)
	);
	SplitFifo_1 REG_T3_EAST_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T3_EAST_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T3_EAST_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T3_EAST_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T3_EAST_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst14_out[0]),
		.end_fifo(REG_T3_EAST_B1_end_value_O[0]),
		.valid0(MUX_SB_T3_EAST_SB_OUT_B1_valid_out),
		.valid1(REG_T3_EAST_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T3_EAST_B1_ready_out),
		.fifo_en(REG_T3_EAST_B1_fifo_value_O[0])
	);
	SliceWrapper_32_4_5 REG_T3_EAST_B1_end_value(
		.I(config_reg_1_O),
		.O(REG_T3_EAST_B1_end_value_O)
	);
	SliceWrapper_32_5_6 REG_T3_EAST_B1_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T3_EAST_B1_fifo_value_O)
	);
	SliceWrapper_32_6_7 REG_T3_EAST_B1_start_value(
		.I(config_reg_1_O),
		.O(REG_T3_EAST_B1_start_value_O)
	);
	SplitFifo_1 REG_T3_NORTH_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T3_NORTH_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T3_NORTH_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T3_NORTH_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T3_NORTH_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst12_out[0]),
		.end_fifo(REG_T3_NORTH_B1_end_value_O[0]),
		.valid0(MUX_SB_T3_NORTH_SB_OUT_B1_valid_out),
		.valid1(REG_T3_NORTH_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T3_NORTH_B1_ready_out),
		.fifo_en(REG_T3_NORTH_B1_fifo_value_O[0])
	);
	SliceWrapper_32_7_8 REG_T3_NORTH_B1_end_value(
		.I(config_reg_1_O),
		.O(REG_T3_NORTH_B1_end_value_O)
	);
	SliceWrapper_32_8_9 REG_T3_NORTH_B1_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T3_NORTH_B1_fifo_value_O)
	);
	SliceWrapper_32_9_10 REG_T3_NORTH_B1_start_value(
		.I(config_reg_1_O),
		.O(REG_T3_NORTH_B1_start_value_O)
	);
	SplitFifo_1 REG_T3_SOUTH_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T3_SOUTH_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T3_SOUTH_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T3_SOUTH_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T3_SOUTH_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst13_out[0]),
		.end_fifo(REG_T3_SOUTH_B1_end_value_O[0]),
		.valid0(MUX_SB_T3_SOUTH_SB_OUT_B1_valid_out),
		.valid1(REG_T3_SOUTH_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T3_SOUTH_B1_ready_out),
		.fifo_en(REG_T3_SOUTH_B1_fifo_value_O[0])
	);
	SliceWrapper_32_10_11 REG_T3_SOUTH_B1_end_value(
		.I(config_reg_1_O),
		.O(REG_T3_SOUTH_B1_end_value_O)
	);
	SliceWrapper_32_11_12 REG_T3_SOUTH_B1_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T3_SOUTH_B1_fifo_value_O)
	);
	SliceWrapper_32_12_13 REG_T3_SOUTH_B1_start_value(
		.I(config_reg_1_O),
		.O(REG_T3_SOUTH_B1_start_value_O)
	);
	SplitFifo_1 REG_T3_WEST_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T3_WEST_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T3_WEST_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T3_WEST_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T3_WEST_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst15_out[0]),
		.end_fifo(REG_T3_WEST_B1_end_value_O[0]),
		.valid0(MUX_SB_T3_WEST_SB_OUT_B1_valid_out),
		.valid1(REG_T3_WEST_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T3_WEST_B1_ready_out),
		.fifo_en(REG_T3_WEST_B1_fifo_value_O[0])
	);
	SliceWrapper_32_13_14 REG_T3_WEST_B1_end_value(
		.I(config_reg_1_O),
		.O(REG_T3_WEST_B1_end_value_O)
	);
	SliceWrapper_32_14_15 REG_T3_WEST_B1_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T3_WEST_B1_fifo_value_O)
	);
	SliceWrapper_32_15_16 REG_T3_WEST_B1_start_value(
		.I(config_reg_1_O),
		.O(REG_T3_WEST_B1_start_value_O)
	);
	SplitFifo_1 REG_T4_EAST_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T4_EAST_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T4_EAST_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T4_EAST_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T4_EAST_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst18_out[0]),
		.end_fifo(REG_T4_EAST_B1_end_value_O[0]),
		.valid0(MUX_SB_T4_EAST_SB_OUT_B1_valid_out),
		.valid1(REG_T4_EAST_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T4_EAST_B1_ready_out),
		.fifo_en(REG_T4_EAST_B1_fifo_value_O[0])
	);
	SliceWrapper_32_16_17 REG_T4_EAST_B1_end_value(
		.I(config_reg_1_O),
		.O(REG_T4_EAST_B1_end_value_O)
	);
	SliceWrapper_32_17_18 REG_T4_EAST_B1_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T4_EAST_B1_fifo_value_O)
	);
	SliceWrapper_32_18_19 REG_T4_EAST_B1_start_value(
		.I(config_reg_1_O),
		.O(REG_T4_EAST_B1_start_value_O)
	);
	SplitFifo_1 REG_T4_NORTH_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T4_NORTH_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T4_NORTH_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T4_NORTH_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T4_NORTH_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst16_out[0]),
		.end_fifo(REG_T4_NORTH_B1_end_value_O[0]),
		.valid0(MUX_SB_T4_NORTH_SB_OUT_B1_valid_out),
		.valid1(REG_T4_NORTH_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T4_NORTH_B1_ready_out),
		.fifo_en(REG_T4_NORTH_B1_fifo_value_O[0])
	);
	SliceWrapper_32_19_20 REG_T4_NORTH_B1_end_value(
		.I(config_reg_1_O),
		.O(REG_T4_NORTH_B1_end_value_O)
	);
	SliceWrapper_32_20_21 REG_T4_NORTH_B1_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T4_NORTH_B1_fifo_value_O)
	);
	SliceWrapper_32_21_22 REG_T4_NORTH_B1_start_value(
		.I(config_reg_1_O),
		.O(REG_T4_NORTH_B1_start_value_O)
	);
	SplitFifo_1 REG_T4_SOUTH_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T4_SOUTH_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T4_SOUTH_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T4_SOUTH_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T4_SOUTH_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst17_out[0]),
		.end_fifo(REG_T4_SOUTH_B1_end_value_O[0]),
		.valid0(MUX_SB_T4_SOUTH_SB_OUT_B1_valid_out),
		.valid1(REG_T4_SOUTH_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T4_SOUTH_B1_ready_out),
		.fifo_en(REG_T4_SOUTH_B1_fifo_value_O[0])
	);
	SliceWrapper_32_22_23 REG_T4_SOUTH_B1_end_value(
		.I(config_reg_1_O),
		.O(REG_T4_SOUTH_B1_end_value_O)
	);
	SliceWrapper_32_23_24 REG_T4_SOUTH_B1_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T4_SOUTH_B1_fifo_value_O)
	);
	SliceWrapper_32_24_25 REG_T4_SOUTH_B1_start_value(
		.I(config_reg_1_O),
		.O(REG_T4_SOUTH_B1_start_value_O)
	);
	SplitFifo_1 REG_T4_WEST_B1$SplitFifo_1_inst0(
		.data_in(MUX_SB_T4_WEST_SB_OUT_B1_O),
		.rst(reset),
		.start_fifo(REG_T4_WEST_B1_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T4_WEST_B1$SplitFifo_1_inst0_ready0),
		.data_out(REG_T4_WEST_B1$SplitFifo_1_inst0_data_out),
		.clk_en(and1_inst19_out[0]),
		.end_fifo(REG_T4_WEST_B1_end_value_O[0]),
		.valid0(MUX_SB_T4_WEST_SB_OUT_B1_valid_out),
		.valid1(REG_T4_WEST_B1$SplitFifo_1_inst0_valid1),
		.ready1(RMUX_T4_WEST_B1_ready_out),
		.fifo_en(REG_T4_WEST_B1_fifo_value_O[0])
	);
	SliceWrapper_32_25_26 REG_T4_WEST_B1_end_value(
		.I(config_reg_1_O),
		.O(REG_T4_WEST_B1_end_value_O)
	);
	SliceWrapper_32_26_27 REG_T4_WEST_B1_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T4_WEST_B1_fifo_value_O)
	);
	SliceWrapper_32_27_28 REG_T4_WEST_B1_start_value(
		.I(config_reg_1_O),
		.O(REG_T4_WEST_B1_start_value_O)
	);
	wire [1:0] RMUX_T0_EAST_B1_I;
	assign RMUX_T0_EAST_B1_I[1+:1] = REG_T0_EAST_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T0_EAST_B1_I[0+:1] = MUX_SB_T0_EAST_SB_OUT_B1_O;
	wire [1:0] RMUX_T0_EAST_B1_valid_in;
	assign RMUX_T0_EAST_B1_valid_in = {REG_T0_EAST_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T0_EAST_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T0_EAST_B1(
		.I(RMUX_T0_EAST_B1_I),
		.O(RMUX_T0_EAST_B1_O),
		.ready_in(SB_T0_EAST_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T0_EAST_B1_ready_out),
		.valid_in(RMUX_T0_EAST_B1_valid_in),
		.valid_out(RMUX_T0_EAST_B1_valid_out),
		.S(RMUX_T0_EAST_B1_sel_value_O),
		.out_sel(RMUX_T0_EAST_B1_out_sel)
	);
	SliceWrapper_32_28_29 RMUX_T0_EAST_B1_sel_value(
		.I(config_reg_1_O),
		.O(RMUX_T0_EAST_B1_sel_value_O)
	);
	wire [1:0] RMUX_T0_NORTH_B1_I;
	assign RMUX_T0_NORTH_B1_I[1+:1] = REG_T0_NORTH_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T0_NORTH_B1_I[0+:1] = MUX_SB_T0_NORTH_SB_OUT_B1_O;
	wire [1:0] RMUX_T0_NORTH_B1_valid_in;
	assign RMUX_T0_NORTH_B1_valid_in = {REG_T0_NORTH_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T0_NORTH_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T0_NORTH_B1(
		.I(RMUX_T0_NORTH_B1_I),
		.O(RMUX_T0_NORTH_B1_O),
		.ready_in(SB_T0_NORTH_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T0_NORTH_B1_ready_out),
		.valid_in(RMUX_T0_NORTH_B1_valid_in),
		.valid_out(RMUX_T0_NORTH_B1_valid_out),
		.S(RMUX_T0_NORTH_B1_sel_value_O),
		.out_sel(RMUX_T0_NORTH_B1_out_sel)
	);
	SliceWrapper_32_29_30 RMUX_T0_NORTH_B1_sel_value(
		.I(config_reg_1_O),
		.O(RMUX_T0_NORTH_B1_sel_value_O)
	);
	wire [1:0] RMUX_T0_SOUTH_B1_I;
	assign RMUX_T0_SOUTH_B1_I[1+:1] = REG_T0_SOUTH_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T0_SOUTH_B1_I[0+:1] = MUX_SB_T0_SOUTH_SB_OUT_B1_O;
	wire [1:0] RMUX_T0_SOUTH_B1_valid_in;
	assign RMUX_T0_SOUTH_B1_valid_in = {REG_T0_SOUTH_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T0_SOUTH_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T0_SOUTH_B1(
		.I(RMUX_T0_SOUTH_B1_I),
		.O(RMUX_T0_SOUTH_B1_O),
		.ready_in(SB_T0_SOUTH_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T0_SOUTH_B1_ready_out),
		.valid_in(RMUX_T0_SOUTH_B1_valid_in),
		.valid_out(RMUX_T0_SOUTH_B1_valid_out),
		.S(RMUX_T0_SOUTH_B1_sel_value_O),
		.out_sel(RMUX_T0_SOUTH_B1_out_sel)
	);
	SliceWrapper_32_30_31 RMUX_T0_SOUTH_B1_sel_value(
		.I(config_reg_1_O),
		.O(RMUX_T0_SOUTH_B1_sel_value_O)
	);
	wire [1:0] RMUX_T0_WEST_B1_I;
	assign RMUX_T0_WEST_B1_I[1+:1] = REG_T0_WEST_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T0_WEST_B1_I[0+:1] = MUX_SB_T0_WEST_SB_OUT_B1_O;
	wire [1:0] RMUX_T0_WEST_B1_valid_in;
	assign RMUX_T0_WEST_B1_valid_in = {REG_T0_WEST_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T0_WEST_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T0_WEST_B1(
		.I(RMUX_T0_WEST_B1_I),
		.O(RMUX_T0_WEST_B1_O),
		.ready_in(SB_T0_WEST_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T0_WEST_B1_ready_out),
		.valid_in(RMUX_T0_WEST_B1_valid_in),
		.valid_out(RMUX_T0_WEST_B1_valid_out),
		.S(RMUX_T0_WEST_B1_sel_value_O),
		.out_sel(RMUX_T0_WEST_B1_out_sel)
	);
	SliceWrapper_32_31_32 RMUX_T0_WEST_B1_sel_value(
		.I(config_reg_1_O),
		.O(RMUX_T0_WEST_B1_sel_value_O)
	);
	wire [1:0] RMUX_T1_EAST_B1_I;
	assign RMUX_T1_EAST_B1_I[1+:1] = REG_T1_EAST_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T1_EAST_B1_I[0+:1] = MUX_SB_T1_EAST_SB_OUT_B1_O;
	wire [1:0] RMUX_T1_EAST_B1_valid_in;
	assign RMUX_T1_EAST_B1_valid_in = {REG_T1_EAST_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T1_EAST_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T1_EAST_B1(
		.I(RMUX_T1_EAST_B1_I),
		.O(RMUX_T1_EAST_B1_O),
		.ready_in(SB_T1_EAST_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T1_EAST_B1_ready_out),
		.valid_in(RMUX_T1_EAST_B1_valid_in),
		.valid_out(RMUX_T1_EAST_B1_valid_out),
		.S(RMUX_T1_EAST_B1_sel_value_O),
		.out_sel(RMUX_T1_EAST_B1_out_sel)
	);
	SliceWrapper_32_0_1 RMUX_T1_EAST_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T1_EAST_B1_sel_value_O)
	);
	wire [1:0] RMUX_T1_NORTH_B1_I;
	assign RMUX_T1_NORTH_B1_I[1+:1] = REG_T1_NORTH_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T1_NORTH_B1_I[0+:1] = MUX_SB_T1_NORTH_SB_OUT_B1_O;
	wire [1:0] RMUX_T1_NORTH_B1_valid_in;
	assign RMUX_T1_NORTH_B1_valid_in = {REG_T1_NORTH_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T1_NORTH_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T1_NORTH_B1(
		.I(RMUX_T1_NORTH_B1_I),
		.O(RMUX_T1_NORTH_B1_O),
		.ready_in(SB_T1_NORTH_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T1_NORTH_B1_ready_out),
		.valid_in(RMUX_T1_NORTH_B1_valid_in),
		.valid_out(RMUX_T1_NORTH_B1_valid_out),
		.S(RMUX_T1_NORTH_B1_sel_value_O),
		.out_sel(RMUX_T1_NORTH_B1_out_sel)
	);
	SliceWrapper_32_1_2 RMUX_T1_NORTH_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T1_NORTH_B1_sel_value_O)
	);
	wire [1:0] RMUX_T1_SOUTH_B1_I;
	assign RMUX_T1_SOUTH_B1_I[1+:1] = REG_T1_SOUTH_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T1_SOUTH_B1_I[0+:1] = MUX_SB_T1_SOUTH_SB_OUT_B1_O;
	wire [1:0] RMUX_T1_SOUTH_B1_valid_in;
	assign RMUX_T1_SOUTH_B1_valid_in = {REG_T1_SOUTH_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T1_SOUTH_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T1_SOUTH_B1(
		.I(RMUX_T1_SOUTH_B1_I),
		.O(RMUX_T1_SOUTH_B1_O),
		.ready_in(SB_T1_SOUTH_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T1_SOUTH_B1_ready_out),
		.valid_in(RMUX_T1_SOUTH_B1_valid_in),
		.valid_out(RMUX_T1_SOUTH_B1_valid_out),
		.S(RMUX_T1_SOUTH_B1_sel_value_O),
		.out_sel(RMUX_T1_SOUTH_B1_out_sel)
	);
	SliceWrapper_32_2_3 RMUX_T1_SOUTH_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T1_SOUTH_B1_sel_value_O)
	);
	wire [1:0] RMUX_T1_WEST_B1_I;
	assign RMUX_T1_WEST_B1_I[1+:1] = REG_T1_WEST_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T1_WEST_B1_I[0+:1] = MUX_SB_T1_WEST_SB_OUT_B1_O;
	wire [1:0] RMUX_T1_WEST_B1_valid_in;
	assign RMUX_T1_WEST_B1_valid_in = {REG_T1_WEST_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T1_WEST_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T1_WEST_B1(
		.I(RMUX_T1_WEST_B1_I),
		.O(RMUX_T1_WEST_B1_O),
		.ready_in(SB_T1_WEST_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T1_WEST_B1_ready_out),
		.valid_in(RMUX_T1_WEST_B1_valid_in),
		.valid_out(RMUX_T1_WEST_B1_valid_out),
		.S(RMUX_T1_WEST_B1_sel_value_O),
		.out_sel(RMUX_T1_WEST_B1_out_sel)
	);
	SliceWrapper_32_3_4 RMUX_T1_WEST_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T1_WEST_B1_sel_value_O)
	);
	wire [1:0] RMUX_T2_EAST_B1_I;
	assign RMUX_T2_EAST_B1_I[1+:1] = REG_T2_EAST_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T2_EAST_B1_I[0+:1] = MUX_SB_T2_EAST_SB_OUT_B1_O;
	wire [1:0] RMUX_T2_EAST_B1_valid_in;
	assign RMUX_T2_EAST_B1_valid_in = {REG_T2_EAST_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T2_EAST_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T2_EAST_B1(
		.I(RMUX_T2_EAST_B1_I),
		.O(RMUX_T2_EAST_B1_O),
		.ready_in(SB_T2_EAST_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T2_EAST_B1_ready_out),
		.valid_in(RMUX_T2_EAST_B1_valid_in),
		.valid_out(RMUX_T2_EAST_B1_valid_out),
		.S(RMUX_T2_EAST_B1_sel_value_O),
		.out_sel(RMUX_T2_EAST_B1_out_sel)
	);
	SliceWrapper_32_4_5 RMUX_T2_EAST_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T2_EAST_B1_sel_value_O)
	);
	wire [1:0] RMUX_T2_NORTH_B1_I;
	assign RMUX_T2_NORTH_B1_I[1+:1] = REG_T2_NORTH_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T2_NORTH_B1_I[0+:1] = MUX_SB_T2_NORTH_SB_OUT_B1_O;
	wire [1:0] RMUX_T2_NORTH_B1_valid_in;
	assign RMUX_T2_NORTH_B1_valid_in = {REG_T2_NORTH_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T2_NORTH_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T2_NORTH_B1(
		.I(RMUX_T2_NORTH_B1_I),
		.O(RMUX_T2_NORTH_B1_O),
		.ready_in(SB_T2_NORTH_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T2_NORTH_B1_ready_out),
		.valid_in(RMUX_T2_NORTH_B1_valid_in),
		.valid_out(RMUX_T2_NORTH_B1_valid_out),
		.S(RMUX_T2_NORTH_B1_sel_value_O),
		.out_sel(RMUX_T2_NORTH_B1_out_sel)
	);
	SliceWrapper_32_5_6 RMUX_T2_NORTH_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T2_NORTH_B1_sel_value_O)
	);
	wire [1:0] RMUX_T2_SOUTH_B1_I;
	assign RMUX_T2_SOUTH_B1_I[1+:1] = REG_T2_SOUTH_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T2_SOUTH_B1_I[0+:1] = MUX_SB_T2_SOUTH_SB_OUT_B1_O;
	wire [1:0] RMUX_T2_SOUTH_B1_valid_in;
	assign RMUX_T2_SOUTH_B1_valid_in = {REG_T2_SOUTH_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T2_SOUTH_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T2_SOUTH_B1(
		.I(RMUX_T2_SOUTH_B1_I),
		.O(RMUX_T2_SOUTH_B1_O),
		.ready_in(SB_T2_SOUTH_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T2_SOUTH_B1_ready_out),
		.valid_in(RMUX_T2_SOUTH_B1_valid_in),
		.valid_out(RMUX_T2_SOUTH_B1_valid_out),
		.S(RMUX_T2_SOUTH_B1_sel_value_O),
		.out_sel(RMUX_T2_SOUTH_B1_out_sel)
	);
	SliceWrapper_32_6_7 RMUX_T2_SOUTH_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T2_SOUTH_B1_sel_value_O)
	);
	wire [1:0] RMUX_T2_WEST_B1_I;
	assign RMUX_T2_WEST_B1_I[1+:1] = REG_T2_WEST_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T2_WEST_B1_I[0+:1] = MUX_SB_T2_WEST_SB_OUT_B1_O;
	wire [1:0] RMUX_T2_WEST_B1_valid_in;
	assign RMUX_T2_WEST_B1_valid_in = {REG_T2_WEST_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T2_WEST_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T2_WEST_B1(
		.I(RMUX_T2_WEST_B1_I),
		.O(RMUX_T2_WEST_B1_O),
		.ready_in(SB_T2_WEST_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T2_WEST_B1_ready_out),
		.valid_in(RMUX_T2_WEST_B1_valid_in),
		.valid_out(RMUX_T2_WEST_B1_valid_out),
		.S(RMUX_T2_WEST_B1_sel_value_O),
		.out_sel(RMUX_T2_WEST_B1_out_sel)
	);
	SliceWrapper_32_7_8 RMUX_T2_WEST_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T2_WEST_B1_sel_value_O)
	);
	wire [1:0] RMUX_T3_EAST_B1_I;
	assign RMUX_T3_EAST_B1_I[1+:1] = REG_T3_EAST_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T3_EAST_B1_I[0+:1] = MUX_SB_T3_EAST_SB_OUT_B1_O;
	wire [1:0] RMUX_T3_EAST_B1_valid_in;
	assign RMUX_T3_EAST_B1_valid_in = {REG_T3_EAST_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T3_EAST_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T3_EAST_B1(
		.I(RMUX_T3_EAST_B1_I),
		.O(RMUX_T3_EAST_B1_O),
		.ready_in(SB_T3_EAST_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T3_EAST_B1_ready_out),
		.valid_in(RMUX_T3_EAST_B1_valid_in),
		.valid_out(RMUX_T3_EAST_B1_valid_out),
		.S(RMUX_T3_EAST_B1_sel_value_O),
		.out_sel(RMUX_T3_EAST_B1_out_sel)
	);
	SliceWrapper_32_8_9 RMUX_T3_EAST_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T3_EAST_B1_sel_value_O)
	);
	wire [1:0] RMUX_T3_NORTH_B1_I;
	assign RMUX_T3_NORTH_B1_I[1+:1] = REG_T3_NORTH_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T3_NORTH_B1_I[0+:1] = MUX_SB_T3_NORTH_SB_OUT_B1_O;
	wire [1:0] RMUX_T3_NORTH_B1_valid_in;
	assign RMUX_T3_NORTH_B1_valid_in = {REG_T3_NORTH_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T3_NORTH_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T3_NORTH_B1(
		.I(RMUX_T3_NORTH_B1_I),
		.O(RMUX_T3_NORTH_B1_O),
		.ready_in(SB_T3_NORTH_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T3_NORTH_B1_ready_out),
		.valid_in(RMUX_T3_NORTH_B1_valid_in),
		.valid_out(RMUX_T3_NORTH_B1_valid_out),
		.S(RMUX_T3_NORTH_B1_sel_value_O),
		.out_sel(RMUX_T3_NORTH_B1_out_sel)
	);
	SliceWrapper_32_9_10 RMUX_T3_NORTH_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T3_NORTH_B1_sel_value_O)
	);
	wire [1:0] RMUX_T3_SOUTH_B1_I;
	assign RMUX_T3_SOUTH_B1_I[1+:1] = REG_T3_SOUTH_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T3_SOUTH_B1_I[0+:1] = MUX_SB_T3_SOUTH_SB_OUT_B1_O;
	wire [1:0] RMUX_T3_SOUTH_B1_valid_in;
	assign RMUX_T3_SOUTH_B1_valid_in = {REG_T3_SOUTH_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T3_SOUTH_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T3_SOUTH_B1(
		.I(RMUX_T3_SOUTH_B1_I),
		.O(RMUX_T3_SOUTH_B1_O),
		.ready_in(SB_T3_SOUTH_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T3_SOUTH_B1_ready_out),
		.valid_in(RMUX_T3_SOUTH_B1_valid_in),
		.valid_out(RMUX_T3_SOUTH_B1_valid_out),
		.S(RMUX_T3_SOUTH_B1_sel_value_O),
		.out_sel(RMUX_T3_SOUTH_B1_out_sel)
	);
	SliceWrapper_32_10_11 RMUX_T3_SOUTH_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T3_SOUTH_B1_sel_value_O)
	);
	wire [1:0] RMUX_T3_WEST_B1_I;
	assign RMUX_T3_WEST_B1_I[1+:1] = REG_T3_WEST_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T3_WEST_B1_I[0+:1] = MUX_SB_T3_WEST_SB_OUT_B1_O;
	wire [1:0] RMUX_T3_WEST_B1_valid_in;
	assign RMUX_T3_WEST_B1_valid_in = {REG_T3_WEST_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T3_WEST_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T3_WEST_B1(
		.I(RMUX_T3_WEST_B1_I),
		.O(RMUX_T3_WEST_B1_O),
		.ready_in(SB_T3_WEST_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T3_WEST_B1_ready_out),
		.valid_in(RMUX_T3_WEST_B1_valid_in),
		.valid_out(RMUX_T3_WEST_B1_valid_out),
		.S(RMUX_T3_WEST_B1_sel_value_O),
		.out_sel(RMUX_T3_WEST_B1_out_sel)
	);
	SliceWrapper_32_11_12 RMUX_T3_WEST_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T3_WEST_B1_sel_value_O)
	);
	wire [1:0] RMUX_T4_EAST_B1_I;
	assign RMUX_T4_EAST_B1_I[1+:1] = REG_T4_EAST_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T4_EAST_B1_I[0+:1] = MUX_SB_T4_EAST_SB_OUT_B1_O;
	wire [1:0] RMUX_T4_EAST_B1_valid_in;
	assign RMUX_T4_EAST_B1_valid_in = {REG_T4_EAST_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T4_EAST_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T4_EAST_B1(
		.I(RMUX_T4_EAST_B1_I),
		.O(RMUX_T4_EAST_B1_O),
		.ready_in(SB_T4_EAST_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T4_EAST_B1_ready_out),
		.valid_in(RMUX_T4_EAST_B1_valid_in),
		.valid_out(RMUX_T4_EAST_B1_valid_out),
		.S(RMUX_T4_EAST_B1_sel_value_O),
		.out_sel(RMUX_T4_EAST_B1_out_sel)
	);
	SliceWrapper_32_12_13 RMUX_T4_EAST_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T4_EAST_B1_sel_value_O)
	);
	wire [1:0] RMUX_T4_NORTH_B1_I;
	assign RMUX_T4_NORTH_B1_I[1+:1] = REG_T4_NORTH_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T4_NORTH_B1_I[0+:1] = MUX_SB_T4_NORTH_SB_OUT_B1_O;
	wire [1:0] RMUX_T4_NORTH_B1_valid_in;
	assign RMUX_T4_NORTH_B1_valid_in = {REG_T4_NORTH_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T4_NORTH_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T4_NORTH_B1(
		.I(RMUX_T4_NORTH_B1_I),
		.O(RMUX_T4_NORTH_B1_O),
		.ready_in(SB_T4_NORTH_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T4_NORTH_B1_ready_out),
		.valid_in(RMUX_T4_NORTH_B1_valid_in),
		.valid_out(RMUX_T4_NORTH_B1_valid_out),
		.S(RMUX_T4_NORTH_B1_sel_value_O),
		.out_sel(RMUX_T4_NORTH_B1_out_sel)
	);
	SliceWrapper_32_13_14 RMUX_T4_NORTH_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T4_NORTH_B1_sel_value_O)
	);
	wire [1:0] RMUX_T4_SOUTH_B1_I;
	assign RMUX_T4_SOUTH_B1_I[1+:1] = REG_T4_SOUTH_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T4_SOUTH_B1_I[0+:1] = MUX_SB_T4_SOUTH_SB_OUT_B1_O;
	wire [1:0] RMUX_T4_SOUTH_B1_valid_in;
	assign RMUX_T4_SOUTH_B1_valid_in = {REG_T4_SOUTH_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T4_SOUTH_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T4_SOUTH_B1(
		.I(RMUX_T4_SOUTH_B1_I),
		.O(RMUX_T4_SOUTH_B1_O),
		.ready_in(SB_T4_SOUTH_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T4_SOUTH_B1_ready_out),
		.valid_in(RMUX_T4_SOUTH_B1_valid_in),
		.valid_out(RMUX_T4_SOUTH_B1_valid_out),
		.S(RMUX_T4_SOUTH_B1_sel_value_O),
		.out_sel(RMUX_T4_SOUTH_B1_out_sel)
	);
	SliceWrapper_32_14_15 RMUX_T4_SOUTH_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T4_SOUTH_B1_sel_value_O)
	);
	wire [1:0] RMUX_T4_WEST_B1_I;
	assign RMUX_T4_WEST_B1_I[1+:1] = REG_T4_WEST_B1$SplitFifo_1_inst0_data_out;
	assign RMUX_T4_WEST_B1_I[0+:1] = MUX_SB_T4_WEST_SB_OUT_B1_O;
	wire [1:0] RMUX_T4_WEST_B1_valid_in;
	assign RMUX_T4_WEST_B1_valid_in = {REG_T4_WEST_B1$SplitFifo_1_inst0_valid1[0], MUX_SB_T4_WEST_SB_OUT_B1_valid_out};
	mux_aoi_ready_valid_2_1 RMUX_T4_WEST_B1(
		.I(RMUX_T4_WEST_B1_I),
		.O(RMUX_T4_WEST_B1_O),
		.ready_in(SB_T4_WEST_SB_OUT_B1_ready_in),
		.ready_out(RMUX_T4_WEST_B1_ready_out),
		.valid_in(RMUX_T4_WEST_B1_valid_in),
		.valid_out(RMUX_T4_WEST_B1_valid_out),
		.S(RMUX_T4_WEST_B1_sel_value_O),
		.out_sel(RMUX_T4_WEST_B1_out_sel)
	);
	SliceWrapper_32_15_16 RMUX_T4_WEST_B1_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T4_WEST_B1_sel_value_O)
	);
	SliceWrapper_32_16_17 SB_T0_EAST_SB_IN_B1_enable_value(
		.I(config_reg_2_O),
		.O(SB_T0_EAST_SB_IN_B1_enable_value_O)
	);
	FanoutHash_4678C6877F96240E SB_T0_EAST_SB_IN_B1_fan_in(
		.E3(MEM_input_width_1_num_0_enable),
		.I5(const_0_1_out),
		.E0(SB_T0_WEST_SB_OUT_B1_enable_value_O),
		.S5(const_0_32_out),
		.S3(MEM_input_width_1_num_0_out_sel),
		.S4(MEM_input_width_1_num_1_out_sel),
		.I3(MEM_input_width_1_num_0_ready),
		.I4(MEM_input_width_1_num_1_ready),
		.S1(MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T0_WEST_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T4_NORTH_SB_OUT_B1_out_sel),
		.E2(SB_T4_NORTH_SB_OUT_B1_enable_value_O),
		.E5(const_0_1_out),
		.E4(MEM_input_width_1_num_1_enable),
		.I2(MUX_SB_T4_NORTH_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out),
		.O(SB_T0_EAST_SB_IN_B1_fan_in_O),
		.E1(SB_T3_SOUTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T0_WEST_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T0_EAST_SB_OUT_B1_FANOUT_I;
	assign SB_T0_EAST_SB_OUT_B1_FANOUT_I = {REG_T0_EAST_B1$SplitFifo_1_inst0_ready0[0], RMUX_T0_EAST_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T0_EAST_SB_OUT_B1_FANOUT(
		.O(SB_T0_EAST_SB_OUT_B1_FANOUT_O),
		.I(SB_T0_EAST_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T0_EAST_B1_out_sel)
	);
	SliceWrapper_32_17_18 SB_T0_EAST_SB_OUT_B1_enable_value(
		.I(config_reg_2_O),
		.O(SB_T0_EAST_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_32_18_21 SB_T0_EAST_SB_OUT_B1_sel_value(
		.I(config_reg_2_O),
		.O(SB_T0_EAST_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_32_21_22 SB_T0_NORTH_SB_IN_B1_enable_value(
		.I(config_reg_2_O),
		.O(SB_T0_NORTH_SB_IN_B1_enable_value_O)
	);
	FanoutHash_F95D10B01D02012 SB_T0_NORTH_SB_IN_B1_fan_in(
		.E3(MEM_input_width_1_num_0_enable),
		.I5(const_0_1_out),
		.E0(SB_T0_WEST_SB_OUT_B1_enable_value_O),
		.S5(const_0_32_out),
		.S3(MEM_input_width_1_num_0_out_sel),
		.S4(MEM_input_width_1_num_1_out_sel),
		.I3(MEM_input_width_1_num_0_ready),
		.I4(MEM_input_width_1_num_1_ready),
		.S1(MUX_SB_T1_EAST_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T0_WEST_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel),
		.E2(SB_T0_SOUTH_SB_OUT_B1_enable_value_O),
		.E5(const_0_1_out),
		.E4(MEM_input_width_1_num_1_enable),
		.I2(MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T1_EAST_SB_OUT_B1_ready_out),
		.O(SB_T0_NORTH_SB_IN_B1_fan_in_O),
		.E1(SB_T1_EAST_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T0_WEST_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T0_NORTH_SB_OUT_B1_FANOUT_I;
	assign SB_T0_NORTH_SB_OUT_B1_FANOUT_I = {REG_T0_NORTH_B1$SplitFifo_1_inst0_ready0[0], RMUX_T0_NORTH_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T0_NORTH_SB_OUT_B1_FANOUT(
		.O(SB_T0_NORTH_SB_OUT_B1_FANOUT_O),
		.I(SB_T0_NORTH_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T0_NORTH_B1_out_sel)
	);
	SliceWrapper_32_22_23 SB_T0_NORTH_SB_OUT_B1_enable_value(
		.I(config_reg_2_O),
		.O(SB_T0_NORTH_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_32_23_26 SB_T0_NORTH_SB_OUT_B1_sel_value(
		.I(config_reg_2_O),
		.O(SB_T0_NORTH_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_32_26_27 SB_T0_SOUTH_SB_IN_B1_enable_value(
		.I(config_reg_2_O),
		.O(SB_T0_SOUTH_SB_IN_B1_enable_value_O)
	);
	FanoutHash_99D793215CEDDD5 SB_T0_SOUTH_SB_IN_B1_fan_in(
		.E3(MEM_input_width_1_num_0_enable),
		.I5(const_0_1_out),
		.E0(SB_T3_EAST_SB_OUT_B1_enable_value_O),
		.S5(const_0_32_out),
		.S3(MEM_input_width_1_num_0_out_sel),
		.S4(MEM_input_width_1_num_1_out_sel),
		.I3(MEM_input_width_1_num_0_ready),
		.I4(MEM_input_width_1_num_1_ready),
		.S1(MUX_SB_T0_NORTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T3_EAST_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T1_WEST_SB_OUT_B1_out_sel),
		.E2(SB_T1_WEST_SB_OUT_B1_enable_value_O),
		.E5(const_0_1_out),
		.E4(MEM_input_width_1_num_1_enable),
		.I2(MUX_SB_T1_WEST_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T0_NORTH_SB_OUT_B1_ready_out),
		.O(SB_T0_SOUTH_SB_IN_B1_fan_in_O),
		.E1(SB_T0_NORTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T3_EAST_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T0_SOUTH_SB_OUT_B1_FANOUT_I;
	assign SB_T0_SOUTH_SB_OUT_B1_FANOUT_I = {REG_T0_SOUTH_B1$SplitFifo_1_inst0_ready0[0], RMUX_T0_SOUTH_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T0_SOUTH_SB_OUT_B1_FANOUT(
		.O(SB_T0_SOUTH_SB_OUT_B1_FANOUT_O),
		.I(SB_T0_SOUTH_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T0_SOUTH_B1_out_sel)
	);
	SliceWrapper_32_27_28 SB_T0_SOUTH_SB_OUT_B1_enable_value(
		.I(config_reg_2_O),
		.O(SB_T0_SOUTH_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_32_28_31 SB_T0_SOUTH_SB_OUT_B1_sel_value(
		.I(config_reg_2_O),
		.O(SB_T0_SOUTH_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_32_31_32 SB_T0_WEST_SB_IN_B1_enable_value(
		.I(config_reg_2_O),
		.O(SB_T0_WEST_SB_IN_B1_enable_value_O)
	);
	FanoutHash_3A0064632A577CF5 SB_T0_WEST_SB_IN_B1_fan_in(
		.E3(MEM_input_width_1_num_0_enable),
		.I5(const_0_1_out),
		.E0(SB_T0_NORTH_SB_OUT_B1_enable_value_O),
		.S5(const_0_32_out),
		.S3(MEM_input_width_1_num_0_out_sel),
		.S4(MEM_input_width_1_num_1_out_sel),
		.I3(MEM_input_width_1_num_0_ready),
		.I4(MEM_input_width_1_num_1_ready),
		.S1(MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T0_NORTH_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T0_EAST_SB_OUT_B1_out_sel),
		.E2(SB_T0_EAST_SB_OUT_B1_enable_value_O),
		.E5(const_0_1_out),
		.E4(MEM_input_width_1_num_1_enable),
		.I2(MUX_SB_T0_EAST_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out),
		.O(SB_T0_WEST_SB_IN_B1_fan_in_O),
		.E1(SB_T4_SOUTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T0_NORTH_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T0_WEST_SB_OUT_B1_FANOUT_I;
	assign SB_T0_WEST_SB_OUT_B1_FANOUT_I = {REG_T0_WEST_B1$SplitFifo_1_inst0_ready0[0], RMUX_T0_WEST_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T0_WEST_SB_OUT_B1_FANOUT(
		.O(SB_T0_WEST_SB_OUT_B1_FANOUT_O),
		.I(SB_T0_WEST_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T0_WEST_B1_out_sel)
	);
	SliceWrapper_31_0_1 SB_T0_WEST_SB_OUT_B1_enable_value(
		.I(config_reg_3_O),
		.O(SB_T0_WEST_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_31_1_4 SB_T0_WEST_SB_OUT_B1_sel_value(
		.I(config_reg_3_O),
		.O(SB_T0_WEST_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_31_4_5 SB_T1_EAST_SB_IN_B1_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_EAST_SB_IN_B1_enable_value_O)
	);
	FanoutHash_1130FCC7DFE98006 SB_T1_EAST_SB_IN_B1_fan_in(
		.E3(MEM_input_width_1_num_0_enable),
		.I5(const_0_1_out),
		.E0(SB_T0_NORTH_SB_OUT_B1_enable_value_O),
		.S5(const_0_32_out),
		.S3(MEM_input_width_1_num_0_out_sel),
		.S4(MEM_input_width_1_num_1_out_sel),
		.I3(MEM_input_width_1_num_0_ready),
		.I4(MEM_input_width_1_num_1_ready),
		.S1(MUX_SB_T1_WEST_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T0_NORTH_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel),
		.E2(SB_T2_SOUTH_SB_OUT_B1_enable_value_O),
		.E5(const_0_1_out),
		.E4(MEM_input_width_1_num_1_enable),
		.I2(MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T1_WEST_SB_OUT_B1_ready_out),
		.O(SB_T1_EAST_SB_IN_B1_fan_in_O),
		.E1(SB_T1_WEST_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T0_NORTH_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T1_EAST_SB_OUT_B1_FANOUT_I;
	assign SB_T1_EAST_SB_OUT_B1_FANOUT_I = {REG_T1_EAST_B1$SplitFifo_1_inst0_ready0[0], RMUX_T1_EAST_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T1_EAST_SB_OUT_B1_FANOUT(
		.O(SB_T1_EAST_SB_OUT_B1_FANOUT_O),
		.I(SB_T1_EAST_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T1_EAST_B1_out_sel)
	);
	SliceWrapper_31_5_6 SB_T1_EAST_SB_OUT_B1_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_EAST_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_31_6_9 SB_T1_EAST_SB_OUT_B1_sel_value(
		.I(config_reg_3_O),
		.O(SB_T1_EAST_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_31_9_10 SB_T1_NORTH_SB_IN_B1_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_NORTH_SB_IN_B1_enable_value_O)
	);
	FanoutHash_31555E0CDC460B97 SB_T1_NORTH_SB_IN_B1_fan_in(
		.E3(MEM_input_width_1_num_0_enable),
		.I5(const_0_1_out),
		.E0(SB_T2_EAST_SB_OUT_B1_enable_value_O),
		.S5(const_0_32_out),
		.S3(MEM_input_width_1_num_0_out_sel),
		.S4(MEM_input_width_1_num_1_out_sel),
		.I3(MEM_input_width_1_num_0_ready),
		.I4(MEM_input_width_1_num_1_ready),
		.S1(MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T2_EAST_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T4_WEST_SB_OUT_B1_out_sel),
		.E2(SB_T4_WEST_SB_OUT_B1_enable_value_O),
		.E5(const_0_1_out),
		.E4(MEM_input_width_1_num_1_enable),
		.I2(MUX_SB_T4_WEST_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out),
		.O(SB_T1_NORTH_SB_IN_B1_fan_in_O),
		.E1(SB_T1_SOUTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T2_EAST_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T1_NORTH_SB_OUT_B1_FANOUT_I;
	assign SB_T1_NORTH_SB_OUT_B1_FANOUT_I = {REG_T1_NORTH_B1$SplitFifo_1_inst0_ready0[0], RMUX_T1_NORTH_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T1_NORTH_SB_OUT_B1_FANOUT(
		.O(SB_T1_NORTH_SB_OUT_B1_FANOUT_O),
		.I(SB_T1_NORTH_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T1_NORTH_B1_out_sel)
	);
	SliceWrapper_31_10_11 SB_T1_NORTH_SB_OUT_B1_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_NORTH_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_31_11_14 SB_T1_NORTH_SB_OUT_B1_sel_value(
		.I(config_reg_3_O),
		.O(SB_T1_NORTH_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_31_14_15 SB_T1_SOUTH_SB_IN_B1_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_SOUTH_SB_IN_B1_enable_value_O)
	);
	FanoutHash_4FF010386DB0B737 SB_T1_SOUTH_SB_IN_B1_fan_in(
		.E3(MEM_input_width_1_num_0_enable),
		.I5(const_0_1_out),
		.E0(SB_T2_EAST_SB_OUT_B1_enable_value_O),
		.S5(const_0_32_out),
		.S3(MEM_input_width_1_num_0_out_sel),
		.S4(MEM_input_width_1_num_1_out_sel),
		.I3(MEM_input_width_1_num_0_ready),
		.I4(MEM_input_width_1_num_1_ready),
		.S1(MUX_SB_T1_NORTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T2_EAST_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T2_WEST_SB_OUT_B1_out_sel),
		.E2(SB_T2_WEST_SB_OUT_B1_enable_value_O),
		.E5(const_0_1_out),
		.E4(MEM_input_width_1_num_1_enable),
		.I2(MUX_SB_T2_WEST_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T1_NORTH_SB_OUT_B1_ready_out),
		.O(SB_T1_SOUTH_SB_IN_B1_fan_in_O),
		.E1(SB_T1_NORTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T2_EAST_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T1_SOUTH_SB_OUT_B1_FANOUT_I;
	assign SB_T1_SOUTH_SB_OUT_B1_FANOUT_I = {REG_T1_SOUTH_B1$SplitFifo_1_inst0_ready0[0], RMUX_T1_SOUTH_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T1_SOUTH_SB_OUT_B1_FANOUT(
		.O(SB_T1_SOUTH_SB_OUT_B1_FANOUT_O),
		.I(SB_T1_SOUTH_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T1_SOUTH_B1_out_sel)
	);
	SliceWrapper_31_15_16 SB_T1_SOUTH_SB_OUT_B1_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_SOUTH_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_31_16_19 SB_T1_SOUTH_SB_OUT_B1_sel_value(
		.I(config_reg_3_O),
		.O(SB_T1_SOUTH_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_31_19_20 SB_T1_WEST_SB_IN_B1_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_WEST_SB_IN_B1_enable_value_O)
	);
	FanoutHash_1A568579D8E9714B SB_T1_WEST_SB_IN_B1_fan_in(
		.E3(MEM_input_width_1_num_0_enable),
		.I5(const_0_1_out),
		.E0(SB_T4_NORTH_SB_OUT_B1_enable_value_O),
		.S5(const_0_32_out),
		.S3(MEM_input_width_1_num_0_out_sel),
		.S4(MEM_input_width_1_num_1_out_sel),
		.I3(MEM_input_width_1_num_0_ready),
		.I4(MEM_input_width_1_num_1_ready),
		.S1(MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T4_NORTH_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T1_EAST_SB_OUT_B1_out_sel),
		.E2(SB_T1_EAST_SB_OUT_B1_enable_value_O),
		.E5(const_0_1_out),
		.E4(MEM_input_width_1_num_1_enable),
		.I2(MUX_SB_T1_EAST_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out),
		.O(SB_T1_WEST_SB_IN_B1_fan_in_O),
		.E1(SB_T0_SOUTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T4_NORTH_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T1_WEST_SB_OUT_B1_FANOUT_I;
	assign SB_T1_WEST_SB_OUT_B1_FANOUT_I = {REG_T1_WEST_B1$SplitFifo_1_inst0_ready0[0], RMUX_T1_WEST_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T1_WEST_SB_OUT_B1_FANOUT(
		.O(SB_T1_WEST_SB_OUT_B1_FANOUT_O),
		.I(SB_T1_WEST_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T1_WEST_B1_out_sel)
	);
	SliceWrapper_31_20_21 SB_T1_WEST_SB_OUT_B1_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_WEST_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_31_21_24 SB_T1_WEST_SB_OUT_B1_sel_value(
		.I(config_reg_3_O),
		.O(SB_T1_WEST_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_31_24_25 SB_T2_EAST_SB_IN_B1_enable_value(
		.I(config_reg_3_O),
		.O(SB_T2_EAST_SB_IN_B1_enable_value_O)
	);
	FanoutHash_278348DB702230E6 SB_T2_EAST_SB_IN_B1_fan_in(
		.E3(MEM_input_width_1_num_0_enable),
		.I5(const_0_1_out),
		.E0(SB_T1_NORTH_SB_OUT_B1_enable_value_O),
		.S5(const_0_32_out),
		.S3(MEM_input_width_1_num_0_out_sel),
		.S4(MEM_input_width_1_num_1_out_sel),
		.I3(MEM_input_width_1_num_0_ready),
		.I4(MEM_input_width_1_num_1_ready),
		.S1(MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T1_NORTH_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T2_WEST_SB_OUT_B1_out_sel),
		.E2(SB_T2_WEST_SB_OUT_B1_enable_value_O),
		.E5(const_0_1_out),
		.E4(MEM_input_width_1_num_1_enable),
		.I2(MUX_SB_T2_WEST_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out),
		.O(SB_T2_EAST_SB_IN_B1_fan_in_O),
		.E1(SB_T1_SOUTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T1_NORTH_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T2_EAST_SB_OUT_B1_FANOUT_I;
	assign SB_T2_EAST_SB_OUT_B1_FANOUT_I = {REG_T2_EAST_B1$SplitFifo_1_inst0_ready0[0], RMUX_T2_EAST_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T2_EAST_SB_OUT_B1_FANOUT(
		.O(SB_T2_EAST_SB_OUT_B1_FANOUT_O),
		.I(SB_T2_EAST_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T2_EAST_B1_out_sel)
	);
	SliceWrapper_31_25_26 SB_T2_EAST_SB_OUT_B1_enable_value(
		.I(config_reg_3_O),
		.O(SB_T2_EAST_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_31_26_29 SB_T2_EAST_SB_OUT_B1_sel_value(
		.I(config_reg_3_O),
		.O(SB_T2_EAST_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_31_29_30 SB_T2_NORTH_SB_IN_B1_enable_value(
		.I(config_reg_3_O),
		.O(SB_T2_NORTH_SB_IN_B1_enable_value_O)
	);
	FanoutHash_6EB42FA08A9B7B5B SB_T2_NORTH_SB_IN_B1_fan_in(
		.E3(MEM_input_width_1_num_0_enable),
		.I5(const_0_1_out),
		.E0(SB_T3_EAST_SB_OUT_B1_enable_value_O),
		.S5(const_0_32_out),
		.S3(MEM_input_width_1_num_0_out_sel),
		.S4(MEM_input_width_1_num_1_out_sel),
		.I3(MEM_input_width_1_num_0_ready),
		.I4(MEM_input_width_1_num_1_ready),
		.S1(MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T3_EAST_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T3_WEST_SB_OUT_B1_out_sel),
		.E2(SB_T3_WEST_SB_OUT_B1_enable_value_O),
		.E5(const_0_1_out),
		.E4(MEM_input_width_1_num_1_enable),
		.I2(MUX_SB_T3_WEST_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out),
		.O(SB_T2_NORTH_SB_IN_B1_fan_in_O),
		.E1(SB_T2_SOUTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T3_EAST_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T2_NORTH_SB_OUT_B1_FANOUT_I;
	assign SB_T2_NORTH_SB_OUT_B1_FANOUT_I = {REG_T2_NORTH_B1$SplitFifo_1_inst0_ready0[0], RMUX_T2_NORTH_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T2_NORTH_SB_OUT_B1_FANOUT(
		.O(SB_T2_NORTH_SB_OUT_B1_FANOUT_O),
		.I(SB_T2_NORTH_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T2_NORTH_B1_out_sel)
	);
	SliceWrapper_31_30_31 SB_T2_NORTH_SB_OUT_B1_enable_value(
		.I(config_reg_3_O),
		.O(SB_T2_NORTH_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_30_0_3 SB_T2_NORTH_SB_OUT_B1_sel_value(
		.I(config_reg_4_O),
		.O(SB_T2_NORTH_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_30_3_4 SB_T2_SOUTH_SB_IN_B1_enable_value(
		.I(config_reg_4_O),
		.O(SB_T2_SOUTH_SB_IN_B1_enable_value_O)
	);
	FanoutHash_308BAC760F688049 SB_T2_SOUTH_SB_IN_B1_fan_in(
		.E3(MEM_input_width_1_num_0_enable),
		.I5(const_0_1_out),
		.E0(SB_T1_EAST_SB_OUT_B1_enable_value_O),
		.S5(const_0_32_out),
		.S3(MEM_input_width_1_num_0_out_sel),
		.S4(MEM_input_width_1_num_1_out_sel),
		.I3(MEM_input_width_1_num_0_ready),
		.I4(MEM_input_width_1_num_1_ready),
		.S1(MUX_SB_T2_NORTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T1_EAST_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T3_WEST_SB_OUT_B1_out_sel),
		.E2(SB_T3_WEST_SB_OUT_B1_enable_value_O),
		.E5(const_0_1_out),
		.E4(MEM_input_width_1_num_1_enable),
		.I2(MUX_SB_T3_WEST_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T2_NORTH_SB_OUT_B1_ready_out),
		.O(SB_T2_SOUTH_SB_IN_B1_fan_in_O),
		.E1(SB_T2_NORTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T1_EAST_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T2_SOUTH_SB_OUT_B1_FANOUT_I;
	assign SB_T2_SOUTH_SB_OUT_B1_FANOUT_I = {REG_T2_SOUTH_B1$SplitFifo_1_inst0_ready0[0], RMUX_T2_SOUTH_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T2_SOUTH_SB_OUT_B1_FANOUT(
		.O(SB_T2_SOUTH_SB_OUT_B1_FANOUT_O),
		.I(SB_T2_SOUTH_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T2_SOUTH_B1_out_sel)
	);
	SliceWrapper_30_4_5 SB_T2_SOUTH_SB_OUT_B1_enable_value(
		.I(config_reg_4_O),
		.O(SB_T2_SOUTH_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_30_5_8 SB_T2_SOUTH_SB_OUT_B1_sel_value(
		.I(config_reg_4_O),
		.O(SB_T2_SOUTH_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_30_8_9 SB_T2_WEST_SB_IN_B1_enable_value(
		.I(config_reg_4_O),
		.O(SB_T2_WEST_SB_IN_B1_enable_value_O)
	);
	FanoutHash_F8E7A0823DC8CDD SB_T2_WEST_SB_IN_B1_fan_in(
		.E3(MEM_input_width_1_num_0_enable),
		.I5(const_0_1_out),
		.E0(SB_T3_NORTH_SB_OUT_B1_enable_value_O),
		.S5(const_0_32_out),
		.S3(MEM_input_width_1_num_0_out_sel),
		.S4(MEM_input_width_1_num_1_out_sel),
		.I3(MEM_input_width_1_num_0_ready),
		.I4(MEM_input_width_1_num_1_ready),
		.S1(MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T3_NORTH_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T2_EAST_SB_OUT_B1_out_sel),
		.E2(SB_T2_EAST_SB_OUT_B1_enable_value_O),
		.E5(const_0_1_out),
		.E4(MEM_input_width_1_num_1_enable),
		.I2(MUX_SB_T2_EAST_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out),
		.O(SB_T2_WEST_SB_IN_B1_fan_in_O),
		.E1(SB_T1_SOUTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T3_NORTH_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T2_WEST_SB_OUT_B1_FANOUT_I;
	assign SB_T2_WEST_SB_OUT_B1_FANOUT_I = {REG_T2_WEST_B1$SplitFifo_1_inst0_ready0[0], RMUX_T2_WEST_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T2_WEST_SB_OUT_B1_FANOUT(
		.O(SB_T2_WEST_SB_OUT_B1_FANOUT_O),
		.I(SB_T2_WEST_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T2_WEST_B1_out_sel)
	);
	SliceWrapper_30_9_10 SB_T2_WEST_SB_OUT_B1_enable_value(
		.I(config_reg_4_O),
		.O(SB_T2_WEST_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_30_10_13 SB_T2_WEST_SB_OUT_B1_sel_value(
		.I(config_reg_4_O),
		.O(SB_T2_WEST_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_30_13_14 SB_T3_EAST_SB_IN_B1_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_EAST_SB_IN_B1_enable_value_O)
	);
	FanoutHash_D70CFBE8EA3CE7F SB_T3_EAST_SB_IN_B1_fan_in(
		.E3(MEM_input_width_1_num_0_enable),
		.I5(const_0_1_out),
		.E0(SB_T0_SOUTH_SB_OUT_B1_enable_value_O),
		.S5(const_0_32_out),
		.S3(MEM_input_width_1_num_0_out_sel),
		.S4(MEM_input_width_1_num_1_out_sel),
		.I3(MEM_input_width_1_num_0_ready),
		.I4(MEM_input_width_1_num_1_ready),
		.S1(MUX_SB_T2_NORTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T3_WEST_SB_OUT_B1_out_sel),
		.E2(SB_T3_WEST_SB_OUT_B1_enable_value_O),
		.E5(const_0_1_out),
		.E4(MEM_input_width_1_num_1_enable),
		.I2(MUX_SB_T3_WEST_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T2_NORTH_SB_OUT_B1_ready_out),
		.O(SB_T3_EAST_SB_IN_B1_fan_in_O),
		.E1(SB_T2_NORTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T3_EAST_SB_OUT_B1_FANOUT_I;
	assign SB_T3_EAST_SB_OUT_B1_FANOUT_I = {REG_T3_EAST_B1$SplitFifo_1_inst0_ready0[0], RMUX_T3_EAST_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T3_EAST_SB_OUT_B1_FANOUT(
		.O(SB_T3_EAST_SB_OUT_B1_FANOUT_O),
		.I(SB_T3_EAST_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T3_EAST_B1_out_sel)
	);
	SliceWrapper_30_14_15 SB_T3_EAST_SB_OUT_B1_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_EAST_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_30_15_18 SB_T3_EAST_SB_OUT_B1_sel_value(
		.I(config_reg_4_O),
		.O(SB_T3_EAST_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_30_18_19 SB_T3_NORTH_SB_IN_B1_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_NORTH_SB_IN_B1_enable_value_O)
	);
	FanoutHash_5DE101F5B6936D07 SB_T3_NORTH_SB_IN_B1_fan_in(
		.E3(MEM_input_width_1_num_0_enable),
		.I5(const_0_1_out),
		.E0(SB_T2_WEST_SB_OUT_B1_enable_value_O),
		.S5(const_0_32_out),
		.S3(MEM_input_width_1_num_0_out_sel),
		.S4(MEM_input_width_1_num_1_out_sel),
		.I3(MEM_input_width_1_num_0_ready),
		.I4(MEM_input_width_1_num_1_ready),
		.S1(MUX_SB_T4_EAST_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T2_WEST_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel),
		.E2(SB_T3_SOUTH_SB_OUT_B1_enable_value_O),
		.E5(const_0_1_out),
		.E4(MEM_input_width_1_num_1_enable),
		.I2(MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T4_EAST_SB_OUT_B1_ready_out),
		.O(SB_T3_NORTH_SB_IN_B1_fan_in_O),
		.E1(SB_T4_EAST_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T2_WEST_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T3_NORTH_SB_OUT_B1_FANOUT_I;
	assign SB_T3_NORTH_SB_OUT_B1_FANOUT_I = {REG_T3_NORTH_B1$SplitFifo_1_inst0_ready0[0], RMUX_T3_NORTH_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T3_NORTH_SB_OUT_B1_FANOUT(
		.O(SB_T3_NORTH_SB_OUT_B1_FANOUT_O),
		.I(SB_T3_NORTH_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T3_NORTH_B1_out_sel)
	);
	SliceWrapper_30_19_20 SB_T3_NORTH_SB_OUT_B1_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_NORTH_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_30_20_23 SB_T3_NORTH_SB_OUT_B1_sel_value(
		.I(config_reg_4_O),
		.O(SB_T3_NORTH_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_30_23_24 SB_T3_SOUTH_SB_IN_B1_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_SOUTH_SB_IN_B1_enable_value_O)
	);
	FanoutHash_13B77C2790BDE4E2 SB_T3_SOUTH_SB_IN_B1_fan_in(
		.E3(MEM_input_width_1_num_0_enable),
		.I5(const_0_1_out),
		.E0(SB_T0_EAST_SB_OUT_B1_enable_value_O),
		.S5(const_0_32_out),
		.S3(MEM_input_width_1_num_0_out_sel),
		.S4(MEM_input_width_1_num_1_out_sel),
		.I3(MEM_input_width_1_num_0_ready),
		.I4(MEM_input_width_1_num_1_ready),
		.S1(MUX_SB_T3_NORTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T0_EAST_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T4_WEST_SB_OUT_B1_out_sel),
		.E2(SB_T4_WEST_SB_OUT_B1_enable_value_O),
		.E5(const_0_1_out),
		.E4(MEM_input_width_1_num_1_enable),
		.I2(MUX_SB_T4_WEST_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T3_NORTH_SB_OUT_B1_ready_out),
		.O(SB_T3_SOUTH_SB_IN_B1_fan_in_O),
		.E1(SB_T3_NORTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T0_EAST_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T3_SOUTH_SB_OUT_B1_FANOUT_I;
	assign SB_T3_SOUTH_SB_OUT_B1_FANOUT_I = {REG_T3_SOUTH_B1$SplitFifo_1_inst0_ready0[0], RMUX_T3_SOUTH_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T3_SOUTH_SB_OUT_B1_FANOUT(
		.O(SB_T3_SOUTH_SB_OUT_B1_FANOUT_O),
		.I(SB_T3_SOUTH_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T3_SOUTH_B1_out_sel)
	);
	SliceWrapper_30_24_25 SB_T3_SOUTH_SB_OUT_B1_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_SOUTH_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_30_25_28 SB_T3_SOUTH_SB_OUT_B1_sel_value(
		.I(config_reg_4_O),
		.O(SB_T3_SOUTH_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_30_28_29 SB_T3_WEST_SB_IN_B1_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_WEST_SB_IN_B1_enable_value_O)
	);
	FanoutHash_7FDF2D3240D4A947 SB_T3_WEST_SB_IN_B1_fan_in(
		.E3(MEM_input_width_1_num_0_enable),
		.I5(const_0_1_out),
		.E0(SB_T2_NORTH_SB_OUT_B1_enable_value_O),
		.S5(const_0_32_out),
		.S3(MEM_input_width_1_num_0_out_sel),
		.S4(MEM_input_width_1_num_1_out_sel),
		.I3(MEM_input_width_1_num_0_ready),
		.I4(MEM_input_width_1_num_1_ready),
		.S1(MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T2_NORTH_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T3_EAST_SB_OUT_B1_out_sel),
		.E2(SB_T3_EAST_SB_OUT_B1_enable_value_O),
		.E5(const_0_1_out),
		.E4(MEM_input_width_1_num_1_enable),
		.I2(MUX_SB_T3_EAST_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out),
		.O(SB_T3_WEST_SB_IN_B1_fan_in_O),
		.E1(SB_T2_SOUTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T2_NORTH_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T3_WEST_SB_OUT_B1_FANOUT_I;
	assign SB_T3_WEST_SB_OUT_B1_FANOUT_I = {REG_T3_WEST_B1$SplitFifo_1_inst0_ready0[0], RMUX_T3_WEST_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T3_WEST_SB_OUT_B1_FANOUT(
		.O(SB_T3_WEST_SB_OUT_B1_FANOUT_O),
		.I(SB_T3_WEST_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T3_WEST_B1_out_sel)
	);
	SliceWrapper_30_29_30 SB_T3_WEST_SB_OUT_B1_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_WEST_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_23_0_3 SB_T3_WEST_SB_OUT_B1_sel_value(
		.I(config_reg_5_O),
		.O(SB_T3_WEST_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_23_3_4 SB_T4_EAST_SB_IN_B1_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_EAST_SB_IN_B1_enable_value_O)
	);
	FanoutHash_11B554A18790BBBC SB_T4_EAST_SB_IN_B1_fan_in(
		.E3(MEM_input_width_1_num_0_enable),
		.I5(const_0_1_out),
		.E0(SB_T3_NORTH_SB_OUT_B1_enable_value_O),
		.S5(const_0_32_out),
		.S3(MEM_input_width_1_num_0_out_sel),
		.S4(MEM_input_width_1_num_1_out_sel),
		.I3(MEM_input_width_1_num_0_ready),
		.I4(MEM_input_width_1_num_1_ready),
		.S1(MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T3_NORTH_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T4_WEST_SB_OUT_B1_out_sel),
		.E2(SB_T4_WEST_SB_OUT_B1_enable_value_O),
		.E5(const_0_1_out),
		.E4(MEM_input_width_1_num_1_enable),
		.I2(MUX_SB_T4_WEST_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out),
		.O(SB_T4_EAST_SB_IN_B1_fan_in_O),
		.E1(SB_T4_SOUTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T3_NORTH_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T4_EAST_SB_OUT_B1_FANOUT_I;
	assign SB_T4_EAST_SB_OUT_B1_FANOUT_I = {REG_T4_EAST_B1$SplitFifo_1_inst0_ready0[0], RMUX_T4_EAST_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T4_EAST_SB_OUT_B1_FANOUT(
		.O(SB_T4_EAST_SB_OUT_B1_FANOUT_O),
		.I(SB_T4_EAST_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T4_EAST_B1_out_sel)
	);
	SliceWrapper_23_4_5 SB_T4_EAST_SB_OUT_B1_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_EAST_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_23_5_8 SB_T4_EAST_SB_OUT_B1_sel_value(
		.I(config_reg_5_O),
		.O(SB_T4_EAST_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_23_8_9 SB_T4_NORTH_SB_IN_B1_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_NORTH_SB_IN_B1_enable_value_O)
	);
	FanoutHash_37B926A0CDF82FCC SB_T4_NORTH_SB_IN_B1_fan_in(
		.E3(MEM_input_width_1_num_0_enable),
		.I5(const_0_1_out),
		.E0(SB_T1_WEST_SB_OUT_B1_enable_value_O),
		.S5(const_0_32_out),
		.S3(MEM_input_width_1_num_0_out_sel),
		.S4(MEM_input_width_1_num_1_out_sel),
		.I3(MEM_input_width_1_num_0_ready),
		.I4(MEM_input_width_1_num_1_ready),
		.S1(MUX_SB_T0_EAST_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T1_WEST_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel),
		.E2(SB_T4_SOUTH_SB_OUT_B1_enable_value_O),
		.E5(const_0_1_out),
		.E4(MEM_input_width_1_num_1_enable),
		.I2(MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T0_EAST_SB_OUT_B1_ready_out),
		.O(SB_T4_NORTH_SB_IN_B1_fan_in_O),
		.E1(SB_T0_EAST_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T1_WEST_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T4_NORTH_SB_OUT_B1_FANOUT_I;
	assign SB_T4_NORTH_SB_OUT_B1_FANOUT_I = {REG_T4_NORTH_B1$SplitFifo_1_inst0_ready0[0], RMUX_T4_NORTH_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T4_NORTH_SB_OUT_B1_FANOUT(
		.O(SB_T4_NORTH_SB_OUT_B1_FANOUT_O),
		.I(SB_T4_NORTH_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T4_NORTH_B1_out_sel)
	);
	SliceWrapper_23_9_10 SB_T4_NORTH_SB_OUT_B1_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_NORTH_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_23_10_13 SB_T4_NORTH_SB_OUT_B1_sel_value(
		.I(config_reg_5_O),
		.O(SB_T4_NORTH_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_23_13_14 SB_T4_SOUTH_SB_IN_B1_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_SOUTH_SB_IN_B1_enable_value_O)
	);
	FanoutHash_1B10C32F008C11AC SB_T4_SOUTH_SB_IN_B1_fan_in(
		.E3(MEM_input_width_1_num_0_enable),
		.I5(const_0_1_out),
		.E0(SB_T0_WEST_SB_OUT_B1_enable_value_O),
		.S5(const_0_32_out),
		.S3(MEM_input_width_1_num_0_out_sel),
		.S4(MEM_input_width_1_num_1_out_sel),
		.I3(MEM_input_width_1_num_0_ready),
		.I4(MEM_input_width_1_num_1_ready),
		.S1(MUX_SB_T4_EAST_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T0_WEST_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T4_NORTH_SB_OUT_B1_out_sel),
		.E2(SB_T4_NORTH_SB_OUT_B1_enable_value_O),
		.E5(const_0_1_out),
		.E4(MEM_input_width_1_num_1_enable),
		.I2(MUX_SB_T4_NORTH_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T4_EAST_SB_OUT_B1_ready_out),
		.O(SB_T4_SOUTH_SB_IN_B1_fan_in_O),
		.E1(SB_T4_EAST_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T0_WEST_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T4_SOUTH_SB_OUT_B1_FANOUT_I;
	assign SB_T4_SOUTH_SB_OUT_B1_FANOUT_I = {REG_T4_SOUTH_B1$SplitFifo_1_inst0_ready0[0], RMUX_T4_SOUTH_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T4_SOUTH_SB_OUT_B1_FANOUT(
		.O(SB_T4_SOUTH_SB_OUT_B1_FANOUT_O),
		.I(SB_T4_SOUTH_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T4_SOUTH_B1_out_sel)
	);
	SliceWrapper_23_14_15 SB_T4_SOUTH_SB_OUT_B1_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_SOUTH_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_23_15_18 SB_T4_SOUTH_SB_OUT_B1_sel_value(
		.I(config_reg_5_O),
		.O(SB_T4_SOUTH_SB_OUT_B1_sel_value_O)
	);
	SliceWrapper_23_18_19 SB_T4_WEST_SB_IN_B1_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_WEST_SB_IN_B1_enable_value_O)
	);
	FanoutHash_660E59B0DDACF452 SB_T4_WEST_SB_IN_B1_fan_in(
		.E3(MEM_input_width_1_num_0_enable),
		.I5(const_0_1_out),
		.E0(SB_T1_NORTH_SB_OUT_B1_enable_value_O),
		.S5(const_0_32_out),
		.S3(MEM_input_width_1_num_0_out_sel),
		.S4(MEM_input_width_1_num_1_out_sel),
		.I3(MEM_input_width_1_num_0_ready),
		.I4(MEM_input_width_1_num_1_ready),
		.S1(MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel),
		.S0(MUX_SB_T1_NORTH_SB_OUT_B1_out_sel),
		.S2(MUX_SB_T4_EAST_SB_OUT_B1_out_sel),
		.E2(SB_T4_EAST_SB_OUT_B1_enable_value_O),
		.E5(const_0_1_out),
		.E4(MEM_input_width_1_num_1_enable),
		.I2(MUX_SB_T4_EAST_SB_OUT_B1_ready_out),
		.I1(MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out),
		.O(SB_T4_WEST_SB_IN_B1_fan_in_O),
		.E1(SB_T3_SOUTH_SB_OUT_B1_enable_value_O),
		.I0(MUX_SB_T1_NORTH_SB_OUT_B1_ready_out)
	);
	wire [1:0] SB_T4_WEST_SB_OUT_B1_FANOUT_I;
	assign SB_T4_WEST_SB_OUT_B1_FANOUT_I = {REG_T4_WEST_B1$SplitFifo_1_inst0_ready0[0], RMUX_T4_WEST_B1_ready_out};
	ExclusiveNodeFanout_H2 SB_T4_WEST_SB_OUT_B1_FANOUT(
		.O(SB_T4_WEST_SB_OUT_B1_FANOUT_O),
		.I(SB_T4_WEST_SB_OUT_B1_FANOUT_I),
		.S(RMUX_T4_WEST_B1_out_sel)
	);
	SliceWrapper_23_19_20 SB_T4_WEST_SB_OUT_B1_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_WEST_SB_OUT_B1_enable_value_O)
	);
	SliceWrapper_23_20_23 SB_T4_WEST_SB_OUT_B1_sel_value(
		.I(config_reg_5_O),
		.O(SB_T4_WEST_SB_OUT_B1_sel_value_O)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T0_EAST_SB_IN_B1(
		.I(SB_T0_EAST_SB_IN_B1),
		.O(WIRE_SB_T0_EAST_SB_IN_B1_O),
		.ready_in(SB_T0_EAST_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T0_EAST_SB_IN_B1_ready_out),
		.valid_in(SB_T0_EAST_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T0_EAST_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T0_NORTH_SB_IN_B1(
		.I(SB_T0_NORTH_SB_IN_B1),
		.O(WIRE_SB_T0_NORTH_SB_IN_B1_O),
		.ready_in(SB_T0_NORTH_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T0_NORTH_SB_IN_B1_ready_out),
		.valid_in(SB_T0_NORTH_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T0_NORTH_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T0_SOUTH_SB_IN_B1(
		.I(SB_T0_SOUTH_SB_IN_B1),
		.O(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
		.ready_in(SB_T0_SOUTH_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T0_SOUTH_SB_IN_B1_ready_out),
		.valid_in(SB_T0_SOUTH_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T0_SOUTH_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T0_WEST_SB_IN_B1(
		.I(SB_T0_WEST_SB_IN_B1),
		.O(WIRE_SB_T0_WEST_SB_IN_B1_O),
		.ready_in(SB_T0_WEST_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T0_WEST_SB_IN_B1_ready_out),
		.valid_in(SB_T0_WEST_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T0_WEST_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T1_EAST_SB_IN_B1(
		.I(SB_T1_EAST_SB_IN_B1),
		.O(WIRE_SB_T1_EAST_SB_IN_B1_O),
		.ready_in(SB_T1_EAST_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T1_EAST_SB_IN_B1_ready_out),
		.valid_in(SB_T1_EAST_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T1_EAST_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T1_NORTH_SB_IN_B1(
		.I(SB_T1_NORTH_SB_IN_B1),
		.O(WIRE_SB_T1_NORTH_SB_IN_B1_O),
		.ready_in(SB_T1_NORTH_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T1_NORTH_SB_IN_B1_ready_out),
		.valid_in(SB_T1_NORTH_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T1_NORTH_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T1_SOUTH_SB_IN_B1(
		.I(SB_T1_SOUTH_SB_IN_B1),
		.O(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
		.ready_in(SB_T1_SOUTH_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T1_SOUTH_SB_IN_B1_ready_out),
		.valid_in(SB_T1_SOUTH_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T1_SOUTH_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T1_WEST_SB_IN_B1(
		.I(SB_T1_WEST_SB_IN_B1),
		.O(WIRE_SB_T1_WEST_SB_IN_B1_O),
		.ready_in(SB_T1_WEST_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T1_WEST_SB_IN_B1_ready_out),
		.valid_in(SB_T1_WEST_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T1_WEST_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T2_EAST_SB_IN_B1(
		.I(SB_T2_EAST_SB_IN_B1),
		.O(WIRE_SB_T2_EAST_SB_IN_B1_O),
		.ready_in(SB_T2_EAST_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T2_EAST_SB_IN_B1_ready_out),
		.valid_in(SB_T2_EAST_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T2_EAST_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T2_NORTH_SB_IN_B1(
		.I(SB_T2_NORTH_SB_IN_B1),
		.O(WIRE_SB_T2_NORTH_SB_IN_B1_O),
		.ready_in(SB_T2_NORTH_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T2_NORTH_SB_IN_B1_ready_out),
		.valid_in(SB_T2_NORTH_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T2_NORTH_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T2_SOUTH_SB_IN_B1(
		.I(SB_T2_SOUTH_SB_IN_B1),
		.O(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
		.ready_in(SB_T2_SOUTH_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T2_SOUTH_SB_IN_B1_ready_out),
		.valid_in(SB_T2_SOUTH_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T2_SOUTH_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T2_WEST_SB_IN_B1(
		.I(SB_T2_WEST_SB_IN_B1),
		.O(WIRE_SB_T2_WEST_SB_IN_B1_O),
		.ready_in(SB_T2_WEST_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T2_WEST_SB_IN_B1_ready_out),
		.valid_in(SB_T2_WEST_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T2_WEST_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T3_EAST_SB_IN_B1(
		.I(SB_T3_EAST_SB_IN_B1),
		.O(WIRE_SB_T3_EAST_SB_IN_B1_O),
		.ready_in(SB_T3_EAST_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T3_EAST_SB_IN_B1_ready_out),
		.valid_in(SB_T3_EAST_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T3_EAST_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T3_NORTH_SB_IN_B1(
		.I(SB_T3_NORTH_SB_IN_B1),
		.O(WIRE_SB_T3_NORTH_SB_IN_B1_O),
		.ready_in(SB_T3_NORTH_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T3_NORTH_SB_IN_B1_ready_out),
		.valid_in(SB_T3_NORTH_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T3_NORTH_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T3_SOUTH_SB_IN_B1(
		.I(SB_T3_SOUTH_SB_IN_B1),
		.O(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
		.ready_in(SB_T3_SOUTH_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T3_SOUTH_SB_IN_B1_ready_out),
		.valid_in(SB_T3_SOUTH_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T3_SOUTH_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T3_WEST_SB_IN_B1(
		.I(SB_T3_WEST_SB_IN_B1),
		.O(WIRE_SB_T3_WEST_SB_IN_B1_O),
		.ready_in(SB_T3_WEST_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T3_WEST_SB_IN_B1_ready_out),
		.valid_in(SB_T3_WEST_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T3_WEST_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T4_EAST_SB_IN_B1(
		.I(SB_T4_EAST_SB_IN_B1),
		.O(WIRE_SB_T4_EAST_SB_IN_B1_O),
		.ready_in(SB_T4_EAST_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T4_EAST_SB_IN_B1_ready_out),
		.valid_in(SB_T4_EAST_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T4_EAST_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T4_NORTH_SB_IN_B1(
		.I(SB_T4_NORTH_SB_IN_B1),
		.O(WIRE_SB_T4_NORTH_SB_IN_B1_O),
		.ready_in(SB_T4_NORTH_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T4_NORTH_SB_IN_B1_ready_out),
		.valid_in(SB_T4_NORTH_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T4_NORTH_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T4_SOUTH_SB_IN_B1(
		.I(SB_T4_SOUTH_SB_IN_B1),
		.O(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
		.ready_in(SB_T4_SOUTH_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T4_SOUTH_SB_IN_B1_ready_out),
		.valid_in(SB_T4_SOUTH_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T4_SOUTH_SB_IN_B1_valid_out)
	);
	MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T4_WEST_SB_IN_B1(
		.I(SB_T4_WEST_SB_IN_B1),
		.O(WIRE_SB_T4_WEST_SB_IN_B1_O),
		.ready_in(SB_T4_WEST_SB_IN_B1_fan_in_O[0]),
		.ready_out(WIRE_SB_T4_WEST_SB_IN_B1_ready_out),
		.valid_in(SB_T4_WEST_SB_IN_B1_valid_in),
		.valid_out(WIRE_SB_T4_WEST_SB_IN_B1_valid_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_23_32_inst0$bit_const_0_None(.out(ZextWrapper_23_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_23_32_inst0$self_O_out;
	assign ZextWrapper_23_32_inst0$self_O_out = {ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, config_reg_5_O};
	mantle_wire__typeBitIn32 ZextWrapper_23_32_inst0$self_O(
		.in(ZextWrapper_23_32_inst0$self_O_in),
		.out(ZextWrapper_23_32_inst0$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_30_32_inst0$bit_const_0_None(.out(ZextWrapper_30_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_30_32_inst0$self_O_out;
	assign ZextWrapper_30_32_inst0$self_O_out = {ZextWrapper_30_32_inst0$bit_const_0_None_out, ZextWrapper_30_32_inst0$bit_const_0_None_out, config_reg_4_O};
	mantle_wire__typeBitIn32 ZextWrapper_30_32_inst0$self_O(
		.in(ZextWrapper_30_32_inst0$self_O_in),
		.out(ZextWrapper_30_32_inst0$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_31_32_inst0$bit_const_0_None(.out(ZextWrapper_31_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_31_32_inst0$self_O_out;
	assign ZextWrapper_31_32_inst0$self_O_out = {ZextWrapper_31_32_inst0$bit_const_0_None_out, config_reg_3_O};
	mantle_wire__typeBitIn32 ZextWrapper_31_32_inst0$self_O(
		.in(ZextWrapper_31_32_inst0$self_O_in),
		.out(ZextWrapper_31_32_inst0$self_O_out)
	);
	coreir_and #(.width(1)) and1_inst0(
		.in0(coreir_eq_1_inst0_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst0_out)
	);
	coreir_and #(.width(1)) and1_inst1(
		.in0(coreir_eq_1_inst1_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst1_out)
	);
	coreir_and #(.width(1)) and1_inst10(
		.in0(coreir_eq_1_inst10_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst10_out)
	);
	coreir_and #(.width(1)) and1_inst11(
		.in0(coreir_eq_1_inst11_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst11_out)
	);
	coreir_and #(.width(1)) and1_inst12(
		.in0(coreir_eq_1_inst12_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst12_out)
	);
	coreir_and #(.width(1)) and1_inst13(
		.in0(coreir_eq_1_inst13_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst13_out)
	);
	coreir_and #(.width(1)) and1_inst14(
		.in0(coreir_eq_1_inst14_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst14_out)
	);
	coreir_and #(.width(1)) and1_inst15(
		.in0(coreir_eq_1_inst15_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst15_out)
	);
	coreir_and #(.width(1)) and1_inst16(
		.in0(coreir_eq_1_inst16_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst16_out)
	);
	coreir_and #(.width(1)) and1_inst17(
		.in0(coreir_eq_1_inst17_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst17_out)
	);
	coreir_and #(.width(1)) and1_inst18(
		.in0(coreir_eq_1_inst18_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst18_out)
	);
	coreir_and #(.width(1)) and1_inst19(
		.in0(coreir_eq_1_inst19_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst19_out)
	);
	coreir_and #(.width(1)) and1_inst2(
		.in0(coreir_eq_1_inst2_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst2_out)
	);
	coreir_and #(.width(1)) and1_inst3(
		.in0(coreir_eq_1_inst3_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst3_out)
	);
	coreir_and #(.width(1)) and1_inst4(
		.in0(coreir_eq_1_inst4_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst4_out)
	);
	coreir_and #(.width(1)) and1_inst5(
		.in0(coreir_eq_1_inst5_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst5_out)
	);
	coreir_and #(.width(1)) and1_inst6(
		.in0(coreir_eq_1_inst6_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst6_out)
	);
	coreir_and #(.width(1)) and1_inst7(
		.in0(coreir_eq_1_inst7_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst7_out)
	);
	coreir_and #(.width(1)) and1_inst8(
		.in0(coreir_eq_1_inst8_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst8_out)
	);
	coreir_and #(.width(1)) and1_inst9(
		.in0(coreir_eq_1_inst9_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst9_out)
	);
	wire [7:0] config_reg_0_config_addr;
	assign config_reg_0_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4], self_config_config_addr_out[3], self_config_config_addr_out[2:0]};
	ConfigRegister_32_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_reg_0_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_1_config_addr;
	assign config_reg_1_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4], self_config_config_addr_out[3], self_config_config_addr_out[2:0]};
	ConfigRegister_32_8_32_1 config_reg_1(
		.clk(clk),
		.reset(reset),
		.O(config_reg_1_O),
		.config_addr(config_reg_1_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_2_config_addr;
	assign config_reg_2_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4], self_config_config_addr_out[3], self_config_config_addr_out[2:0]};
	ConfigRegister_32_8_32_2 config_reg_2(
		.clk(clk),
		.reset(reset),
		.O(config_reg_2_O),
		.config_addr(config_reg_2_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_3_config_addr;
	assign config_reg_3_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4], self_config_config_addr_out[3], self_config_config_addr_out[2:0]};
	ConfigRegister_31_8_32_3 config_reg_3(
		.clk(clk),
		.reset(reset),
		.O(config_reg_3_O),
		.config_addr(config_reg_3_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_4_config_addr;
	assign config_reg_4_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4], self_config_config_addr_out[3], self_config_config_addr_out[2:0]};
	ConfigRegister_30_8_32_4 config_reg_4(
		.clk(clk),
		.reset(reset),
		.O(config_reg_4_O),
		.config_addr(config_reg_4_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_5_config_addr;
	assign config_reg_5_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4], self_config_config_addr_out[3], self_config_config_addr_out[2:0]};
	ConfigRegister_23_8_32_5 config_reg_5(
		.clk(clk),
		.reset(reset),
		.O(config_reg_5_O),
		.config_addr(config_reg_5_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	coreir_const #(
		.value(1'h0),
		.width(1)
	) const_0_1(.out(const_0_1_out));
	coreir_const #(
		.value(32'h00000000),
		.width(32)
	) const_0_32(.out(const_0_32_out));
	coreir_const #(
		.value(1'h1),
		.width(1)
	) const_1_1(.out(const_1_1_out));
	coreir_eq #(.width(1)) coreir_eq_1_inst0(
		.in0(const_1_1_out),
		.in1(RMUX_T0_NORTH_B1_sel_value_O),
		.out(coreir_eq_1_inst0_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst1(
		.in0(const_1_1_out),
		.in1(RMUX_T0_SOUTH_B1_sel_value_O),
		.out(coreir_eq_1_inst1_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst10(
		.in0(const_1_1_out),
		.in1(RMUX_T2_EAST_B1_sel_value_O),
		.out(coreir_eq_1_inst10_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst11(
		.in0(const_1_1_out),
		.in1(RMUX_T2_WEST_B1_sel_value_O),
		.out(coreir_eq_1_inst11_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst12(
		.in0(const_1_1_out),
		.in1(RMUX_T3_NORTH_B1_sel_value_O),
		.out(coreir_eq_1_inst12_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst13(
		.in0(const_1_1_out),
		.in1(RMUX_T3_SOUTH_B1_sel_value_O),
		.out(coreir_eq_1_inst13_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst14(
		.in0(const_1_1_out),
		.in1(RMUX_T3_EAST_B1_sel_value_O),
		.out(coreir_eq_1_inst14_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst15(
		.in0(const_1_1_out),
		.in1(RMUX_T3_WEST_B1_sel_value_O),
		.out(coreir_eq_1_inst15_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst16(
		.in0(const_1_1_out),
		.in1(RMUX_T4_NORTH_B1_sel_value_O),
		.out(coreir_eq_1_inst16_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst17(
		.in0(const_1_1_out),
		.in1(RMUX_T4_SOUTH_B1_sel_value_O),
		.out(coreir_eq_1_inst17_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst18(
		.in0(const_1_1_out),
		.in1(RMUX_T4_EAST_B1_sel_value_O),
		.out(coreir_eq_1_inst18_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst19(
		.in0(const_1_1_out),
		.in1(RMUX_T4_WEST_B1_sel_value_O),
		.out(coreir_eq_1_inst19_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst2(
		.in0(const_1_1_out),
		.in1(RMUX_T0_EAST_B1_sel_value_O),
		.out(coreir_eq_1_inst2_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst3(
		.in0(const_1_1_out),
		.in1(RMUX_T0_WEST_B1_sel_value_O),
		.out(coreir_eq_1_inst3_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst4(
		.in0(const_1_1_out),
		.in1(RMUX_T1_NORTH_B1_sel_value_O),
		.out(coreir_eq_1_inst4_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst5(
		.in0(const_1_1_out),
		.in1(RMUX_T1_SOUTH_B1_sel_value_O),
		.out(coreir_eq_1_inst5_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst6(
		.in0(const_1_1_out),
		.in1(RMUX_T1_EAST_B1_sel_value_O),
		.out(coreir_eq_1_inst6_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst7(
		.in0(const_1_1_out),
		.in1(RMUX_T1_WEST_B1_sel_value_O),
		.out(coreir_eq_1_inst7_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst8(
		.in0(const_1_1_out),
		.in1(RMUX_T2_NORTH_B1_sel_value_O),
		.out(coreir_eq_1_inst8_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst9(
		.in0(const_1_1_out),
		.in1(RMUX_T2_SOUTH_B1_sel_value_O),
		.out(coreir_eq_1_inst9_out)
	);
	wire [191:0] mux_aoi_6_32_inst0_I;
	assign mux_aoi_6_32_inst0_I[160+:32] = ZextWrapper_23_32_inst0$self_O_in;
	assign mux_aoi_6_32_inst0_I[128+:32] = ZextWrapper_30_32_inst0$self_O_in;
	assign mux_aoi_6_32_inst0_I[96+:32] = ZextWrapper_31_32_inst0$self_O_in;
	assign mux_aoi_6_32_inst0_I[64+:32] = config_reg_2_O;
	assign mux_aoi_6_32_inst0_I[32+:32] = config_reg_1_O;
	assign mux_aoi_6_32_inst0_I[0+:32] = config_reg_0_O;
	mux_aoi_6_32 mux_aoi_6_32_inst0(
		.I(mux_aoi_6_32_inst0_I),
		.O(mux_aoi_6_32_inst0_O),
		.S(self_config_config_addr_out[2:0]),
		.out_sel(mux_aoi_6_32_inst0_out_sel)
	);
	mantle_wire__typeBit8 self_config_config_addr(
		.in(config_config_addr),
		.out(self_config_config_addr_out)
	);
	assign MEM_output_width_1_num_0_ready_out = CB_MEM_output_width_1_num_0_fan_in_O[0];
	assign MEM_output_width_1_num_1_ready_out = CB_MEM_output_width_1_num_1_fan_in_O[0];
	assign MEM_output_width_1_num_2_ready_out = CB_MEM_output_width_1_num_2_fan_in_O[0];
	assign SB_T0_EAST_SB_IN_B1_enable = SB_T0_EAST_SB_IN_B1_enable_value_O[0];
	assign SB_T0_EAST_SB_IN_B1_ready_out = WIRE_SB_T0_EAST_SB_IN_B1_ready_out;
	assign SB_T0_EAST_SB_OUT_B1 = RMUX_T0_EAST_B1_O;
	assign SB_T0_EAST_SB_OUT_B1_enable = SB_T0_EAST_SB_OUT_B1_enable_value_O[0];
	assign SB_T0_EAST_SB_OUT_B1_valid_out = RMUX_T0_EAST_B1_valid_out;
	assign SB_T0_NORTH_SB_IN_B1_enable = SB_T0_NORTH_SB_IN_B1_enable_value_O[0];
	assign SB_T0_NORTH_SB_IN_B1_ready_out = WIRE_SB_T0_NORTH_SB_IN_B1_ready_out;
	assign SB_T0_NORTH_SB_OUT_B1 = RMUX_T0_NORTH_B1_O;
	assign SB_T0_NORTH_SB_OUT_B1_enable = SB_T0_NORTH_SB_OUT_B1_enable_value_O[0];
	assign SB_T0_NORTH_SB_OUT_B1_valid_out = RMUX_T0_NORTH_B1_valid_out;
	assign SB_T0_SOUTH_SB_IN_B1_enable = SB_T0_SOUTH_SB_IN_B1_enable_value_O[0];
	assign SB_T0_SOUTH_SB_IN_B1_ready_out = WIRE_SB_T0_SOUTH_SB_IN_B1_ready_out;
	assign SB_T0_SOUTH_SB_OUT_B1 = RMUX_T0_SOUTH_B1_O;
	assign SB_T0_SOUTH_SB_OUT_B1_enable = SB_T0_SOUTH_SB_OUT_B1_enable_value_O[0];
	assign SB_T0_SOUTH_SB_OUT_B1_valid_out = RMUX_T0_SOUTH_B1_valid_out;
	assign SB_T0_WEST_SB_IN_B1_enable = SB_T0_WEST_SB_IN_B1_enable_value_O[0];
	assign SB_T0_WEST_SB_IN_B1_ready_out = WIRE_SB_T0_WEST_SB_IN_B1_ready_out;
	assign SB_T0_WEST_SB_OUT_B1 = RMUX_T0_WEST_B1_O;
	assign SB_T0_WEST_SB_OUT_B1_enable = SB_T0_WEST_SB_OUT_B1_enable_value_O[0];
	assign SB_T0_WEST_SB_OUT_B1_valid_out = RMUX_T0_WEST_B1_valid_out;
	assign SB_T1_EAST_SB_IN_B1_enable = SB_T1_EAST_SB_IN_B1_enable_value_O[0];
	assign SB_T1_EAST_SB_IN_B1_ready_out = WIRE_SB_T1_EAST_SB_IN_B1_ready_out;
	assign SB_T1_EAST_SB_OUT_B1 = RMUX_T1_EAST_B1_O;
	assign SB_T1_EAST_SB_OUT_B1_enable = SB_T1_EAST_SB_OUT_B1_enable_value_O[0];
	assign SB_T1_EAST_SB_OUT_B1_valid_out = RMUX_T1_EAST_B1_valid_out;
	assign SB_T1_NORTH_SB_IN_B1_enable = SB_T1_NORTH_SB_IN_B1_enable_value_O[0];
	assign SB_T1_NORTH_SB_IN_B1_ready_out = WIRE_SB_T1_NORTH_SB_IN_B1_ready_out;
	assign SB_T1_NORTH_SB_OUT_B1 = RMUX_T1_NORTH_B1_O;
	assign SB_T1_NORTH_SB_OUT_B1_enable = SB_T1_NORTH_SB_OUT_B1_enable_value_O[0];
	assign SB_T1_NORTH_SB_OUT_B1_valid_out = RMUX_T1_NORTH_B1_valid_out;
	assign SB_T1_SOUTH_SB_IN_B1_enable = SB_T1_SOUTH_SB_IN_B1_enable_value_O[0];
	assign SB_T1_SOUTH_SB_IN_B1_ready_out = WIRE_SB_T1_SOUTH_SB_IN_B1_ready_out;
	assign SB_T1_SOUTH_SB_OUT_B1 = RMUX_T1_SOUTH_B1_O;
	assign SB_T1_SOUTH_SB_OUT_B1_enable = SB_T1_SOUTH_SB_OUT_B1_enable_value_O[0];
	assign SB_T1_SOUTH_SB_OUT_B1_valid_out = RMUX_T1_SOUTH_B1_valid_out;
	assign SB_T1_WEST_SB_IN_B1_enable = SB_T1_WEST_SB_IN_B1_enable_value_O[0];
	assign SB_T1_WEST_SB_IN_B1_ready_out = WIRE_SB_T1_WEST_SB_IN_B1_ready_out;
	assign SB_T1_WEST_SB_OUT_B1 = RMUX_T1_WEST_B1_O;
	assign SB_T1_WEST_SB_OUT_B1_enable = SB_T1_WEST_SB_OUT_B1_enable_value_O[0];
	assign SB_T1_WEST_SB_OUT_B1_valid_out = RMUX_T1_WEST_B1_valid_out;
	assign SB_T2_EAST_SB_IN_B1_enable = SB_T2_EAST_SB_IN_B1_enable_value_O[0];
	assign SB_T2_EAST_SB_IN_B1_ready_out = WIRE_SB_T2_EAST_SB_IN_B1_ready_out;
	assign SB_T2_EAST_SB_OUT_B1 = RMUX_T2_EAST_B1_O;
	assign SB_T2_EAST_SB_OUT_B1_enable = SB_T2_EAST_SB_OUT_B1_enable_value_O[0];
	assign SB_T2_EAST_SB_OUT_B1_valid_out = RMUX_T2_EAST_B1_valid_out;
	assign SB_T2_NORTH_SB_IN_B1_enable = SB_T2_NORTH_SB_IN_B1_enable_value_O[0];
	assign SB_T2_NORTH_SB_IN_B1_ready_out = WIRE_SB_T2_NORTH_SB_IN_B1_ready_out;
	assign SB_T2_NORTH_SB_OUT_B1 = RMUX_T2_NORTH_B1_O;
	assign SB_T2_NORTH_SB_OUT_B1_enable = SB_T2_NORTH_SB_OUT_B1_enable_value_O[0];
	assign SB_T2_NORTH_SB_OUT_B1_valid_out = RMUX_T2_NORTH_B1_valid_out;
	assign SB_T2_SOUTH_SB_IN_B1_enable = SB_T2_SOUTH_SB_IN_B1_enable_value_O[0];
	assign SB_T2_SOUTH_SB_IN_B1_ready_out = WIRE_SB_T2_SOUTH_SB_IN_B1_ready_out;
	assign SB_T2_SOUTH_SB_OUT_B1 = RMUX_T2_SOUTH_B1_O;
	assign SB_T2_SOUTH_SB_OUT_B1_enable = SB_T2_SOUTH_SB_OUT_B1_enable_value_O[0];
	assign SB_T2_SOUTH_SB_OUT_B1_valid_out = RMUX_T2_SOUTH_B1_valid_out;
	assign SB_T2_WEST_SB_IN_B1_enable = SB_T2_WEST_SB_IN_B1_enable_value_O[0];
	assign SB_T2_WEST_SB_IN_B1_ready_out = WIRE_SB_T2_WEST_SB_IN_B1_ready_out;
	assign SB_T2_WEST_SB_OUT_B1 = RMUX_T2_WEST_B1_O;
	assign SB_T2_WEST_SB_OUT_B1_enable = SB_T2_WEST_SB_OUT_B1_enable_value_O[0];
	assign SB_T2_WEST_SB_OUT_B1_valid_out = RMUX_T2_WEST_B1_valid_out;
	assign SB_T3_EAST_SB_IN_B1_enable = SB_T3_EAST_SB_IN_B1_enable_value_O[0];
	assign SB_T3_EAST_SB_IN_B1_ready_out = WIRE_SB_T3_EAST_SB_IN_B1_ready_out;
	assign SB_T3_EAST_SB_OUT_B1 = RMUX_T3_EAST_B1_O;
	assign SB_T3_EAST_SB_OUT_B1_enable = SB_T3_EAST_SB_OUT_B1_enable_value_O[0];
	assign SB_T3_EAST_SB_OUT_B1_valid_out = RMUX_T3_EAST_B1_valid_out;
	assign SB_T3_NORTH_SB_IN_B1_enable = SB_T3_NORTH_SB_IN_B1_enable_value_O[0];
	assign SB_T3_NORTH_SB_IN_B1_ready_out = WIRE_SB_T3_NORTH_SB_IN_B1_ready_out;
	assign SB_T3_NORTH_SB_OUT_B1 = RMUX_T3_NORTH_B1_O;
	assign SB_T3_NORTH_SB_OUT_B1_enable = SB_T3_NORTH_SB_OUT_B1_enable_value_O[0];
	assign SB_T3_NORTH_SB_OUT_B1_valid_out = RMUX_T3_NORTH_B1_valid_out;
	assign SB_T3_SOUTH_SB_IN_B1_enable = SB_T3_SOUTH_SB_IN_B1_enable_value_O[0];
	assign SB_T3_SOUTH_SB_IN_B1_ready_out = WIRE_SB_T3_SOUTH_SB_IN_B1_ready_out;
	assign SB_T3_SOUTH_SB_OUT_B1 = RMUX_T3_SOUTH_B1_O;
	assign SB_T3_SOUTH_SB_OUT_B1_enable = SB_T3_SOUTH_SB_OUT_B1_enable_value_O[0];
	assign SB_T3_SOUTH_SB_OUT_B1_valid_out = RMUX_T3_SOUTH_B1_valid_out;
	assign SB_T3_WEST_SB_IN_B1_enable = SB_T3_WEST_SB_IN_B1_enable_value_O[0];
	assign SB_T3_WEST_SB_IN_B1_ready_out = WIRE_SB_T3_WEST_SB_IN_B1_ready_out;
	assign SB_T3_WEST_SB_OUT_B1 = RMUX_T3_WEST_B1_O;
	assign SB_T3_WEST_SB_OUT_B1_enable = SB_T3_WEST_SB_OUT_B1_enable_value_O[0];
	assign SB_T3_WEST_SB_OUT_B1_valid_out = RMUX_T3_WEST_B1_valid_out;
	assign SB_T4_EAST_SB_IN_B1_enable = SB_T4_EAST_SB_IN_B1_enable_value_O[0];
	assign SB_T4_EAST_SB_IN_B1_ready_out = WIRE_SB_T4_EAST_SB_IN_B1_ready_out;
	assign SB_T4_EAST_SB_OUT_B1 = RMUX_T4_EAST_B1_O;
	assign SB_T4_EAST_SB_OUT_B1_enable = SB_T4_EAST_SB_OUT_B1_enable_value_O[0];
	assign SB_T4_EAST_SB_OUT_B1_valid_out = RMUX_T4_EAST_B1_valid_out;
	assign SB_T4_NORTH_SB_IN_B1_enable = SB_T4_NORTH_SB_IN_B1_enable_value_O[0];
	assign SB_T4_NORTH_SB_IN_B1_ready_out = WIRE_SB_T4_NORTH_SB_IN_B1_ready_out;
	assign SB_T4_NORTH_SB_OUT_B1 = RMUX_T4_NORTH_B1_O;
	assign SB_T4_NORTH_SB_OUT_B1_enable = SB_T4_NORTH_SB_OUT_B1_enable_value_O[0];
	assign SB_T4_NORTH_SB_OUT_B1_valid_out = RMUX_T4_NORTH_B1_valid_out;
	assign SB_T4_SOUTH_SB_IN_B1_enable = SB_T4_SOUTH_SB_IN_B1_enable_value_O[0];
	assign SB_T4_SOUTH_SB_IN_B1_ready_out = WIRE_SB_T4_SOUTH_SB_IN_B1_ready_out;
	assign SB_T4_SOUTH_SB_OUT_B1 = RMUX_T4_SOUTH_B1_O;
	assign SB_T4_SOUTH_SB_OUT_B1_enable = SB_T4_SOUTH_SB_OUT_B1_enable_value_O[0];
	assign SB_T4_SOUTH_SB_OUT_B1_valid_out = RMUX_T4_SOUTH_B1_valid_out;
	assign SB_T4_WEST_SB_IN_B1_enable = SB_T4_WEST_SB_IN_B1_enable_value_O[0];
	assign SB_T4_WEST_SB_IN_B1_ready_out = WIRE_SB_T4_WEST_SB_IN_B1_ready_out;
	assign SB_T4_WEST_SB_OUT_B1 = RMUX_T4_WEST_B1_O;
	assign SB_T4_WEST_SB_OUT_B1_enable = SB_T4_WEST_SB_OUT_B1_enable_value_O[0];
	assign SB_T4_WEST_SB_OUT_B1_valid_out = RMUX_T4_WEST_B1_valid_out;
	assign read_config_data = mux_aoi_6_32_inst0_O;
endmodule
module SB_ID0_5TRACKS_B17_PE (
	PE_input_width_17_num_0_enable,
	PE_input_width_17_num_0_out_sel,
	PE_input_width_17_num_0_ready,
	PE_input_width_17_num_1_enable,
	PE_input_width_17_num_1_out_sel,
	PE_input_width_17_num_1_ready,
	PE_input_width_17_num_2_enable,
	PE_input_width_17_num_2_out_sel,
	PE_input_width_17_num_2_ready,
	PE_input_width_17_num_3_enable,
	PE_input_width_17_num_3_out_sel,
	PE_input_width_17_num_3_ready,
	PE_output_width_17_num_0,
	PE_output_width_17_num_0_ready_out,
	PE_output_width_17_num_0_valid,
	PE_output_width_17_num_1,
	PE_output_width_17_num_1_ready_out,
	PE_output_width_17_num_1_valid,
	PE_output_width_17_num_2,
	PE_output_width_17_num_2_ready_out,
	PE_output_width_17_num_2_valid,
	PondTop_input_width_17_num_0_enable,
	PondTop_input_width_17_num_0_out_sel,
	PondTop_input_width_17_num_0_ready,
	PondTop_input_width_17_num_1_enable,
	PondTop_input_width_17_num_1_out_sel,
	PondTop_input_width_17_num_1_ready,
	PondTop_output_width_17_num_0_ready_out,
	PondTop_output_width_17_num_0_valid,
	PondTop_output_width_17_num_1,
	PondTop_output_width_17_num_1_ready_out,
	PondTop_output_width_17_num_1_valid,
	SB_T0_EAST_SB_IN_B17,
	SB_T0_EAST_SB_IN_B17_enable,
	SB_T0_EAST_SB_IN_B17_ready_out,
	SB_T0_EAST_SB_IN_B17_valid_in,
	SB_T0_EAST_SB_OUT_B17,
	SB_T0_EAST_SB_OUT_B17_enable,
	SB_T0_EAST_SB_OUT_B17_ready_in,
	SB_T0_EAST_SB_OUT_B17_valid_out,
	SB_T0_NORTH_SB_IN_B17,
	SB_T0_NORTH_SB_IN_B17_enable,
	SB_T0_NORTH_SB_IN_B17_ready_out,
	SB_T0_NORTH_SB_IN_B17_valid_in,
	SB_T0_NORTH_SB_OUT_B17,
	SB_T0_NORTH_SB_OUT_B17_enable,
	SB_T0_NORTH_SB_OUT_B17_ready_in,
	SB_T0_NORTH_SB_OUT_B17_valid_out,
	SB_T0_SOUTH_SB_IN_B17,
	SB_T0_SOUTH_SB_IN_B17_enable,
	SB_T0_SOUTH_SB_IN_B17_ready_out,
	SB_T0_SOUTH_SB_IN_B17_valid_in,
	SB_T0_SOUTH_SB_OUT_B17,
	SB_T0_SOUTH_SB_OUT_B17_enable,
	SB_T0_SOUTH_SB_OUT_B17_ready_in,
	SB_T0_SOUTH_SB_OUT_B17_valid_out,
	SB_T0_WEST_SB_IN_B17,
	SB_T0_WEST_SB_IN_B17_enable,
	SB_T0_WEST_SB_IN_B17_ready_out,
	SB_T0_WEST_SB_IN_B17_valid_in,
	SB_T0_WEST_SB_OUT_B17,
	SB_T0_WEST_SB_OUT_B17_enable,
	SB_T0_WEST_SB_OUT_B17_ready_in,
	SB_T0_WEST_SB_OUT_B17_valid_out,
	SB_T1_EAST_SB_IN_B17,
	SB_T1_EAST_SB_IN_B17_enable,
	SB_T1_EAST_SB_IN_B17_ready_out,
	SB_T1_EAST_SB_IN_B17_valid_in,
	SB_T1_EAST_SB_OUT_B17,
	SB_T1_EAST_SB_OUT_B17_enable,
	SB_T1_EAST_SB_OUT_B17_ready_in,
	SB_T1_EAST_SB_OUT_B17_valid_out,
	SB_T1_NORTH_SB_IN_B17,
	SB_T1_NORTH_SB_IN_B17_enable,
	SB_T1_NORTH_SB_IN_B17_ready_out,
	SB_T1_NORTH_SB_IN_B17_valid_in,
	SB_T1_NORTH_SB_OUT_B17,
	SB_T1_NORTH_SB_OUT_B17_enable,
	SB_T1_NORTH_SB_OUT_B17_ready_in,
	SB_T1_NORTH_SB_OUT_B17_valid_out,
	SB_T1_SOUTH_SB_IN_B17,
	SB_T1_SOUTH_SB_IN_B17_enable,
	SB_T1_SOUTH_SB_IN_B17_ready_out,
	SB_T1_SOUTH_SB_IN_B17_valid_in,
	SB_T1_SOUTH_SB_OUT_B17,
	SB_T1_SOUTH_SB_OUT_B17_enable,
	SB_T1_SOUTH_SB_OUT_B17_ready_in,
	SB_T1_SOUTH_SB_OUT_B17_valid_out,
	SB_T1_WEST_SB_IN_B17,
	SB_T1_WEST_SB_IN_B17_enable,
	SB_T1_WEST_SB_IN_B17_ready_out,
	SB_T1_WEST_SB_IN_B17_valid_in,
	SB_T1_WEST_SB_OUT_B17,
	SB_T1_WEST_SB_OUT_B17_enable,
	SB_T1_WEST_SB_OUT_B17_ready_in,
	SB_T1_WEST_SB_OUT_B17_valid_out,
	SB_T2_EAST_SB_IN_B17,
	SB_T2_EAST_SB_IN_B17_enable,
	SB_T2_EAST_SB_IN_B17_ready_out,
	SB_T2_EAST_SB_IN_B17_valid_in,
	SB_T2_EAST_SB_OUT_B17,
	SB_T2_EAST_SB_OUT_B17_enable,
	SB_T2_EAST_SB_OUT_B17_ready_in,
	SB_T2_EAST_SB_OUT_B17_valid_out,
	SB_T2_NORTH_SB_IN_B17,
	SB_T2_NORTH_SB_IN_B17_enable,
	SB_T2_NORTH_SB_IN_B17_ready_out,
	SB_T2_NORTH_SB_IN_B17_valid_in,
	SB_T2_NORTH_SB_OUT_B17,
	SB_T2_NORTH_SB_OUT_B17_enable,
	SB_T2_NORTH_SB_OUT_B17_ready_in,
	SB_T2_NORTH_SB_OUT_B17_valid_out,
	SB_T2_SOUTH_SB_IN_B17,
	SB_T2_SOUTH_SB_IN_B17_enable,
	SB_T2_SOUTH_SB_IN_B17_ready_out,
	SB_T2_SOUTH_SB_IN_B17_valid_in,
	SB_T2_SOUTH_SB_OUT_B17,
	SB_T2_SOUTH_SB_OUT_B17_enable,
	SB_T2_SOUTH_SB_OUT_B17_ready_in,
	SB_T2_SOUTH_SB_OUT_B17_valid_out,
	SB_T2_WEST_SB_IN_B17,
	SB_T2_WEST_SB_IN_B17_enable,
	SB_T2_WEST_SB_IN_B17_ready_out,
	SB_T2_WEST_SB_IN_B17_valid_in,
	SB_T2_WEST_SB_OUT_B17,
	SB_T2_WEST_SB_OUT_B17_enable,
	SB_T2_WEST_SB_OUT_B17_ready_in,
	SB_T2_WEST_SB_OUT_B17_valid_out,
	SB_T3_EAST_SB_IN_B17,
	SB_T3_EAST_SB_IN_B17_enable,
	SB_T3_EAST_SB_IN_B17_ready_out,
	SB_T3_EAST_SB_IN_B17_valid_in,
	SB_T3_EAST_SB_OUT_B17,
	SB_T3_EAST_SB_OUT_B17_enable,
	SB_T3_EAST_SB_OUT_B17_ready_in,
	SB_T3_EAST_SB_OUT_B17_valid_out,
	SB_T3_NORTH_SB_IN_B17,
	SB_T3_NORTH_SB_IN_B17_enable,
	SB_T3_NORTH_SB_IN_B17_ready_out,
	SB_T3_NORTH_SB_IN_B17_valid_in,
	SB_T3_NORTH_SB_OUT_B17,
	SB_T3_NORTH_SB_OUT_B17_enable,
	SB_T3_NORTH_SB_OUT_B17_ready_in,
	SB_T3_NORTH_SB_OUT_B17_valid_out,
	SB_T3_SOUTH_SB_IN_B17,
	SB_T3_SOUTH_SB_IN_B17_enable,
	SB_T3_SOUTH_SB_IN_B17_ready_out,
	SB_T3_SOUTH_SB_IN_B17_valid_in,
	SB_T3_SOUTH_SB_OUT_B17,
	SB_T3_SOUTH_SB_OUT_B17_enable,
	SB_T3_SOUTH_SB_OUT_B17_ready_in,
	SB_T3_SOUTH_SB_OUT_B17_valid_out,
	SB_T3_WEST_SB_IN_B17,
	SB_T3_WEST_SB_IN_B17_enable,
	SB_T3_WEST_SB_IN_B17_ready_out,
	SB_T3_WEST_SB_IN_B17_valid_in,
	SB_T3_WEST_SB_OUT_B17,
	SB_T3_WEST_SB_OUT_B17_enable,
	SB_T3_WEST_SB_OUT_B17_ready_in,
	SB_T3_WEST_SB_OUT_B17_valid_out,
	SB_T4_EAST_SB_IN_B17,
	SB_T4_EAST_SB_IN_B17_enable,
	SB_T4_EAST_SB_IN_B17_ready_out,
	SB_T4_EAST_SB_IN_B17_valid_in,
	SB_T4_EAST_SB_OUT_B17,
	SB_T4_EAST_SB_OUT_B17_enable,
	SB_T4_EAST_SB_OUT_B17_ready_in,
	SB_T4_EAST_SB_OUT_B17_valid_out,
	SB_T4_NORTH_SB_IN_B17,
	SB_T4_NORTH_SB_IN_B17_enable,
	SB_T4_NORTH_SB_IN_B17_ready_out,
	SB_T4_NORTH_SB_IN_B17_valid_in,
	SB_T4_NORTH_SB_OUT_B17,
	SB_T4_NORTH_SB_OUT_B17_enable,
	SB_T4_NORTH_SB_OUT_B17_ready_in,
	SB_T4_NORTH_SB_OUT_B17_valid_out,
	SB_T4_SOUTH_SB_IN_B17,
	SB_T4_SOUTH_SB_IN_B17_enable,
	SB_T4_SOUTH_SB_IN_B17_ready_out,
	SB_T4_SOUTH_SB_IN_B17_valid_in,
	SB_T4_SOUTH_SB_OUT_B17,
	SB_T4_SOUTH_SB_OUT_B17_enable,
	SB_T4_SOUTH_SB_OUT_B17_ready_in,
	SB_T4_SOUTH_SB_OUT_B17_valid_out,
	SB_T4_WEST_SB_IN_B17,
	SB_T4_WEST_SB_IN_B17_enable,
	SB_T4_WEST_SB_IN_B17_ready_out,
	SB_T4_WEST_SB_IN_B17_valid_in,
	SB_T4_WEST_SB_OUT_B17,
	SB_T4_WEST_SB_OUT_B17_enable,
	SB_T4_WEST_SB_OUT_B17_ready_in,
	SB_T4_WEST_SB_OUT_B17_valid_out,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	read_config_data,
	reset,
	stall
);
	input [0:0] PE_input_width_17_num_0_enable;
	input [31:0] PE_input_width_17_num_0_out_sel;
	input PE_input_width_17_num_0_ready;
	input [0:0] PE_input_width_17_num_1_enable;
	input [31:0] PE_input_width_17_num_1_out_sel;
	input PE_input_width_17_num_1_ready;
	input [0:0] PE_input_width_17_num_2_enable;
	input [31:0] PE_input_width_17_num_2_out_sel;
	input PE_input_width_17_num_2_ready;
	input [0:0] PE_input_width_17_num_3_enable;
	input [31:0] PE_input_width_17_num_3_out_sel;
	input PE_input_width_17_num_3_ready;
	input [16:0] PE_output_width_17_num_0;
	output wire PE_output_width_17_num_0_ready_out;
	input PE_output_width_17_num_0_valid;
	input [16:0] PE_output_width_17_num_1;
	output wire PE_output_width_17_num_1_ready_out;
	input PE_output_width_17_num_1_valid;
	input [16:0] PE_output_width_17_num_2;
	output wire PE_output_width_17_num_2_ready_out;
	input PE_output_width_17_num_2_valid;
	input [0:0] PondTop_input_width_17_num_0_enable;
	input [31:0] PondTop_input_width_17_num_0_out_sel;
	input PondTop_input_width_17_num_0_ready;
	input [0:0] PondTop_input_width_17_num_1_enable;
	input [31:0] PondTop_input_width_17_num_1_out_sel;
	input PondTop_input_width_17_num_1_ready;
	output wire PondTop_output_width_17_num_0_ready_out;
	input PondTop_output_width_17_num_0_valid;
	input [16:0] PondTop_output_width_17_num_1;
	output wire PondTop_output_width_17_num_1_ready_out;
	input PondTop_output_width_17_num_1_valid;
	input [16:0] SB_T0_EAST_SB_IN_B17;
	output wire SB_T0_EAST_SB_IN_B17_enable;
	output wire SB_T0_EAST_SB_IN_B17_ready_out;
	input SB_T0_EAST_SB_IN_B17_valid_in;
	output wire [16:0] SB_T0_EAST_SB_OUT_B17;
	output wire SB_T0_EAST_SB_OUT_B17_enable;
	input SB_T0_EAST_SB_OUT_B17_ready_in;
	output wire SB_T0_EAST_SB_OUT_B17_valid_out;
	input [16:0] SB_T0_NORTH_SB_IN_B17;
	output wire SB_T0_NORTH_SB_IN_B17_enable;
	output wire SB_T0_NORTH_SB_IN_B17_ready_out;
	input SB_T0_NORTH_SB_IN_B17_valid_in;
	output wire [16:0] SB_T0_NORTH_SB_OUT_B17;
	output wire SB_T0_NORTH_SB_OUT_B17_enable;
	input SB_T0_NORTH_SB_OUT_B17_ready_in;
	output wire SB_T0_NORTH_SB_OUT_B17_valid_out;
	input [16:0] SB_T0_SOUTH_SB_IN_B17;
	output wire SB_T0_SOUTH_SB_IN_B17_enable;
	output wire SB_T0_SOUTH_SB_IN_B17_ready_out;
	input SB_T0_SOUTH_SB_IN_B17_valid_in;
	output wire [16:0] SB_T0_SOUTH_SB_OUT_B17;
	output wire SB_T0_SOUTH_SB_OUT_B17_enable;
	input SB_T0_SOUTH_SB_OUT_B17_ready_in;
	output wire SB_T0_SOUTH_SB_OUT_B17_valid_out;
	input [16:0] SB_T0_WEST_SB_IN_B17;
	output wire SB_T0_WEST_SB_IN_B17_enable;
	output wire SB_T0_WEST_SB_IN_B17_ready_out;
	input SB_T0_WEST_SB_IN_B17_valid_in;
	output wire [16:0] SB_T0_WEST_SB_OUT_B17;
	output wire SB_T0_WEST_SB_OUT_B17_enable;
	input SB_T0_WEST_SB_OUT_B17_ready_in;
	output wire SB_T0_WEST_SB_OUT_B17_valid_out;
	input [16:0] SB_T1_EAST_SB_IN_B17;
	output wire SB_T1_EAST_SB_IN_B17_enable;
	output wire SB_T1_EAST_SB_IN_B17_ready_out;
	input SB_T1_EAST_SB_IN_B17_valid_in;
	output wire [16:0] SB_T1_EAST_SB_OUT_B17;
	output wire SB_T1_EAST_SB_OUT_B17_enable;
	input SB_T1_EAST_SB_OUT_B17_ready_in;
	output wire SB_T1_EAST_SB_OUT_B17_valid_out;
	input [16:0] SB_T1_NORTH_SB_IN_B17;
	output wire SB_T1_NORTH_SB_IN_B17_enable;
	output wire SB_T1_NORTH_SB_IN_B17_ready_out;
	input SB_T1_NORTH_SB_IN_B17_valid_in;
	output wire [16:0] SB_T1_NORTH_SB_OUT_B17;
	output wire SB_T1_NORTH_SB_OUT_B17_enable;
	input SB_T1_NORTH_SB_OUT_B17_ready_in;
	output wire SB_T1_NORTH_SB_OUT_B17_valid_out;
	input [16:0] SB_T1_SOUTH_SB_IN_B17;
	output wire SB_T1_SOUTH_SB_IN_B17_enable;
	output wire SB_T1_SOUTH_SB_IN_B17_ready_out;
	input SB_T1_SOUTH_SB_IN_B17_valid_in;
	output wire [16:0] SB_T1_SOUTH_SB_OUT_B17;
	output wire SB_T1_SOUTH_SB_OUT_B17_enable;
	input SB_T1_SOUTH_SB_OUT_B17_ready_in;
	output wire SB_T1_SOUTH_SB_OUT_B17_valid_out;
	input [16:0] SB_T1_WEST_SB_IN_B17;
	output wire SB_T1_WEST_SB_IN_B17_enable;
	output wire SB_T1_WEST_SB_IN_B17_ready_out;
	input SB_T1_WEST_SB_IN_B17_valid_in;
	output wire [16:0] SB_T1_WEST_SB_OUT_B17;
	output wire SB_T1_WEST_SB_OUT_B17_enable;
	input SB_T1_WEST_SB_OUT_B17_ready_in;
	output wire SB_T1_WEST_SB_OUT_B17_valid_out;
	input [16:0] SB_T2_EAST_SB_IN_B17;
	output wire SB_T2_EAST_SB_IN_B17_enable;
	output wire SB_T2_EAST_SB_IN_B17_ready_out;
	input SB_T2_EAST_SB_IN_B17_valid_in;
	output wire [16:0] SB_T2_EAST_SB_OUT_B17;
	output wire SB_T2_EAST_SB_OUT_B17_enable;
	input SB_T2_EAST_SB_OUT_B17_ready_in;
	output wire SB_T2_EAST_SB_OUT_B17_valid_out;
	input [16:0] SB_T2_NORTH_SB_IN_B17;
	output wire SB_T2_NORTH_SB_IN_B17_enable;
	output wire SB_T2_NORTH_SB_IN_B17_ready_out;
	input SB_T2_NORTH_SB_IN_B17_valid_in;
	output wire [16:0] SB_T2_NORTH_SB_OUT_B17;
	output wire SB_T2_NORTH_SB_OUT_B17_enable;
	input SB_T2_NORTH_SB_OUT_B17_ready_in;
	output wire SB_T2_NORTH_SB_OUT_B17_valid_out;
	input [16:0] SB_T2_SOUTH_SB_IN_B17;
	output wire SB_T2_SOUTH_SB_IN_B17_enable;
	output wire SB_T2_SOUTH_SB_IN_B17_ready_out;
	input SB_T2_SOUTH_SB_IN_B17_valid_in;
	output wire [16:0] SB_T2_SOUTH_SB_OUT_B17;
	output wire SB_T2_SOUTH_SB_OUT_B17_enable;
	input SB_T2_SOUTH_SB_OUT_B17_ready_in;
	output wire SB_T2_SOUTH_SB_OUT_B17_valid_out;
	input [16:0] SB_T2_WEST_SB_IN_B17;
	output wire SB_T2_WEST_SB_IN_B17_enable;
	output wire SB_T2_WEST_SB_IN_B17_ready_out;
	input SB_T2_WEST_SB_IN_B17_valid_in;
	output wire [16:0] SB_T2_WEST_SB_OUT_B17;
	output wire SB_T2_WEST_SB_OUT_B17_enable;
	input SB_T2_WEST_SB_OUT_B17_ready_in;
	output wire SB_T2_WEST_SB_OUT_B17_valid_out;
	input [16:0] SB_T3_EAST_SB_IN_B17;
	output wire SB_T3_EAST_SB_IN_B17_enable;
	output wire SB_T3_EAST_SB_IN_B17_ready_out;
	input SB_T3_EAST_SB_IN_B17_valid_in;
	output wire [16:0] SB_T3_EAST_SB_OUT_B17;
	output wire SB_T3_EAST_SB_OUT_B17_enable;
	input SB_T3_EAST_SB_OUT_B17_ready_in;
	output wire SB_T3_EAST_SB_OUT_B17_valid_out;
	input [16:0] SB_T3_NORTH_SB_IN_B17;
	output wire SB_T3_NORTH_SB_IN_B17_enable;
	output wire SB_T3_NORTH_SB_IN_B17_ready_out;
	input SB_T3_NORTH_SB_IN_B17_valid_in;
	output wire [16:0] SB_T3_NORTH_SB_OUT_B17;
	output wire SB_T3_NORTH_SB_OUT_B17_enable;
	input SB_T3_NORTH_SB_OUT_B17_ready_in;
	output wire SB_T3_NORTH_SB_OUT_B17_valid_out;
	input [16:0] SB_T3_SOUTH_SB_IN_B17;
	output wire SB_T3_SOUTH_SB_IN_B17_enable;
	output wire SB_T3_SOUTH_SB_IN_B17_ready_out;
	input SB_T3_SOUTH_SB_IN_B17_valid_in;
	output wire [16:0] SB_T3_SOUTH_SB_OUT_B17;
	output wire SB_T3_SOUTH_SB_OUT_B17_enable;
	input SB_T3_SOUTH_SB_OUT_B17_ready_in;
	output wire SB_T3_SOUTH_SB_OUT_B17_valid_out;
	input [16:0] SB_T3_WEST_SB_IN_B17;
	output wire SB_T3_WEST_SB_IN_B17_enable;
	output wire SB_T3_WEST_SB_IN_B17_ready_out;
	input SB_T3_WEST_SB_IN_B17_valid_in;
	output wire [16:0] SB_T3_WEST_SB_OUT_B17;
	output wire SB_T3_WEST_SB_OUT_B17_enable;
	input SB_T3_WEST_SB_OUT_B17_ready_in;
	output wire SB_T3_WEST_SB_OUT_B17_valid_out;
	input [16:0] SB_T4_EAST_SB_IN_B17;
	output wire SB_T4_EAST_SB_IN_B17_enable;
	output wire SB_T4_EAST_SB_IN_B17_ready_out;
	input SB_T4_EAST_SB_IN_B17_valid_in;
	output wire [16:0] SB_T4_EAST_SB_OUT_B17;
	output wire SB_T4_EAST_SB_OUT_B17_enable;
	input SB_T4_EAST_SB_OUT_B17_ready_in;
	output wire SB_T4_EAST_SB_OUT_B17_valid_out;
	input [16:0] SB_T4_NORTH_SB_IN_B17;
	output wire SB_T4_NORTH_SB_IN_B17_enable;
	output wire SB_T4_NORTH_SB_IN_B17_ready_out;
	input SB_T4_NORTH_SB_IN_B17_valid_in;
	output wire [16:0] SB_T4_NORTH_SB_OUT_B17;
	output wire SB_T4_NORTH_SB_OUT_B17_enable;
	input SB_T4_NORTH_SB_OUT_B17_ready_in;
	output wire SB_T4_NORTH_SB_OUT_B17_valid_out;
	input [16:0] SB_T4_SOUTH_SB_IN_B17;
	output wire SB_T4_SOUTH_SB_IN_B17_enable;
	output wire SB_T4_SOUTH_SB_IN_B17_ready_out;
	input SB_T4_SOUTH_SB_IN_B17_valid_in;
	output wire [16:0] SB_T4_SOUTH_SB_OUT_B17;
	output wire SB_T4_SOUTH_SB_OUT_B17_enable;
	input SB_T4_SOUTH_SB_OUT_B17_ready_in;
	output wire SB_T4_SOUTH_SB_OUT_B17_valid_out;
	input [16:0] SB_T4_WEST_SB_IN_B17;
	output wire SB_T4_WEST_SB_IN_B17_enable;
	output wire SB_T4_WEST_SB_IN_B17_ready_out;
	input SB_T4_WEST_SB_IN_B17_valid_in;
	output wire [16:0] SB_T4_WEST_SB_OUT_B17;
	output wire SB_T4_WEST_SB_OUT_B17_enable;
	input SB_T4_WEST_SB_OUT_B17_ready_in;
	output wire SB_T4_WEST_SB_OUT_B17_valid_out;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output wire [31:0] read_config_data;
	input reset;
	input [0:0] stall;
	wire [0:0] CB_PE_output_width_17_num_0_fan_in_O;
	wire [0:0] CB_PE_output_width_17_num_1_fan_in_O;
	wire [0:0] CB_PE_output_width_17_num_2_fan_in_O;
	wire [0:0] CB_PondTop_output_width_17_num_0_fan_in_O;
	wire [0:0] CB_PondTop_output_width_17_num_1_fan_in_O;
	wire [0:0] Invert1_inst0_out;
	wire [16:0] MUX_SB_T0_EAST_SB_OUT_B17_O;
	wire MUX_SB_T0_EAST_SB_OUT_B17_ready_out;
	wire MUX_SB_T0_EAST_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T0_EAST_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T0_NORTH_SB_OUT_B17_O;
	wire MUX_SB_T0_NORTH_SB_OUT_B17_ready_out;
	wire MUX_SB_T0_NORTH_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T0_NORTH_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T0_SOUTH_SB_OUT_B17_O;
	wire MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out;
	wire MUX_SB_T0_SOUTH_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T0_WEST_SB_OUT_B17_O;
	wire MUX_SB_T0_WEST_SB_OUT_B17_ready_out;
	wire MUX_SB_T0_WEST_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T0_WEST_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T1_EAST_SB_OUT_B17_O;
	wire MUX_SB_T1_EAST_SB_OUT_B17_ready_out;
	wire MUX_SB_T1_EAST_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T1_EAST_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T1_NORTH_SB_OUT_B17_O;
	wire MUX_SB_T1_NORTH_SB_OUT_B17_ready_out;
	wire MUX_SB_T1_NORTH_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T1_NORTH_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T1_SOUTH_SB_OUT_B17_O;
	wire MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out;
	wire MUX_SB_T1_SOUTH_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T1_WEST_SB_OUT_B17_O;
	wire MUX_SB_T1_WEST_SB_OUT_B17_ready_out;
	wire MUX_SB_T1_WEST_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T1_WEST_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T2_EAST_SB_OUT_B17_O;
	wire MUX_SB_T2_EAST_SB_OUT_B17_ready_out;
	wire MUX_SB_T2_EAST_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T2_EAST_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T2_NORTH_SB_OUT_B17_O;
	wire MUX_SB_T2_NORTH_SB_OUT_B17_ready_out;
	wire MUX_SB_T2_NORTH_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T2_NORTH_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T2_SOUTH_SB_OUT_B17_O;
	wire MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out;
	wire MUX_SB_T2_SOUTH_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T2_WEST_SB_OUT_B17_O;
	wire MUX_SB_T2_WEST_SB_OUT_B17_ready_out;
	wire MUX_SB_T2_WEST_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T2_WEST_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T3_EAST_SB_OUT_B17_O;
	wire MUX_SB_T3_EAST_SB_OUT_B17_ready_out;
	wire MUX_SB_T3_EAST_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T3_EAST_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T3_NORTH_SB_OUT_B17_O;
	wire MUX_SB_T3_NORTH_SB_OUT_B17_ready_out;
	wire MUX_SB_T3_NORTH_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T3_NORTH_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T3_SOUTH_SB_OUT_B17_O;
	wire MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out;
	wire MUX_SB_T3_SOUTH_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T3_WEST_SB_OUT_B17_O;
	wire MUX_SB_T3_WEST_SB_OUT_B17_ready_out;
	wire MUX_SB_T3_WEST_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T3_WEST_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T4_EAST_SB_OUT_B17_O;
	wire MUX_SB_T4_EAST_SB_OUT_B17_ready_out;
	wire MUX_SB_T4_EAST_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T4_EAST_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T4_NORTH_SB_OUT_B17_O;
	wire MUX_SB_T4_NORTH_SB_OUT_B17_ready_out;
	wire MUX_SB_T4_NORTH_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T4_NORTH_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T4_SOUTH_SB_OUT_B17_O;
	wire MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out;
	wire MUX_SB_T4_SOUTH_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T4_WEST_SB_OUT_B17_O;
	wire MUX_SB_T4_WEST_SB_OUT_B17_ready_out;
	wire MUX_SB_T4_WEST_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T4_WEST_SB_OUT_B17_out_sel;
	wire [0:0] REG_T0_EAST_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T0_EAST_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T0_EAST_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T0_EAST_B17_end_value_O;
	wire [0:0] REG_T0_EAST_B17_fifo_value_O;
	wire [0:0] REG_T0_EAST_B17_start_value_O;
	wire [0:0] REG_T0_NORTH_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T0_NORTH_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T0_NORTH_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T0_NORTH_B17_end_value_O;
	wire [0:0] REG_T0_NORTH_B17_fifo_value_O;
	wire [0:0] REG_T0_NORTH_B17_start_value_O;
	wire [0:0] REG_T0_SOUTH_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T0_SOUTH_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T0_SOUTH_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T0_SOUTH_B17_end_value_O;
	wire [0:0] REG_T0_SOUTH_B17_fifo_value_O;
	wire [0:0] REG_T0_SOUTH_B17_start_value_O;
	wire [0:0] REG_T0_WEST_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T0_WEST_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T0_WEST_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T0_WEST_B17_end_value_O;
	wire [0:0] REG_T0_WEST_B17_fifo_value_O;
	wire [0:0] REG_T0_WEST_B17_start_value_O;
	wire [0:0] REG_T1_EAST_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T1_EAST_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T1_EAST_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T1_EAST_B17_end_value_O;
	wire [0:0] REG_T1_EAST_B17_fifo_value_O;
	wire [0:0] REG_T1_EAST_B17_start_value_O;
	wire [0:0] REG_T1_NORTH_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T1_NORTH_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T1_NORTH_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T1_NORTH_B17_end_value_O;
	wire [0:0] REG_T1_NORTH_B17_fifo_value_O;
	wire [0:0] REG_T1_NORTH_B17_start_value_O;
	wire [0:0] REG_T1_SOUTH_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T1_SOUTH_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T1_SOUTH_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T1_SOUTH_B17_end_value_O;
	wire [0:0] REG_T1_SOUTH_B17_fifo_value_O;
	wire [0:0] REG_T1_SOUTH_B17_start_value_O;
	wire [0:0] REG_T1_WEST_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T1_WEST_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T1_WEST_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T1_WEST_B17_end_value_O;
	wire [0:0] REG_T1_WEST_B17_fifo_value_O;
	wire [0:0] REG_T1_WEST_B17_start_value_O;
	wire [0:0] REG_T2_EAST_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T2_EAST_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T2_EAST_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T2_EAST_B17_end_value_O;
	wire [0:0] REG_T2_EAST_B17_fifo_value_O;
	wire [0:0] REG_T2_EAST_B17_start_value_O;
	wire [0:0] REG_T2_NORTH_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T2_NORTH_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T2_NORTH_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T2_NORTH_B17_end_value_O;
	wire [0:0] REG_T2_NORTH_B17_fifo_value_O;
	wire [0:0] REG_T2_NORTH_B17_start_value_O;
	wire [0:0] REG_T2_SOUTH_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T2_SOUTH_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T2_SOUTH_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T2_SOUTH_B17_end_value_O;
	wire [0:0] REG_T2_SOUTH_B17_fifo_value_O;
	wire [0:0] REG_T2_SOUTH_B17_start_value_O;
	wire [0:0] REG_T2_WEST_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T2_WEST_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T2_WEST_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T2_WEST_B17_end_value_O;
	wire [0:0] REG_T2_WEST_B17_fifo_value_O;
	wire [0:0] REG_T2_WEST_B17_start_value_O;
	wire [0:0] REG_T3_EAST_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T3_EAST_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T3_EAST_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T3_EAST_B17_end_value_O;
	wire [0:0] REG_T3_EAST_B17_fifo_value_O;
	wire [0:0] REG_T3_EAST_B17_start_value_O;
	wire [0:0] REG_T3_NORTH_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T3_NORTH_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T3_NORTH_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T3_NORTH_B17_end_value_O;
	wire [0:0] REG_T3_NORTH_B17_fifo_value_O;
	wire [0:0] REG_T3_NORTH_B17_start_value_O;
	wire [0:0] REG_T3_SOUTH_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T3_SOUTH_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T3_SOUTH_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T3_SOUTH_B17_end_value_O;
	wire [0:0] REG_T3_SOUTH_B17_fifo_value_O;
	wire [0:0] REG_T3_SOUTH_B17_start_value_O;
	wire [0:0] REG_T3_WEST_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T3_WEST_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T3_WEST_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T3_WEST_B17_end_value_O;
	wire [0:0] REG_T3_WEST_B17_fifo_value_O;
	wire [0:0] REG_T3_WEST_B17_start_value_O;
	wire [0:0] REG_T4_EAST_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T4_EAST_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T4_EAST_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T4_EAST_B17_end_value_O;
	wire [0:0] REG_T4_EAST_B17_fifo_value_O;
	wire [0:0] REG_T4_EAST_B17_start_value_O;
	wire [0:0] REG_T4_NORTH_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T4_NORTH_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T4_NORTH_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T4_NORTH_B17_end_value_O;
	wire [0:0] REG_T4_NORTH_B17_fifo_value_O;
	wire [0:0] REG_T4_NORTH_B17_start_value_O;
	wire [0:0] REG_T4_SOUTH_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T4_SOUTH_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T4_SOUTH_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T4_SOUTH_B17_end_value_O;
	wire [0:0] REG_T4_SOUTH_B17_fifo_value_O;
	wire [0:0] REG_T4_SOUTH_B17_start_value_O;
	wire [0:0] REG_T4_WEST_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T4_WEST_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T4_WEST_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T4_WEST_B17_end_value_O;
	wire [0:0] REG_T4_WEST_B17_fifo_value_O;
	wire [0:0] REG_T4_WEST_B17_start_value_O;
	wire [16:0] RMUX_T0_EAST_B17_O;
	wire RMUX_T0_EAST_B17_ready_out;
	wire RMUX_T0_EAST_B17_valid_out;
	wire [1:0] RMUX_T0_EAST_B17_out_sel;
	wire [0:0] RMUX_T0_EAST_B17_sel_value_O;
	wire [16:0] RMUX_T0_NORTH_B17_O;
	wire RMUX_T0_NORTH_B17_ready_out;
	wire RMUX_T0_NORTH_B17_valid_out;
	wire [1:0] RMUX_T0_NORTH_B17_out_sel;
	wire [0:0] RMUX_T0_NORTH_B17_sel_value_O;
	wire [16:0] RMUX_T0_SOUTH_B17_O;
	wire RMUX_T0_SOUTH_B17_ready_out;
	wire RMUX_T0_SOUTH_B17_valid_out;
	wire [1:0] RMUX_T0_SOUTH_B17_out_sel;
	wire [0:0] RMUX_T0_SOUTH_B17_sel_value_O;
	wire [16:0] RMUX_T0_WEST_B17_O;
	wire RMUX_T0_WEST_B17_ready_out;
	wire RMUX_T0_WEST_B17_valid_out;
	wire [1:0] RMUX_T0_WEST_B17_out_sel;
	wire [0:0] RMUX_T0_WEST_B17_sel_value_O;
	wire [16:0] RMUX_T1_EAST_B17_O;
	wire RMUX_T1_EAST_B17_ready_out;
	wire RMUX_T1_EAST_B17_valid_out;
	wire [1:0] RMUX_T1_EAST_B17_out_sel;
	wire [0:0] RMUX_T1_EAST_B17_sel_value_O;
	wire [16:0] RMUX_T1_NORTH_B17_O;
	wire RMUX_T1_NORTH_B17_ready_out;
	wire RMUX_T1_NORTH_B17_valid_out;
	wire [1:0] RMUX_T1_NORTH_B17_out_sel;
	wire [0:0] RMUX_T1_NORTH_B17_sel_value_O;
	wire [16:0] RMUX_T1_SOUTH_B17_O;
	wire RMUX_T1_SOUTH_B17_ready_out;
	wire RMUX_T1_SOUTH_B17_valid_out;
	wire [1:0] RMUX_T1_SOUTH_B17_out_sel;
	wire [0:0] RMUX_T1_SOUTH_B17_sel_value_O;
	wire [16:0] RMUX_T1_WEST_B17_O;
	wire RMUX_T1_WEST_B17_ready_out;
	wire RMUX_T1_WEST_B17_valid_out;
	wire [1:0] RMUX_T1_WEST_B17_out_sel;
	wire [0:0] RMUX_T1_WEST_B17_sel_value_O;
	wire [16:0] RMUX_T2_EAST_B17_O;
	wire RMUX_T2_EAST_B17_ready_out;
	wire RMUX_T2_EAST_B17_valid_out;
	wire [1:0] RMUX_T2_EAST_B17_out_sel;
	wire [0:0] RMUX_T2_EAST_B17_sel_value_O;
	wire [16:0] RMUX_T2_NORTH_B17_O;
	wire RMUX_T2_NORTH_B17_ready_out;
	wire RMUX_T2_NORTH_B17_valid_out;
	wire [1:0] RMUX_T2_NORTH_B17_out_sel;
	wire [0:0] RMUX_T2_NORTH_B17_sel_value_O;
	wire [16:0] RMUX_T2_SOUTH_B17_O;
	wire RMUX_T2_SOUTH_B17_ready_out;
	wire RMUX_T2_SOUTH_B17_valid_out;
	wire [1:0] RMUX_T2_SOUTH_B17_out_sel;
	wire [0:0] RMUX_T2_SOUTH_B17_sel_value_O;
	wire [16:0] RMUX_T2_WEST_B17_O;
	wire RMUX_T2_WEST_B17_ready_out;
	wire RMUX_T2_WEST_B17_valid_out;
	wire [1:0] RMUX_T2_WEST_B17_out_sel;
	wire [0:0] RMUX_T2_WEST_B17_sel_value_O;
	wire [16:0] RMUX_T3_EAST_B17_O;
	wire RMUX_T3_EAST_B17_ready_out;
	wire RMUX_T3_EAST_B17_valid_out;
	wire [1:0] RMUX_T3_EAST_B17_out_sel;
	wire [0:0] RMUX_T3_EAST_B17_sel_value_O;
	wire [16:0] RMUX_T3_NORTH_B17_O;
	wire RMUX_T3_NORTH_B17_ready_out;
	wire RMUX_T3_NORTH_B17_valid_out;
	wire [1:0] RMUX_T3_NORTH_B17_out_sel;
	wire [0:0] RMUX_T3_NORTH_B17_sel_value_O;
	wire [16:0] RMUX_T3_SOUTH_B17_O;
	wire RMUX_T3_SOUTH_B17_ready_out;
	wire RMUX_T3_SOUTH_B17_valid_out;
	wire [1:0] RMUX_T3_SOUTH_B17_out_sel;
	wire [0:0] RMUX_T3_SOUTH_B17_sel_value_O;
	wire [16:0] RMUX_T3_WEST_B17_O;
	wire RMUX_T3_WEST_B17_ready_out;
	wire RMUX_T3_WEST_B17_valid_out;
	wire [1:0] RMUX_T3_WEST_B17_out_sel;
	wire [0:0] RMUX_T3_WEST_B17_sel_value_O;
	wire [16:0] RMUX_T4_EAST_B17_O;
	wire RMUX_T4_EAST_B17_ready_out;
	wire RMUX_T4_EAST_B17_valid_out;
	wire [1:0] RMUX_T4_EAST_B17_out_sel;
	wire [0:0] RMUX_T4_EAST_B17_sel_value_O;
	wire [16:0] RMUX_T4_NORTH_B17_O;
	wire RMUX_T4_NORTH_B17_ready_out;
	wire RMUX_T4_NORTH_B17_valid_out;
	wire [1:0] RMUX_T4_NORTH_B17_out_sel;
	wire [0:0] RMUX_T4_NORTH_B17_sel_value_O;
	wire [16:0] RMUX_T4_SOUTH_B17_O;
	wire RMUX_T4_SOUTH_B17_ready_out;
	wire RMUX_T4_SOUTH_B17_valid_out;
	wire [1:0] RMUX_T4_SOUTH_B17_out_sel;
	wire [0:0] RMUX_T4_SOUTH_B17_sel_value_O;
	wire [16:0] RMUX_T4_WEST_B17_O;
	wire RMUX_T4_WEST_B17_ready_out;
	wire RMUX_T4_WEST_B17_valid_out;
	wire [1:0] RMUX_T4_WEST_B17_out_sel;
	wire [0:0] RMUX_T4_WEST_B17_sel_value_O;
	wire [0:0] SB_T0_EAST_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T0_EAST_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T0_EAST_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T0_EAST_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T0_EAST_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T0_NORTH_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T0_NORTH_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T0_NORTH_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T0_NORTH_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T0_NORTH_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T0_SOUTH_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T0_SOUTH_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T0_SOUTH_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T0_SOUTH_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T0_SOUTH_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T0_WEST_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T0_WEST_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T0_WEST_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T0_WEST_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T0_WEST_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T1_EAST_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T1_EAST_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T1_EAST_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T1_EAST_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T1_EAST_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T1_NORTH_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T1_NORTH_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T1_NORTH_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T1_NORTH_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T1_NORTH_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T1_SOUTH_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T1_SOUTH_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T1_SOUTH_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T1_SOUTH_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T1_SOUTH_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T1_WEST_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T1_WEST_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T1_WEST_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T1_WEST_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T1_WEST_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T2_EAST_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T2_EAST_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T2_EAST_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T2_EAST_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T2_EAST_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T2_NORTH_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T2_NORTH_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T2_NORTH_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T2_NORTH_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T2_NORTH_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T2_SOUTH_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T2_SOUTH_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T2_SOUTH_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T2_SOUTH_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T2_SOUTH_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T2_WEST_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T2_WEST_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T2_WEST_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T2_WEST_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T2_WEST_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T3_EAST_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T3_EAST_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T3_EAST_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T3_EAST_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T3_EAST_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T3_NORTH_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T3_NORTH_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T3_NORTH_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T3_NORTH_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T3_NORTH_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T3_SOUTH_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T3_SOUTH_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T3_SOUTH_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T3_SOUTH_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T3_SOUTH_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T3_WEST_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T3_WEST_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T3_WEST_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T3_WEST_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T3_WEST_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T4_EAST_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T4_EAST_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T4_EAST_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T4_EAST_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T4_EAST_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T4_NORTH_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T4_NORTH_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T4_NORTH_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T4_NORTH_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T4_NORTH_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T4_SOUTH_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T4_SOUTH_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T4_SOUTH_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T4_SOUTH_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T4_SOUTH_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T4_WEST_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T4_WEST_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T4_WEST_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T4_WEST_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T4_WEST_SB_OUT_B17_sel_value_O;
	wire [16:0] WIRE_SB_T0_EAST_SB_IN_B17_O;
	wire WIRE_SB_T0_EAST_SB_IN_B17_ready_out;
	wire WIRE_SB_T0_EAST_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T0_NORTH_SB_IN_B17_O;
	wire WIRE_SB_T0_NORTH_SB_IN_B17_ready_out;
	wire WIRE_SB_T0_NORTH_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T0_SOUTH_SB_IN_B17_O;
	wire WIRE_SB_T0_SOUTH_SB_IN_B17_ready_out;
	wire WIRE_SB_T0_SOUTH_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T0_WEST_SB_IN_B17_O;
	wire WIRE_SB_T0_WEST_SB_IN_B17_ready_out;
	wire WIRE_SB_T0_WEST_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T1_EAST_SB_IN_B17_O;
	wire WIRE_SB_T1_EAST_SB_IN_B17_ready_out;
	wire WIRE_SB_T1_EAST_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T1_NORTH_SB_IN_B17_O;
	wire WIRE_SB_T1_NORTH_SB_IN_B17_ready_out;
	wire WIRE_SB_T1_NORTH_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T1_SOUTH_SB_IN_B17_O;
	wire WIRE_SB_T1_SOUTH_SB_IN_B17_ready_out;
	wire WIRE_SB_T1_SOUTH_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T1_WEST_SB_IN_B17_O;
	wire WIRE_SB_T1_WEST_SB_IN_B17_ready_out;
	wire WIRE_SB_T1_WEST_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T2_EAST_SB_IN_B17_O;
	wire WIRE_SB_T2_EAST_SB_IN_B17_ready_out;
	wire WIRE_SB_T2_EAST_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T2_NORTH_SB_IN_B17_O;
	wire WIRE_SB_T2_NORTH_SB_IN_B17_ready_out;
	wire WIRE_SB_T2_NORTH_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T2_SOUTH_SB_IN_B17_O;
	wire WIRE_SB_T2_SOUTH_SB_IN_B17_ready_out;
	wire WIRE_SB_T2_SOUTH_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T2_WEST_SB_IN_B17_O;
	wire WIRE_SB_T2_WEST_SB_IN_B17_ready_out;
	wire WIRE_SB_T2_WEST_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T3_EAST_SB_IN_B17_O;
	wire WIRE_SB_T3_EAST_SB_IN_B17_ready_out;
	wire WIRE_SB_T3_EAST_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T3_NORTH_SB_IN_B17_O;
	wire WIRE_SB_T3_NORTH_SB_IN_B17_ready_out;
	wire WIRE_SB_T3_NORTH_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T3_SOUTH_SB_IN_B17_O;
	wire WIRE_SB_T3_SOUTH_SB_IN_B17_ready_out;
	wire WIRE_SB_T3_SOUTH_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T3_WEST_SB_IN_B17_O;
	wire WIRE_SB_T3_WEST_SB_IN_B17_ready_out;
	wire WIRE_SB_T3_WEST_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T4_EAST_SB_IN_B17_O;
	wire WIRE_SB_T4_EAST_SB_IN_B17_ready_out;
	wire WIRE_SB_T4_EAST_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T4_NORTH_SB_IN_B17_O;
	wire WIRE_SB_T4_NORTH_SB_IN_B17_ready_out;
	wire WIRE_SB_T4_NORTH_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T4_SOUTH_SB_IN_B17_O;
	wire WIRE_SB_T4_SOUTH_SB_IN_B17_ready_out;
	wire WIRE_SB_T4_SOUTH_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T4_WEST_SB_IN_B17_O;
	wire WIRE_SB_T4_WEST_SB_IN_B17_ready_out;
	wire WIRE_SB_T4_WEST_SB_IN_B17_valid_out;
	wire ZextWrapper_23_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_23_32_inst0$self_O_in;
	wire ZextWrapper_30_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_30_32_inst0$self_O_in;
	wire ZextWrapper_31_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_31_32_inst0$self_O_in;
	wire [0:0] and1_inst0_out;
	wire [0:0] and1_inst1_out;
	wire [0:0] and1_inst10_out;
	wire [0:0] and1_inst11_out;
	wire [0:0] and1_inst12_out;
	wire [0:0] and1_inst13_out;
	wire [0:0] and1_inst14_out;
	wire [0:0] and1_inst15_out;
	wire [0:0] and1_inst16_out;
	wire [0:0] and1_inst17_out;
	wire [0:0] and1_inst18_out;
	wire [0:0] and1_inst19_out;
	wire [0:0] and1_inst2_out;
	wire [0:0] and1_inst3_out;
	wire [0:0] and1_inst4_out;
	wire [0:0] and1_inst5_out;
	wire [0:0] and1_inst6_out;
	wire [0:0] and1_inst7_out;
	wire [0:0] and1_inst8_out;
	wire [0:0] and1_inst9_out;
	wire [31:0] config_reg_0_O;
	wire [31:0] config_reg_1_O;
	wire [31:0] config_reg_2_O;
	wire [30:0] config_reg_3_O;
	wire [29:0] config_reg_4_O;
	wire [22:0] config_reg_5_O;
	wire [0:0] const_1_1_out;
	wire coreir_eq_1_inst0_out;
	wire coreir_eq_1_inst1_out;
	wire coreir_eq_1_inst10_out;
	wire coreir_eq_1_inst11_out;
	wire coreir_eq_1_inst12_out;
	wire coreir_eq_1_inst13_out;
	wire coreir_eq_1_inst14_out;
	wire coreir_eq_1_inst15_out;
	wire coreir_eq_1_inst16_out;
	wire coreir_eq_1_inst17_out;
	wire coreir_eq_1_inst18_out;
	wire coreir_eq_1_inst19_out;
	wire coreir_eq_1_inst2_out;
	wire coreir_eq_1_inst3_out;
	wire coreir_eq_1_inst4_out;
	wire coreir_eq_1_inst5_out;
	wire coreir_eq_1_inst6_out;
	wire coreir_eq_1_inst7_out;
	wire coreir_eq_1_inst8_out;
	wire coreir_eq_1_inst9_out;
	wire [31:0] mux_aoi_6_32_inst0_O;
	wire [7:0] mux_aoi_6_32_inst0_out_sel;
	wire [7:0] self_config_config_addr_out;
	FanoutHash_330DF95D65589621 CB_PE_output_width_17_num_0_fan_in(
		.I13(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
		.E8(SB_T2_NORTH_SB_OUT_B17_enable_value_O),
		.E17(SB_T4_SOUTH_SB_OUT_B17_enable_value_O),
		.I15(MUX_SB_T3_WEST_SB_OUT_B17_ready_out),
		.I12(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out),
		.E6(SB_T1_EAST_SB_OUT_B17_enable_value_O),
		.I9(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
		.I16(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
		.E3(SB_T0_WEST_SB_OUT_B17_enable_value_O),
		.S14(MUX_SB_T3_EAST_SB_OUT_B17_out_sel),
		.E10(SB_T2_EAST_SB_OUT_B17_enable_value_O),
		.I20(PondTop_input_width_17_num_0_ready),
		.I5(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
		.S6(MUX_SB_T1_EAST_SB_OUT_B17_out_sel),
		.E0(SB_T0_NORTH_SB_OUT_B17_enable_value_O),
		.E18(SB_T4_EAST_SB_OUT_B17_enable_value_O),
		.I19(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
		.I10(MUX_SB_T2_EAST_SB_OUT_B17_ready_out),
		.S5(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel),
		.I6(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
		.I8(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
		.S3(MUX_SB_T0_WEST_SB_OUT_B17_out_sel),
		.S10(MUX_SB_T2_EAST_SB_OUT_B17_out_sel),
		.E16(SB_T4_NORTH_SB_OUT_B17_enable_value_O),
		.S4(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel),
		.E11(SB_T2_WEST_SB_OUT_B17_enable_value_O),
		.S19(MUX_SB_T4_WEST_SB_OUT_B17_out_sel),
		.E15(SB_T3_WEST_SB_OUT_B17_enable_value_O),
		.E19(SB_T4_WEST_SB_OUT_B17_enable_value_O),
		.I3(MUX_SB_T0_WEST_SB_OUT_B17_ready_out),
		.I4(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out),
		.S1(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel),
		.S21(PondTop_input_width_17_num_1_out_sel),
		.E13(SB_T3_SOUTH_SB_OUT_B17_enable_value_O),
		.S0(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T0_EAST_SB_OUT_B17_out_sel),
		.I11(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
		.S8(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel),
		.E2(SB_T0_EAST_SB_OUT_B17_enable_value_O),
		.E14(SB_T3_EAST_SB_OUT_B17_enable_value_O),
		.S17(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel),
		.E5(SB_T1_SOUTH_SB_OUT_B17_enable_value_O),
		.E4(SB_T1_NORTH_SB_OUT_B17_enable_value_O),
		.E21(PondTop_input_width_17_num_1_enable),
		.I1(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
		.I2(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
		.I17(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
		.O(CB_PE_output_width_17_num_0_fan_in_O),
		.E9(SB_T2_SOUTH_SB_OUT_B17_enable_value_O),
		.S13(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel),
		.I21(PondTop_input_width_17_num_1_ready),
		.S11(MUX_SB_T2_WEST_SB_OUT_B17_out_sel),
		.S20(PondTop_input_width_17_num_0_out_sel),
		.E1(SB_T0_SOUTH_SB_OUT_B17_enable_value_O),
		.E20(PondTop_input_width_17_num_0_enable),
		.S15(MUX_SB_T3_WEST_SB_OUT_B17_out_sel),
		.S7(MUX_SB_T1_WEST_SB_OUT_B17_out_sel),
		.S9(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel),
		.S18(MUX_SB_T4_EAST_SB_OUT_B17_out_sel),
		.S12(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel),
		.I14(MUX_SB_T3_EAST_SB_OUT_B17_ready_out),
		.I7(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
		.S16(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel),
		.E12(SB_T3_NORTH_SB_OUT_B17_enable_value_O),
		.I0(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out),
		.E7(SB_T1_WEST_SB_OUT_B17_enable_value_O),
		.I18(MUX_SB_T4_EAST_SB_OUT_B17_ready_out)
	);
	FanoutHash_82899D6851EDC11 CB_PE_output_width_17_num_1_fan_in(
		.I13(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
		.E8(SB_T2_NORTH_SB_OUT_B17_enable_value_O),
		.E17(SB_T4_SOUTH_SB_OUT_B17_enable_value_O),
		.I15(MUX_SB_T3_WEST_SB_OUT_B17_ready_out),
		.I12(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out),
		.E6(SB_T1_EAST_SB_OUT_B17_enable_value_O),
		.I9(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
		.I16(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
		.E3(SB_T0_WEST_SB_OUT_B17_enable_value_O),
		.S14(MUX_SB_T3_EAST_SB_OUT_B17_out_sel),
		.E10(SB_T2_EAST_SB_OUT_B17_enable_value_O),
		.I5(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
		.S6(MUX_SB_T1_EAST_SB_OUT_B17_out_sel),
		.E0(SB_T0_NORTH_SB_OUT_B17_enable_value_O),
		.E18(SB_T4_EAST_SB_OUT_B17_enable_value_O),
		.I19(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
		.I10(MUX_SB_T2_EAST_SB_OUT_B17_ready_out),
		.S5(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel),
		.I6(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
		.I8(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
		.S3(MUX_SB_T0_WEST_SB_OUT_B17_out_sel),
		.S10(MUX_SB_T2_EAST_SB_OUT_B17_out_sel),
		.E16(SB_T4_NORTH_SB_OUT_B17_enable_value_O),
		.S4(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel),
		.E11(SB_T2_WEST_SB_OUT_B17_enable_value_O),
		.S19(MUX_SB_T4_WEST_SB_OUT_B17_out_sel),
		.E15(SB_T3_WEST_SB_OUT_B17_enable_value_O),
		.E19(SB_T4_WEST_SB_OUT_B17_enable_value_O),
		.I3(MUX_SB_T0_WEST_SB_OUT_B17_ready_out),
		.I4(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out),
		.S1(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel),
		.E13(SB_T3_SOUTH_SB_OUT_B17_enable_value_O),
		.S0(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T0_EAST_SB_OUT_B17_out_sel),
		.I11(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
		.S8(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel),
		.E2(SB_T0_EAST_SB_OUT_B17_enable_value_O),
		.E14(SB_T3_EAST_SB_OUT_B17_enable_value_O),
		.S17(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel),
		.E5(SB_T1_SOUTH_SB_OUT_B17_enable_value_O),
		.E4(SB_T1_NORTH_SB_OUT_B17_enable_value_O),
		.I1(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
		.I2(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
		.I17(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
		.O(CB_PE_output_width_17_num_1_fan_in_O),
		.E9(SB_T2_SOUTH_SB_OUT_B17_enable_value_O),
		.S13(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel),
		.S11(MUX_SB_T2_WEST_SB_OUT_B17_out_sel),
		.S7(MUX_SB_T1_WEST_SB_OUT_B17_out_sel),
		.E1(SB_T0_SOUTH_SB_OUT_B17_enable_value_O),
		.S15(MUX_SB_T3_WEST_SB_OUT_B17_out_sel),
		.S9(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel),
		.S18(MUX_SB_T4_EAST_SB_OUT_B17_out_sel),
		.S12(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel),
		.I14(MUX_SB_T3_EAST_SB_OUT_B17_ready_out),
		.I7(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
		.S16(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel),
		.E12(SB_T3_NORTH_SB_OUT_B17_enable_value_O),
		.I0(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out),
		.E7(SB_T1_WEST_SB_OUT_B17_enable_value_O),
		.I18(MUX_SB_T4_EAST_SB_OUT_B17_ready_out)
	);
	FanoutHash_CE1AA874B742213 CB_PE_output_width_17_num_2_fan_in(
		.I13(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
		.E8(SB_T2_NORTH_SB_OUT_B17_enable_value_O),
		.E17(SB_T4_SOUTH_SB_OUT_B17_enable_value_O),
		.I15(MUX_SB_T3_WEST_SB_OUT_B17_ready_out),
		.I12(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out),
		.E6(SB_T1_EAST_SB_OUT_B17_enable_value_O),
		.I9(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
		.I16(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
		.E3(SB_T0_WEST_SB_OUT_B17_enable_value_O),
		.S14(MUX_SB_T3_EAST_SB_OUT_B17_out_sel),
		.E10(SB_T2_EAST_SB_OUT_B17_enable_value_O),
		.I5(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
		.S6(MUX_SB_T1_EAST_SB_OUT_B17_out_sel),
		.E0(SB_T0_NORTH_SB_OUT_B17_enable_value_O),
		.E18(SB_T4_EAST_SB_OUT_B17_enable_value_O),
		.I19(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
		.I10(MUX_SB_T2_EAST_SB_OUT_B17_ready_out),
		.S5(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel),
		.I6(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
		.I8(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
		.S3(MUX_SB_T0_WEST_SB_OUT_B17_out_sel),
		.S10(MUX_SB_T2_EAST_SB_OUT_B17_out_sel),
		.E16(SB_T4_NORTH_SB_OUT_B17_enable_value_O),
		.S4(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel),
		.E11(SB_T2_WEST_SB_OUT_B17_enable_value_O),
		.S19(MUX_SB_T4_WEST_SB_OUT_B17_out_sel),
		.E15(SB_T3_WEST_SB_OUT_B17_enable_value_O),
		.E19(SB_T4_WEST_SB_OUT_B17_enable_value_O),
		.I3(MUX_SB_T0_WEST_SB_OUT_B17_ready_out),
		.I4(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out),
		.S1(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel),
		.E13(SB_T3_SOUTH_SB_OUT_B17_enable_value_O),
		.S0(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T0_EAST_SB_OUT_B17_out_sel),
		.I11(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
		.S8(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel),
		.E2(SB_T0_EAST_SB_OUT_B17_enable_value_O),
		.E14(SB_T3_EAST_SB_OUT_B17_enable_value_O),
		.S17(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel),
		.E5(SB_T1_SOUTH_SB_OUT_B17_enable_value_O),
		.E4(SB_T1_NORTH_SB_OUT_B17_enable_value_O),
		.I1(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
		.I2(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
		.I17(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
		.O(CB_PE_output_width_17_num_2_fan_in_O),
		.E9(SB_T2_SOUTH_SB_OUT_B17_enable_value_O),
		.S13(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel),
		.S11(MUX_SB_T2_WEST_SB_OUT_B17_out_sel),
		.S7(MUX_SB_T1_WEST_SB_OUT_B17_out_sel),
		.E1(SB_T0_SOUTH_SB_OUT_B17_enable_value_O),
		.S15(MUX_SB_T3_WEST_SB_OUT_B17_out_sel),
		.S9(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel),
		.S18(MUX_SB_T4_EAST_SB_OUT_B17_out_sel),
		.S12(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel),
		.I14(MUX_SB_T3_EAST_SB_OUT_B17_ready_out),
		.I7(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
		.S16(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel),
		.E12(SB_T3_NORTH_SB_OUT_B17_enable_value_O),
		.I0(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out),
		.E7(SB_T1_WEST_SB_OUT_B17_enable_value_O),
		.I18(MUX_SB_T4_EAST_SB_OUT_B17_ready_out)
	);
	FanoutHash_14EBE1E8E49CA541 CB_PondTop_output_width_17_num_0_fan_in(
		.E0(PE_input_width_17_num_0_enable),
		.S0(PE_input_width_17_num_0_out_sel),
		.E1(PE_input_width_17_num_1_enable),
		.S2(PE_input_width_17_num_2_out_sel),
		.I2(PE_input_width_17_num_2_ready),
		.E2(PE_input_width_17_num_2_enable),
		.S1(PE_input_width_17_num_1_out_sel),
		.I1(PE_input_width_17_num_1_ready),
		.I0(PE_input_width_17_num_0_ready),
		.O(CB_PondTop_output_width_17_num_0_fan_in_O)
	);
	FanoutHash_1EBD0270673B29D7 CB_PondTop_output_width_17_num_1_fan_in(
		.I13(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
		.E8(SB_T2_NORTH_SB_OUT_B17_enable_value_O),
		.E17(SB_T4_SOUTH_SB_OUT_B17_enable_value_O),
		.I15(MUX_SB_T3_WEST_SB_OUT_B17_ready_out),
		.I12(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out),
		.E6(SB_T1_EAST_SB_OUT_B17_enable_value_O),
		.I9(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
		.I16(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
		.E3(SB_T0_WEST_SB_OUT_B17_enable_value_O),
		.S14(MUX_SB_T3_EAST_SB_OUT_B17_out_sel),
		.E10(SB_T2_EAST_SB_OUT_B17_enable_value_O),
		.I5(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
		.S6(MUX_SB_T1_EAST_SB_OUT_B17_out_sel),
		.E0(SB_T0_NORTH_SB_OUT_B17_enable_value_O),
		.E18(SB_T4_EAST_SB_OUT_B17_enable_value_O),
		.I19(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
		.I10(MUX_SB_T2_EAST_SB_OUT_B17_ready_out),
		.S5(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel),
		.I6(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
		.I8(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
		.S3(MUX_SB_T0_WEST_SB_OUT_B17_out_sel),
		.S10(MUX_SB_T2_EAST_SB_OUT_B17_out_sel),
		.E16(SB_T4_NORTH_SB_OUT_B17_enable_value_O),
		.S4(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel),
		.E11(SB_T2_WEST_SB_OUT_B17_enable_value_O),
		.S19(MUX_SB_T4_WEST_SB_OUT_B17_out_sel),
		.E15(SB_T3_WEST_SB_OUT_B17_enable_value_O),
		.E19(SB_T4_WEST_SB_OUT_B17_enable_value_O),
		.I3(MUX_SB_T0_WEST_SB_OUT_B17_ready_out),
		.I4(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out),
		.S1(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel),
		.E13(SB_T3_SOUTH_SB_OUT_B17_enable_value_O),
		.S0(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T0_EAST_SB_OUT_B17_out_sel),
		.I11(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
		.S8(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel),
		.E2(SB_T0_EAST_SB_OUT_B17_enable_value_O),
		.E14(SB_T3_EAST_SB_OUT_B17_enable_value_O),
		.S17(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel),
		.E5(SB_T1_SOUTH_SB_OUT_B17_enable_value_O),
		.E4(SB_T1_NORTH_SB_OUT_B17_enable_value_O),
		.I1(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
		.I2(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
		.I17(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
		.O(CB_PondTop_output_width_17_num_1_fan_in_O),
		.E9(SB_T2_SOUTH_SB_OUT_B17_enable_value_O),
		.S13(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel),
		.S11(MUX_SB_T2_WEST_SB_OUT_B17_out_sel),
		.S7(MUX_SB_T1_WEST_SB_OUT_B17_out_sel),
		.E1(SB_T0_SOUTH_SB_OUT_B17_enable_value_O),
		.S15(MUX_SB_T3_WEST_SB_OUT_B17_out_sel),
		.S9(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel),
		.S18(MUX_SB_T4_EAST_SB_OUT_B17_out_sel),
		.S12(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel),
		.I14(MUX_SB_T3_EAST_SB_OUT_B17_ready_out),
		.I7(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
		.S16(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel),
		.E12(SB_T3_NORTH_SB_OUT_B17_enable_value_O),
		.I0(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out),
		.E7(SB_T1_WEST_SB_OUT_B17_enable_value_O),
		.I18(MUX_SB_T4_EAST_SB_OUT_B17_ready_out)
	);
	coreir_not #(.width(1)) Invert1_inst0(
		.in(stall),
		.out(Invert1_inst0_out)
	);
	wire [118:0] MUX_SB_T0_EAST_SB_OUT_B17_I;
	assign MUX_SB_T0_EAST_SB_OUT_B17_I[102+:17] = PondTop_output_width_17_num_1;
	assign MUX_SB_T0_EAST_SB_OUT_B17_I[85+:17] = PE_output_width_17_num_2;
	assign MUX_SB_T0_EAST_SB_OUT_B17_I[68+:17] = PE_output_width_17_num_1;
	assign MUX_SB_T0_EAST_SB_OUT_B17_I[51+:17] = PE_output_width_17_num_0;
	assign MUX_SB_T0_EAST_SB_OUT_B17_I[34+:17] = WIRE_SB_T4_NORTH_SB_IN_B17_O;
	assign MUX_SB_T0_EAST_SB_OUT_B17_I[17+:17] = WIRE_SB_T3_SOUTH_SB_IN_B17_O;
	assign MUX_SB_T0_EAST_SB_OUT_B17_I[0+:17] = WIRE_SB_T0_WEST_SB_IN_B17_O;
	wire [6:0] MUX_SB_T0_EAST_SB_OUT_B17_valid_in;
	assign MUX_SB_T0_EAST_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid, PE_output_width_17_num_2_valid, PE_output_width_17_num_1_valid, PE_output_width_17_num_0_valid, WIRE_SB_T4_NORTH_SB_IN_B17_valid_out, WIRE_SB_T3_SOUTH_SB_IN_B17_valid_out, WIRE_SB_T0_WEST_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_7_17 MUX_SB_T0_EAST_SB_OUT_B17(
		.I(MUX_SB_T0_EAST_SB_OUT_B17_I),
		.O(MUX_SB_T0_EAST_SB_OUT_B17_O),
		.ready_in(SB_T0_EAST_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T0_EAST_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T0_EAST_SB_OUT_B17_valid_out),
		.S(SB_T0_EAST_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T0_EAST_SB_OUT_B17_out_sel)
	);
	wire [118:0] MUX_SB_T0_NORTH_SB_OUT_B17_I;
	assign MUX_SB_T0_NORTH_SB_OUT_B17_I[102+:17] = PondTop_output_width_17_num_1;
	assign MUX_SB_T0_NORTH_SB_OUT_B17_I[85+:17] = PE_output_width_17_num_2;
	assign MUX_SB_T0_NORTH_SB_OUT_B17_I[68+:17] = PE_output_width_17_num_1;
	assign MUX_SB_T0_NORTH_SB_OUT_B17_I[51+:17] = PE_output_width_17_num_0;
	assign MUX_SB_T0_NORTH_SB_OUT_B17_I[34+:17] = WIRE_SB_T0_SOUTH_SB_IN_B17_O;
	assign MUX_SB_T0_NORTH_SB_OUT_B17_I[17+:17] = WIRE_SB_T1_EAST_SB_IN_B17_O;
	assign MUX_SB_T0_NORTH_SB_OUT_B17_I[0+:17] = WIRE_SB_T0_WEST_SB_IN_B17_O;
	wire [6:0] MUX_SB_T0_NORTH_SB_OUT_B17_valid_in;
	assign MUX_SB_T0_NORTH_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid, PE_output_width_17_num_2_valid, PE_output_width_17_num_1_valid, PE_output_width_17_num_0_valid, WIRE_SB_T0_SOUTH_SB_IN_B17_valid_out, WIRE_SB_T1_EAST_SB_IN_B17_valid_out, WIRE_SB_T0_WEST_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_7_17 MUX_SB_T0_NORTH_SB_OUT_B17(
		.I(MUX_SB_T0_NORTH_SB_OUT_B17_I),
		.O(MUX_SB_T0_NORTH_SB_OUT_B17_O),
		.ready_in(SB_T0_NORTH_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T0_NORTH_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T0_NORTH_SB_OUT_B17_valid_out),
		.S(SB_T0_NORTH_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel)
	);
	wire [118:0] MUX_SB_T0_SOUTH_SB_OUT_B17_I;
	assign MUX_SB_T0_SOUTH_SB_OUT_B17_I[102+:17] = PondTop_output_width_17_num_1;
	assign MUX_SB_T0_SOUTH_SB_OUT_B17_I[85+:17] = PE_output_width_17_num_2;
	assign MUX_SB_T0_SOUTH_SB_OUT_B17_I[68+:17] = PE_output_width_17_num_1;
	assign MUX_SB_T0_SOUTH_SB_OUT_B17_I[51+:17] = PE_output_width_17_num_0;
	assign MUX_SB_T0_SOUTH_SB_OUT_B17_I[34+:17] = WIRE_SB_T1_WEST_SB_IN_B17_O;
	assign MUX_SB_T0_SOUTH_SB_OUT_B17_I[17+:17] = WIRE_SB_T0_NORTH_SB_IN_B17_O;
	assign MUX_SB_T0_SOUTH_SB_OUT_B17_I[0+:17] = WIRE_SB_T3_EAST_SB_IN_B17_O;
	wire [6:0] MUX_SB_T0_SOUTH_SB_OUT_B17_valid_in;
	assign MUX_SB_T0_SOUTH_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid, PE_output_width_17_num_2_valid, PE_output_width_17_num_1_valid, PE_output_width_17_num_0_valid, WIRE_SB_T1_WEST_SB_IN_B17_valid_out, WIRE_SB_T0_NORTH_SB_IN_B17_valid_out, WIRE_SB_T3_EAST_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_7_17 MUX_SB_T0_SOUTH_SB_OUT_B17(
		.I(MUX_SB_T0_SOUTH_SB_OUT_B17_I),
		.O(MUX_SB_T0_SOUTH_SB_OUT_B17_O),
		.ready_in(SB_T0_SOUTH_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T0_SOUTH_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T0_SOUTH_SB_OUT_B17_valid_out),
		.S(SB_T0_SOUTH_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel)
	);
	wire [118:0] MUX_SB_T0_WEST_SB_OUT_B17_I;
	assign MUX_SB_T0_WEST_SB_OUT_B17_I[102+:17] = PondTop_output_width_17_num_1;
	assign MUX_SB_T0_WEST_SB_OUT_B17_I[85+:17] = PE_output_width_17_num_2;
	assign MUX_SB_T0_WEST_SB_OUT_B17_I[68+:17] = PE_output_width_17_num_1;
	assign MUX_SB_T0_WEST_SB_OUT_B17_I[51+:17] = PE_output_width_17_num_0;
	assign MUX_SB_T0_WEST_SB_OUT_B17_I[34+:17] = WIRE_SB_T0_EAST_SB_IN_B17_O;
	assign MUX_SB_T0_WEST_SB_OUT_B17_I[17+:17] = WIRE_SB_T4_SOUTH_SB_IN_B17_O;
	assign MUX_SB_T0_WEST_SB_OUT_B17_I[0+:17] = WIRE_SB_T0_NORTH_SB_IN_B17_O;
	wire [6:0] MUX_SB_T0_WEST_SB_OUT_B17_valid_in;
	assign MUX_SB_T0_WEST_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid, PE_output_width_17_num_2_valid, PE_output_width_17_num_1_valid, PE_output_width_17_num_0_valid, WIRE_SB_T0_EAST_SB_IN_B17_valid_out, WIRE_SB_T4_SOUTH_SB_IN_B17_valid_out, WIRE_SB_T0_NORTH_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_7_17 MUX_SB_T0_WEST_SB_OUT_B17(
		.I(MUX_SB_T0_WEST_SB_OUT_B17_I),
		.O(MUX_SB_T0_WEST_SB_OUT_B17_O),
		.ready_in(SB_T0_WEST_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T0_WEST_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T0_WEST_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T0_WEST_SB_OUT_B17_valid_out),
		.S(SB_T0_WEST_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T0_WEST_SB_OUT_B17_out_sel)
	);
	wire [118:0] MUX_SB_T1_EAST_SB_OUT_B17_I;
	assign MUX_SB_T1_EAST_SB_OUT_B17_I[102+:17] = PondTop_output_width_17_num_1;
	assign MUX_SB_T1_EAST_SB_OUT_B17_I[85+:17] = PE_output_width_17_num_2;
	assign MUX_SB_T1_EAST_SB_OUT_B17_I[68+:17] = PE_output_width_17_num_1;
	assign MUX_SB_T1_EAST_SB_OUT_B17_I[51+:17] = PE_output_width_17_num_0;
	assign MUX_SB_T1_EAST_SB_OUT_B17_I[34+:17] = WIRE_SB_T2_SOUTH_SB_IN_B17_O;
	assign MUX_SB_T1_EAST_SB_OUT_B17_I[17+:17] = WIRE_SB_T1_WEST_SB_IN_B17_O;
	assign MUX_SB_T1_EAST_SB_OUT_B17_I[0+:17] = WIRE_SB_T0_NORTH_SB_IN_B17_O;
	wire [6:0] MUX_SB_T1_EAST_SB_OUT_B17_valid_in;
	assign MUX_SB_T1_EAST_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid, PE_output_width_17_num_2_valid, PE_output_width_17_num_1_valid, PE_output_width_17_num_0_valid, WIRE_SB_T2_SOUTH_SB_IN_B17_valid_out, WIRE_SB_T1_WEST_SB_IN_B17_valid_out, WIRE_SB_T0_NORTH_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_7_17 MUX_SB_T1_EAST_SB_OUT_B17(
		.I(MUX_SB_T1_EAST_SB_OUT_B17_I),
		.O(MUX_SB_T1_EAST_SB_OUT_B17_O),
		.ready_in(SB_T1_EAST_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T1_EAST_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T1_EAST_SB_OUT_B17_valid_out),
		.S(SB_T1_EAST_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T1_EAST_SB_OUT_B17_out_sel)
	);
	wire [118:0] MUX_SB_T1_NORTH_SB_OUT_B17_I;
	assign MUX_SB_T1_NORTH_SB_OUT_B17_I[102+:17] = PondTop_output_width_17_num_1;
	assign MUX_SB_T1_NORTH_SB_OUT_B17_I[85+:17] = PE_output_width_17_num_2;
	assign MUX_SB_T1_NORTH_SB_OUT_B17_I[68+:17] = PE_output_width_17_num_1;
	assign MUX_SB_T1_NORTH_SB_OUT_B17_I[51+:17] = PE_output_width_17_num_0;
	assign MUX_SB_T1_NORTH_SB_OUT_B17_I[34+:17] = WIRE_SB_T4_WEST_SB_IN_B17_O;
	assign MUX_SB_T1_NORTH_SB_OUT_B17_I[17+:17] = WIRE_SB_T1_SOUTH_SB_IN_B17_O;
	assign MUX_SB_T1_NORTH_SB_OUT_B17_I[0+:17] = WIRE_SB_T2_EAST_SB_IN_B17_O;
	wire [6:0] MUX_SB_T1_NORTH_SB_OUT_B17_valid_in;
	assign MUX_SB_T1_NORTH_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid, PE_output_width_17_num_2_valid, PE_output_width_17_num_1_valid, PE_output_width_17_num_0_valid, WIRE_SB_T4_WEST_SB_IN_B17_valid_out, WIRE_SB_T1_SOUTH_SB_IN_B17_valid_out, WIRE_SB_T2_EAST_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_7_17 MUX_SB_T1_NORTH_SB_OUT_B17(
		.I(MUX_SB_T1_NORTH_SB_OUT_B17_I),
		.O(MUX_SB_T1_NORTH_SB_OUT_B17_O),
		.ready_in(SB_T1_NORTH_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T1_NORTH_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T1_NORTH_SB_OUT_B17_valid_out),
		.S(SB_T1_NORTH_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel)
	);
	wire [118:0] MUX_SB_T1_SOUTH_SB_OUT_B17_I;
	assign MUX_SB_T1_SOUTH_SB_OUT_B17_I[102+:17] = PondTop_output_width_17_num_1;
	assign MUX_SB_T1_SOUTH_SB_OUT_B17_I[85+:17] = PE_output_width_17_num_2;
	assign MUX_SB_T1_SOUTH_SB_OUT_B17_I[68+:17] = PE_output_width_17_num_1;
	assign MUX_SB_T1_SOUTH_SB_OUT_B17_I[51+:17] = PE_output_width_17_num_0;
	assign MUX_SB_T1_SOUTH_SB_OUT_B17_I[34+:17] = WIRE_SB_T2_WEST_SB_IN_B17_O;
	assign MUX_SB_T1_SOUTH_SB_OUT_B17_I[17+:17] = WIRE_SB_T1_NORTH_SB_IN_B17_O;
	assign MUX_SB_T1_SOUTH_SB_OUT_B17_I[0+:17] = WIRE_SB_T2_EAST_SB_IN_B17_O;
	wire [6:0] MUX_SB_T1_SOUTH_SB_OUT_B17_valid_in;
	assign MUX_SB_T1_SOUTH_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid, PE_output_width_17_num_2_valid, PE_output_width_17_num_1_valid, PE_output_width_17_num_0_valid, WIRE_SB_T2_WEST_SB_IN_B17_valid_out, WIRE_SB_T1_NORTH_SB_IN_B17_valid_out, WIRE_SB_T2_EAST_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_7_17 MUX_SB_T1_SOUTH_SB_OUT_B17(
		.I(MUX_SB_T1_SOUTH_SB_OUT_B17_I),
		.O(MUX_SB_T1_SOUTH_SB_OUT_B17_O),
		.ready_in(SB_T1_SOUTH_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T1_SOUTH_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T1_SOUTH_SB_OUT_B17_valid_out),
		.S(SB_T1_SOUTH_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel)
	);
	wire [118:0] MUX_SB_T1_WEST_SB_OUT_B17_I;
	assign MUX_SB_T1_WEST_SB_OUT_B17_I[102+:17] = PondTop_output_width_17_num_1;
	assign MUX_SB_T1_WEST_SB_OUT_B17_I[85+:17] = PE_output_width_17_num_2;
	assign MUX_SB_T1_WEST_SB_OUT_B17_I[68+:17] = PE_output_width_17_num_1;
	assign MUX_SB_T1_WEST_SB_OUT_B17_I[51+:17] = PE_output_width_17_num_0;
	assign MUX_SB_T1_WEST_SB_OUT_B17_I[34+:17] = WIRE_SB_T1_EAST_SB_IN_B17_O;
	assign MUX_SB_T1_WEST_SB_OUT_B17_I[17+:17] = WIRE_SB_T0_SOUTH_SB_IN_B17_O;
	assign MUX_SB_T1_WEST_SB_OUT_B17_I[0+:17] = WIRE_SB_T4_NORTH_SB_IN_B17_O;
	wire [6:0] MUX_SB_T1_WEST_SB_OUT_B17_valid_in;
	assign MUX_SB_T1_WEST_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid, PE_output_width_17_num_2_valid, PE_output_width_17_num_1_valid, PE_output_width_17_num_0_valid, WIRE_SB_T1_EAST_SB_IN_B17_valid_out, WIRE_SB_T0_SOUTH_SB_IN_B17_valid_out, WIRE_SB_T4_NORTH_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_7_17 MUX_SB_T1_WEST_SB_OUT_B17(
		.I(MUX_SB_T1_WEST_SB_OUT_B17_I),
		.O(MUX_SB_T1_WEST_SB_OUT_B17_O),
		.ready_in(SB_T1_WEST_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T1_WEST_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T1_WEST_SB_OUT_B17_valid_out),
		.S(SB_T1_WEST_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T1_WEST_SB_OUT_B17_out_sel)
	);
	wire [118:0] MUX_SB_T2_EAST_SB_OUT_B17_I;
	assign MUX_SB_T2_EAST_SB_OUT_B17_I[102+:17] = PondTop_output_width_17_num_1;
	assign MUX_SB_T2_EAST_SB_OUT_B17_I[85+:17] = PE_output_width_17_num_2;
	assign MUX_SB_T2_EAST_SB_OUT_B17_I[68+:17] = PE_output_width_17_num_1;
	assign MUX_SB_T2_EAST_SB_OUT_B17_I[51+:17] = PE_output_width_17_num_0;
	assign MUX_SB_T2_EAST_SB_OUT_B17_I[34+:17] = WIRE_SB_T2_WEST_SB_IN_B17_O;
	assign MUX_SB_T2_EAST_SB_OUT_B17_I[17+:17] = WIRE_SB_T1_SOUTH_SB_IN_B17_O;
	assign MUX_SB_T2_EAST_SB_OUT_B17_I[0+:17] = WIRE_SB_T1_NORTH_SB_IN_B17_O;
	wire [6:0] MUX_SB_T2_EAST_SB_OUT_B17_valid_in;
	assign MUX_SB_T2_EAST_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid, PE_output_width_17_num_2_valid, PE_output_width_17_num_1_valid, PE_output_width_17_num_0_valid, WIRE_SB_T2_WEST_SB_IN_B17_valid_out, WIRE_SB_T1_SOUTH_SB_IN_B17_valid_out, WIRE_SB_T1_NORTH_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_7_17 MUX_SB_T2_EAST_SB_OUT_B17(
		.I(MUX_SB_T2_EAST_SB_OUT_B17_I),
		.O(MUX_SB_T2_EAST_SB_OUT_B17_O),
		.ready_in(SB_T2_EAST_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T2_EAST_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T2_EAST_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T2_EAST_SB_OUT_B17_valid_out),
		.S(SB_T2_EAST_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T2_EAST_SB_OUT_B17_out_sel)
	);
	wire [118:0] MUX_SB_T2_NORTH_SB_OUT_B17_I;
	assign MUX_SB_T2_NORTH_SB_OUT_B17_I[102+:17] = PondTop_output_width_17_num_1;
	assign MUX_SB_T2_NORTH_SB_OUT_B17_I[85+:17] = PE_output_width_17_num_2;
	assign MUX_SB_T2_NORTH_SB_OUT_B17_I[68+:17] = PE_output_width_17_num_1;
	assign MUX_SB_T2_NORTH_SB_OUT_B17_I[51+:17] = PE_output_width_17_num_0;
	assign MUX_SB_T2_NORTH_SB_OUT_B17_I[34+:17] = WIRE_SB_T3_WEST_SB_IN_B17_O;
	assign MUX_SB_T2_NORTH_SB_OUT_B17_I[17+:17] = WIRE_SB_T2_SOUTH_SB_IN_B17_O;
	assign MUX_SB_T2_NORTH_SB_OUT_B17_I[0+:17] = WIRE_SB_T3_EAST_SB_IN_B17_O;
	wire [6:0] MUX_SB_T2_NORTH_SB_OUT_B17_valid_in;
	assign MUX_SB_T2_NORTH_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid, PE_output_width_17_num_2_valid, PE_output_width_17_num_1_valid, PE_output_width_17_num_0_valid, WIRE_SB_T3_WEST_SB_IN_B17_valid_out, WIRE_SB_T2_SOUTH_SB_IN_B17_valid_out, WIRE_SB_T3_EAST_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_7_17 MUX_SB_T2_NORTH_SB_OUT_B17(
		.I(MUX_SB_T2_NORTH_SB_OUT_B17_I),
		.O(MUX_SB_T2_NORTH_SB_OUT_B17_O),
		.ready_in(SB_T2_NORTH_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T2_NORTH_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T2_NORTH_SB_OUT_B17_valid_out),
		.S(SB_T2_NORTH_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel)
	);
	wire [118:0] MUX_SB_T2_SOUTH_SB_OUT_B17_I;
	assign MUX_SB_T2_SOUTH_SB_OUT_B17_I[102+:17] = PondTop_output_width_17_num_1;
	assign MUX_SB_T2_SOUTH_SB_OUT_B17_I[85+:17] = PE_output_width_17_num_2;
	assign MUX_SB_T2_SOUTH_SB_OUT_B17_I[68+:17] = PE_output_width_17_num_1;
	assign MUX_SB_T2_SOUTH_SB_OUT_B17_I[51+:17] = PE_output_width_17_num_0;
	assign MUX_SB_T2_SOUTH_SB_OUT_B17_I[34+:17] = WIRE_SB_T3_WEST_SB_IN_B17_O;
	assign MUX_SB_T2_SOUTH_SB_OUT_B17_I[17+:17] = WIRE_SB_T2_NORTH_SB_IN_B17_O;
	assign MUX_SB_T2_SOUTH_SB_OUT_B17_I[0+:17] = WIRE_SB_T1_EAST_SB_IN_B17_O;
	wire [6:0] MUX_SB_T2_SOUTH_SB_OUT_B17_valid_in;
	assign MUX_SB_T2_SOUTH_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid, PE_output_width_17_num_2_valid, PE_output_width_17_num_1_valid, PE_output_width_17_num_0_valid, WIRE_SB_T3_WEST_SB_IN_B17_valid_out, WIRE_SB_T2_NORTH_SB_IN_B17_valid_out, WIRE_SB_T1_EAST_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_7_17 MUX_SB_T2_SOUTH_SB_OUT_B17(
		.I(MUX_SB_T2_SOUTH_SB_OUT_B17_I),
		.O(MUX_SB_T2_SOUTH_SB_OUT_B17_O),
		.ready_in(SB_T2_SOUTH_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T2_SOUTH_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T2_SOUTH_SB_OUT_B17_valid_out),
		.S(SB_T2_SOUTH_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel)
	);
	wire [118:0] MUX_SB_T2_WEST_SB_OUT_B17_I;
	assign MUX_SB_T2_WEST_SB_OUT_B17_I[102+:17] = PondTop_output_width_17_num_1;
	assign MUX_SB_T2_WEST_SB_OUT_B17_I[85+:17] = PE_output_width_17_num_2;
	assign MUX_SB_T2_WEST_SB_OUT_B17_I[68+:17] = PE_output_width_17_num_1;
	assign MUX_SB_T2_WEST_SB_OUT_B17_I[51+:17] = PE_output_width_17_num_0;
	assign MUX_SB_T2_WEST_SB_OUT_B17_I[34+:17] = WIRE_SB_T2_EAST_SB_IN_B17_O;
	assign MUX_SB_T2_WEST_SB_OUT_B17_I[17+:17] = WIRE_SB_T1_SOUTH_SB_IN_B17_O;
	assign MUX_SB_T2_WEST_SB_OUT_B17_I[0+:17] = WIRE_SB_T3_NORTH_SB_IN_B17_O;
	wire [6:0] MUX_SB_T2_WEST_SB_OUT_B17_valid_in;
	assign MUX_SB_T2_WEST_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid, PE_output_width_17_num_2_valid, PE_output_width_17_num_1_valid, PE_output_width_17_num_0_valid, WIRE_SB_T2_EAST_SB_IN_B17_valid_out, WIRE_SB_T1_SOUTH_SB_IN_B17_valid_out, WIRE_SB_T3_NORTH_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_7_17 MUX_SB_T2_WEST_SB_OUT_B17(
		.I(MUX_SB_T2_WEST_SB_OUT_B17_I),
		.O(MUX_SB_T2_WEST_SB_OUT_B17_O),
		.ready_in(SB_T2_WEST_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T2_WEST_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T2_WEST_SB_OUT_B17_valid_out),
		.S(SB_T2_WEST_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T2_WEST_SB_OUT_B17_out_sel)
	);
	wire [118:0] MUX_SB_T3_EAST_SB_OUT_B17_I;
	assign MUX_SB_T3_EAST_SB_OUT_B17_I[102+:17] = PondTop_output_width_17_num_1;
	assign MUX_SB_T3_EAST_SB_OUT_B17_I[85+:17] = PE_output_width_17_num_2;
	assign MUX_SB_T3_EAST_SB_OUT_B17_I[68+:17] = PE_output_width_17_num_1;
	assign MUX_SB_T3_EAST_SB_OUT_B17_I[51+:17] = PE_output_width_17_num_0;
	assign MUX_SB_T3_EAST_SB_OUT_B17_I[34+:17] = WIRE_SB_T3_WEST_SB_IN_B17_O;
	assign MUX_SB_T3_EAST_SB_OUT_B17_I[17+:17] = WIRE_SB_T2_NORTH_SB_IN_B17_O;
	assign MUX_SB_T3_EAST_SB_OUT_B17_I[0+:17] = WIRE_SB_T0_SOUTH_SB_IN_B17_O;
	wire [6:0] MUX_SB_T3_EAST_SB_OUT_B17_valid_in;
	assign MUX_SB_T3_EAST_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid, PE_output_width_17_num_2_valid, PE_output_width_17_num_1_valid, PE_output_width_17_num_0_valid, WIRE_SB_T3_WEST_SB_IN_B17_valid_out, WIRE_SB_T2_NORTH_SB_IN_B17_valid_out, WIRE_SB_T0_SOUTH_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_7_17 MUX_SB_T3_EAST_SB_OUT_B17(
		.I(MUX_SB_T3_EAST_SB_OUT_B17_I),
		.O(MUX_SB_T3_EAST_SB_OUT_B17_O),
		.ready_in(SB_T3_EAST_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T3_EAST_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T3_EAST_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T3_EAST_SB_OUT_B17_valid_out),
		.S(SB_T3_EAST_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T3_EAST_SB_OUT_B17_out_sel)
	);
	wire [118:0] MUX_SB_T3_NORTH_SB_OUT_B17_I;
	assign MUX_SB_T3_NORTH_SB_OUT_B17_I[102+:17] = PondTop_output_width_17_num_1;
	assign MUX_SB_T3_NORTH_SB_OUT_B17_I[85+:17] = PE_output_width_17_num_2;
	assign MUX_SB_T3_NORTH_SB_OUT_B17_I[68+:17] = PE_output_width_17_num_1;
	assign MUX_SB_T3_NORTH_SB_OUT_B17_I[51+:17] = PE_output_width_17_num_0;
	assign MUX_SB_T3_NORTH_SB_OUT_B17_I[34+:17] = WIRE_SB_T3_SOUTH_SB_IN_B17_O;
	assign MUX_SB_T3_NORTH_SB_OUT_B17_I[17+:17] = WIRE_SB_T4_EAST_SB_IN_B17_O;
	assign MUX_SB_T3_NORTH_SB_OUT_B17_I[0+:17] = WIRE_SB_T2_WEST_SB_IN_B17_O;
	wire [6:0] MUX_SB_T3_NORTH_SB_OUT_B17_valid_in;
	assign MUX_SB_T3_NORTH_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid, PE_output_width_17_num_2_valid, PE_output_width_17_num_1_valid, PE_output_width_17_num_0_valid, WIRE_SB_T3_SOUTH_SB_IN_B17_valid_out, WIRE_SB_T4_EAST_SB_IN_B17_valid_out, WIRE_SB_T2_WEST_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_7_17 MUX_SB_T3_NORTH_SB_OUT_B17(
		.I(MUX_SB_T3_NORTH_SB_OUT_B17_I),
		.O(MUX_SB_T3_NORTH_SB_OUT_B17_O),
		.ready_in(SB_T3_NORTH_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T3_NORTH_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T3_NORTH_SB_OUT_B17_valid_out),
		.S(SB_T3_NORTH_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel)
	);
	wire [118:0] MUX_SB_T3_SOUTH_SB_OUT_B17_I;
	assign MUX_SB_T3_SOUTH_SB_OUT_B17_I[102+:17] = PondTop_output_width_17_num_1;
	assign MUX_SB_T3_SOUTH_SB_OUT_B17_I[85+:17] = PE_output_width_17_num_2;
	assign MUX_SB_T3_SOUTH_SB_OUT_B17_I[68+:17] = PE_output_width_17_num_1;
	assign MUX_SB_T3_SOUTH_SB_OUT_B17_I[51+:17] = PE_output_width_17_num_0;
	assign MUX_SB_T3_SOUTH_SB_OUT_B17_I[34+:17] = WIRE_SB_T4_WEST_SB_IN_B17_O;
	assign MUX_SB_T3_SOUTH_SB_OUT_B17_I[17+:17] = WIRE_SB_T3_NORTH_SB_IN_B17_O;
	assign MUX_SB_T3_SOUTH_SB_OUT_B17_I[0+:17] = WIRE_SB_T0_EAST_SB_IN_B17_O;
	wire [6:0] MUX_SB_T3_SOUTH_SB_OUT_B17_valid_in;
	assign MUX_SB_T3_SOUTH_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid, PE_output_width_17_num_2_valid, PE_output_width_17_num_1_valid, PE_output_width_17_num_0_valid, WIRE_SB_T4_WEST_SB_IN_B17_valid_out, WIRE_SB_T3_NORTH_SB_IN_B17_valid_out, WIRE_SB_T0_EAST_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_7_17 MUX_SB_T3_SOUTH_SB_OUT_B17(
		.I(MUX_SB_T3_SOUTH_SB_OUT_B17_I),
		.O(MUX_SB_T3_SOUTH_SB_OUT_B17_O),
		.ready_in(SB_T3_SOUTH_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T3_SOUTH_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T3_SOUTH_SB_OUT_B17_valid_out),
		.S(SB_T3_SOUTH_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel)
	);
	wire [118:0] MUX_SB_T3_WEST_SB_OUT_B17_I;
	assign MUX_SB_T3_WEST_SB_OUT_B17_I[102+:17] = PondTop_output_width_17_num_1;
	assign MUX_SB_T3_WEST_SB_OUT_B17_I[85+:17] = PE_output_width_17_num_2;
	assign MUX_SB_T3_WEST_SB_OUT_B17_I[68+:17] = PE_output_width_17_num_1;
	assign MUX_SB_T3_WEST_SB_OUT_B17_I[51+:17] = PE_output_width_17_num_0;
	assign MUX_SB_T3_WEST_SB_OUT_B17_I[34+:17] = WIRE_SB_T3_EAST_SB_IN_B17_O;
	assign MUX_SB_T3_WEST_SB_OUT_B17_I[17+:17] = WIRE_SB_T2_SOUTH_SB_IN_B17_O;
	assign MUX_SB_T3_WEST_SB_OUT_B17_I[0+:17] = WIRE_SB_T2_NORTH_SB_IN_B17_O;
	wire [6:0] MUX_SB_T3_WEST_SB_OUT_B17_valid_in;
	assign MUX_SB_T3_WEST_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid, PE_output_width_17_num_2_valid, PE_output_width_17_num_1_valid, PE_output_width_17_num_0_valid, WIRE_SB_T3_EAST_SB_IN_B17_valid_out, WIRE_SB_T2_SOUTH_SB_IN_B17_valid_out, WIRE_SB_T2_NORTH_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_7_17 MUX_SB_T3_WEST_SB_OUT_B17(
		.I(MUX_SB_T3_WEST_SB_OUT_B17_I),
		.O(MUX_SB_T3_WEST_SB_OUT_B17_O),
		.ready_in(SB_T3_WEST_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T3_WEST_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T3_WEST_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T3_WEST_SB_OUT_B17_valid_out),
		.S(SB_T3_WEST_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T3_WEST_SB_OUT_B17_out_sel)
	);
	wire [118:0] MUX_SB_T4_EAST_SB_OUT_B17_I;
	assign MUX_SB_T4_EAST_SB_OUT_B17_I[102+:17] = PondTop_output_width_17_num_1;
	assign MUX_SB_T4_EAST_SB_OUT_B17_I[85+:17] = PE_output_width_17_num_2;
	assign MUX_SB_T4_EAST_SB_OUT_B17_I[68+:17] = PE_output_width_17_num_1;
	assign MUX_SB_T4_EAST_SB_OUT_B17_I[51+:17] = PE_output_width_17_num_0;
	assign MUX_SB_T4_EAST_SB_OUT_B17_I[34+:17] = WIRE_SB_T4_WEST_SB_IN_B17_O;
	assign MUX_SB_T4_EAST_SB_OUT_B17_I[17+:17] = WIRE_SB_T4_SOUTH_SB_IN_B17_O;
	assign MUX_SB_T4_EAST_SB_OUT_B17_I[0+:17] = WIRE_SB_T3_NORTH_SB_IN_B17_O;
	wire [6:0] MUX_SB_T4_EAST_SB_OUT_B17_valid_in;
	assign MUX_SB_T4_EAST_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid, PE_output_width_17_num_2_valid, PE_output_width_17_num_1_valid, PE_output_width_17_num_0_valid, WIRE_SB_T4_WEST_SB_IN_B17_valid_out, WIRE_SB_T4_SOUTH_SB_IN_B17_valid_out, WIRE_SB_T3_NORTH_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_7_17 MUX_SB_T4_EAST_SB_OUT_B17(
		.I(MUX_SB_T4_EAST_SB_OUT_B17_I),
		.O(MUX_SB_T4_EAST_SB_OUT_B17_O),
		.ready_in(SB_T4_EAST_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T4_EAST_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T4_EAST_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T4_EAST_SB_OUT_B17_valid_out),
		.S(SB_T4_EAST_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T4_EAST_SB_OUT_B17_out_sel)
	);
	wire [118:0] MUX_SB_T4_NORTH_SB_OUT_B17_I;
	assign MUX_SB_T4_NORTH_SB_OUT_B17_I[102+:17] = PondTop_output_width_17_num_1;
	assign MUX_SB_T4_NORTH_SB_OUT_B17_I[85+:17] = PE_output_width_17_num_2;
	assign MUX_SB_T4_NORTH_SB_OUT_B17_I[68+:17] = PE_output_width_17_num_1;
	assign MUX_SB_T4_NORTH_SB_OUT_B17_I[51+:17] = PE_output_width_17_num_0;
	assign MUX_SB_T4_NORTH_SB_OUT_B17_I[34+:17] = WIRE_SB_T4_SOUTH_SB_IN_B17_O;
	assign MUX_SB_T4_NORTH_SB_OUT_B17_I[17+:17] = WIRE_SB_T0_EAST_SB_IN_B17_O;
	assign MUX_SB_T4_NORTH_SB_OUT_B17_I[0+:17] = WIRE_SB_T1_WEST_SB_IN_B17_O;
	wire [6:0] MUX_SB_T4_NORTH_SB_OUT_B17_valid_in;
	assign MUX_SB_T4_NORTH_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid, PE_output_width_17_num_2_valid, PE_output_width_17_num_1_valid, PE_output_width_17_num_0_valid, WIRE_SB_T4_SOUTH_SB_IN_B17_valid_out, WIRE_SB_T0_EAST_SB_IN_B17_valid_out, WIRE_SB_T1_WEST_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_7_17 MUX_SB_T4_NORTH_SB_OUT_B17(
		.I(MUX_SB_T4_NORTH_SB_OUT_B17_I),
		.O(MUX_SB_T4_NORTH_SB_OUT_B17_O),
		.ready_in(SB_T4_NORTH_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T4_NORTH_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T4_NORTH_SB_OUT_B17_valid_out),
		.S(SB_T4_NORTH_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel)
	);
	wire [118:0] MUX_SB_T4_SOUTH_SB_OUT_B17_I;
	assign MUX_SB_T4_SOUTH_SB_OUT_B17_I[102+:17] = PondTop_output_width_17_num_1;
	assign MUX_SB_T4_SOUTH_SB_OUT_B17_I[85+:17] = PE_output_width_17_num_2;
	assign MUX_SB_T4_SOUTH_SB_OUT_B17_I[68+:17] = PE_output_width_17_num_1;
	assign MUX_SB_T4_SOUTH_SB_OUT_B17_I[51+:17] = PE_output_width_17_num_0;
	assign MUX_SB_T4_SOUTH_SB_OUT_B17_I[34+:17] = WIRE_SB_T4_NORTH_SB_IN_B17_O;
	assign MUX_SB_T4_SOUTH_SB_OUT_B17_I[17+:17] = WIRE_SB_T4_EAST_SB_IN_B17_O;
	assign MUX_SB_T4_SOUTH_SB_OUT_B17_I[0+:17] = WIRE_SB_T0_WEST_SB_IN_B17_O;
	wire [6:0] MUX_SB_T4_SOUTH_SB_OUT_B17_valid_in;
	assign MUX_SB_T4_SOUTH_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid, PE_output_width_17_num_2_valid, PE_output_width_17_num_1_valid, PE_output_width_17_num_0_valid, WIRE_SB_T4_NORTH_SB_IN_B17_valid_out, WIRE_SB_T4_EAST_SB_IN_B17_valid_out, WIRE_SB_T0_WEST_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_7_17 MUX_SB_T4_SOUTH_SB_OUT_B17(
		.I(MUX_SB_T4_SOUTH_SB_OUT_B17_I),
		.O(MUX_SB_T4_SOUTH_SB_OUT_B17_O),
		.ready_in(SB_T4_SOUTH_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T4_SOUTH_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T4_SOUTH_SB_OUT_B17_valid_out),
		.S(SB_T4_SOUTH_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel)
	);
	wire [118:0] MUX_SB_T4_WEST_SB_OUT_B17_I;
	assign MUX_SB_T4_WEST_SB_OUT_B17_I[102+:17] = PondTop_output_width_17_num_1;
	assign MUX_SB_T4_WEST_SB_OUT_B17_I[85+:17] = PE_output_width_17_num_2;
	assign MUX_SB_T4_WEST_SB_OUT_B17_I[68+:17] = PE_output_width_17_num_1;
	assign MUX_SB_T4_WEST_SB_OUT_B17_I[51+:17] = PE_output_width_17_num_0;
	assign MUX_SB_T4_WEST_SB_OUT_B17_I[34+:17] = WIRE_SB_T4_EAST_SB_IN_B17_O;
	assign MUX_SB_T4_WEST_SB_OUT_B17_I[17+:17] = WIRE_SB_T3_SOUTH_SB_IN_B17_O;
	assign MUX_SB_T4_WEST_SB_OUT_B17_I[0+:17] = WIRE_SB_T1_NORTH_SB_IN_B17_O;
	wire [6:0] MUX_SB_T4_WEST_SB_OUT_B17_valid_in;
	assign MUX_SB_T4_WEST_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid, PE_output_width_17_num_2_valid, PE_output_width_17_num_1_valid, PE_output_width_17_num_0_valid, WIRE_SB_T4_EAST_SB_IN_B17_valid_out, WIRE_SB_T3_SOUTH_SB_IN_B17_valid_out, WIRE_SB_T1_NORTH_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_7_17 MUX_SB_T4_WEST_SB_OUT_B17(
		.I(MUX_SB_T4_WEST_SB_OUT_B17_I),
		.O(MUX_SB_T4_WEST_SB_OUT_B17_O),
		.ready_in(SB_T4_WEST_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T4_WEST_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T4_WEST_SB_OUT_B17_valid_out),
		.S(SB_T4_WEST_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T4_WEST_SB_OUT_B17_out_sel)
	);
	SplitFifo_17 REG_T0_EAST_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T0_EAST_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T0_EAST_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T0_EAST_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T0_EAST_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst2_out[0]),
		.end_fifo(REG_T0_EAST_B17_end_value_O[0]),
		.valid0(MUX_SB_T0_EAST_SB_OUT_B17_valid_out),
		.valid1(REG_T0_EAST_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T0_EAST_B17_ready_out),
		.fifo_en(REG_T0_EAST_B17_fifo_value_O[0])
	);
	SliceWrapper_32_0_1 REG_T0_EAST_B17_end_value(
		.I(config_reg_0_O),
		.O(REG_T0_EAST_B17_end_value_O)
	);
	SliceWrapper_32_1_2 REG_T0_EAST_B17_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T0_EAST_B17_fifo_value_O)
	);
	SliceWrapper_32_2_3 REG_T0_EAST_B17_start_value(
		.I(config_reg_0_O),
		.O(REG_T0_EAST_B17_start_value_O)
	);
	SplitFifo_17 REG_T0_NORTH_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T0_NORTH_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T0_NORTH_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T0_NORTH_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T0_NORTH_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst0_out[0]),
		.end_fifo(REG_T0_NORTH_B17_end_value_O[0]),
		.valid0(MUX_SB_T0_NORTH_SB_OUT_B17_valid_out),
		.valid1(REG_T0_NORTH_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T0_NORTH_B17_ready_out),
		.fifo_en(REG_T0_NORTH_B17_fifo_value_O[0])
	);
	SliceWrapper_32_3_4 REG_T0_NORTH_B17_end_value(
		.I(config_reg_0_O),
		.O(REG_T0_NORTH_B17_end_value_O)
	);
	SliceWrapper_32_4_5 REG_T0_NORTH_B17_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T0_NORTH_B17_fifo_value_O)
	);
	SliceWrapper_32_5_6 REG_T0_NORTH_B17_start_value(
		.I(config_reg_0_O),
		.O(REG_T0_NORTH_B17_start_value_O)
	);
	SplitFifo_17 REG_T0_SOUTH_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T0_SOUTH_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T0_SOUTH_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T0_SOUTH_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T0_SOUTH_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst1_out[0]),
		.end_fifo(REG_T0_SOUTH_B17_end_value_O[0]),
		.valid0(MUX_SB_T0_SOUTH_SB_OUT_B17_valid_out),
		.valid1(REG_T0_SOUTH_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T0_SOUTH_B17_ready_out),
		.fifo_en(REG_T0_SOUTH_B17_fifo_value_O[0])
	);
	SliceWrapper_32_6_7 REG_T0_SOUTH_B17_end_value(
		.I(config_reg_0_O),
		.O(REG_T0_SOUTH_B17_end_value_O)
	);
	SliceWrapper_32_7_8 REG_T0_SOUTH_B17_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T0_SOUTH_B17_fifo_value_O)
	);
	SliceWrapper_32_8_9 REG_T0_SOUTH_B17_start_value(
		.I(config_reg_0_O),
		.O(REG_T0_SOUTH_B17_start_value_O)
	);
	SplitFifo_17 REG_T0_WEST_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T0_WEST_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T0_WEST_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T0_WEST_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T0_WEST_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst3_out[0]),
		.end_fifo(REG_T0_WEST_B17_end_value_O[0]),
		.valid0(MUX_SB_T0_WEST_SB_OUT_B17_valid_out),
		.valid1(REG_T0_WEST_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T0_WEST_B17_ready_out),
		.fifo_en(REG_T0_WEST_B17_fifo_value_O[0])
	);
	SliceWrapper_32_9_10 REG_T0_WEST_B17_end_value(
		.I(config_reg_0_O),
		.O(REG_T0_WEST_B17_end_value_O)
	);
	SliceWrapper_32_10_11 REG_T0_WEST_B17_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T0_WEST_B17_fifo_value_O)
	);
	SliceWrapper_32_11_12 REG_T0_WEST_B17_start_value(
		.I(config_reg_0_O),
		.O(REG_T0_WEST_B17_start_value_O)
	);
	SplitFifo_17 REG_T1_EAST_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T1_EAST_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T1_EAST_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T1_EAST_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T1_EAST_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst6_out[0]),
		.end_fifo(REG_T1_EAST_B17_end_value_O[0]),
		.valid0(MUX_SB_T1_EAST_SB_OUT_B17_valid_out),
		.valid1(REG_T1_EAST_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T1_EAST_B17_ready_out),
		.fifo_en(REG_T1_EAST_B17_fifo_value_O[0])
	);
	SliceWrapper_32_12_13 REG_T1_EAST_B17_end_value(
		.I(config_reg_0_O),
		.O(REG_T1_EAST_B17_end_value_O)
	);
	SliceWrapper_32_13_14 REG_T1_EAST_B17_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T1_EAST_B17_fifo_value_O)
	);
	SliceWrapper_32_14_15 REG_T1_EAST_B17_start_value(
		.I(config_reg_0_O),
		.O(REG_T1_EAST_B17_start_value_O)
	);
	SplitFifo_17 REG_T1_NORTH_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T1_NORTH_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T1_NORTH_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T1_NORTH_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T1_NORTH_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst4_out[0]),
		.end_fifo(REG_T1_NORTH_B17_end_value_O[0]),
		.valid0(MUX_SB_T1_NORTH_SB_OUT_B17_valid_out),
		.valid1(REG_T1_NORTH_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T1_NORTH_B17_ready_out),
		.fifo_en(REG_T1_NORTH_B17_fifo_value_O[0])
	);
	SliceWrapper_32_15_16 REG_T1_NORTH_B17_end_value(
		.I(config_reg_0_O),
		.O(REG_T1_NORTH_B17_end_value_O)
	);
	SliceWrapper_32_16_17 REG_T1_NORTH_B17_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T1_NORTH_B17_fifo_value_O)
	);
	SliceWrapper_32_17_18 REG_T1_NORTH_B17_start_value(
		.I(config_reg_0_O),
		.O(REG_T1_NORTH_B17_start_value_O)
	);
	SplitFifo_17 REG_T1_SOUTH_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T1_SOUTH_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T1_SOUTH_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T1_SOUTH_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T1_SOUTH_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst5_out[0]),
		.end_fifo(REG_T1_SOUTH_B17_end_value_O[0]),
		.valid0(MUX_SB_T1_SOUTH_SB_OUT_B17_valid_out),
		.valid1(REG_T1_SOUTH_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T1_SOUTH_B17_ready_out),
		.fifo_en(REG_T1_SOUTH_B17_fifo_value_O[0])
	);
	SliceWrapper_32_18_19 REG_T1_SOUTH_B17_end_value(
		.I(config_reg_0_O),
		.O(REG_T1_SOUTH_B17_end_value_O)
	);
	SliceWrapper_32_19_20 REG_T1_SOUTH_B17_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T1_SOUTH_B17_fifo_value_O)
	);
	SliceWrapper_32_20_21 REG_T1_SOUTH_B17_start_value(
		.I(config_reg_0_O),
		.O(REG_T1_SOUTH_B17_start_value_O)
	);
	SplitFifo_17 REG_T1_WEST_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T1_WEST_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T1_WEST_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T1_WEST_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T1_WEST_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst7_out[0]),
		.end_fifo(REG_T1_WEST_B17_end_value_O[0]),
		.valid0(MUX_SB_T1_WEST_SB_OUT_B17_valid_out),
		.valid1(REG_T1_WEST_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T1_WEST_B17_ready_out),
		.fifo_en(REG_T1_WEST_B17_fifo_value_O[0])
	);
	SliceWrapper_32_21_22 REG_T1_WEST_B17_end_value(
		.I(config_reg_0_O),
		.O(REG_T1_WEST_B17_end_value_O)
	);
	SliceWrapper_32_22_23 REG_T1_WEST_B17_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T1_WEST_B17_fifo_value_O)
	);
	SliceWrapper_32_23_24 REG_T1_WEST_B17_start_value(
		.I(config_reg_0_O),
		.O(REG_T1_WEST_B17_start_value_O)
	);
	SplitFifo_17 REG_T2_EAST_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T2_EAST_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T2_EAST_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T2_EAST_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T2_EAST_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst10_out[0]),
		.end_fifo(REG_T2_EAST_B17_end_value_O[0]),
		.valid0(MUX_SB_T2_EAST_SB_OUT_B17_valid_out),
		.valid1(REG_T2_EAST_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T2_EAST_B17_ready_out),
		.fifo_en(REG_T2_EAST_B17_fifo_value_O[0])
	);
	SliceWrapper_32_24_25 REG_T2_EAST_B17_end_value(
		.I(config_reg_0_O),
		.O(REG_T2_EAST_B17_end_value_O)
	);
	SliceWrapper_32_25_26 REG_T2_EAST_B17_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T2_EAST_B17_fifo_value_O)
	);
	SliceWrapper_32_26_27 REG_T2_EAST_B17_start_value(
		.I(config_reg_0_O),
		.O(REG_T2_EAST_B17_start_value_O)
	);
	SplitFifo_17 REG_T2_NORTH_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T2_NORTH_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T2_NORTH_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T2_NORTH_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T2_NORTH_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst8_out[0]),
		.end_fifo(REG_T2_NORTH_B17_end_value_O[0]),
		.valid0(MUX_SB_T2_NORTH_SB_OUT_B17_valid_out),
		.valid1(REG_T2_NORTH_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T2_NORTH_B17_ready_out),
		.fifo_en(REG_T2_NORTH_B17_fifo_value_O[0])
	);
	SliceWrapper_32_27_28 REG_T2_NORTH_B17_end_value(
		.I(config_reg_0_O),
		.O(REG_T2_NORTH_B17_end_value_O)
	);
	SliceWrapper_32_28_29 REG_T2_NORTH_B17_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T2_NORTH_B17_fifo_value_O)
	);
	SliceWrapper_32_29_30 REG_T2_NORTH_B17_start_value(
		.I(config_reg_0_O),
		.O(REG_T2_NORTH_B17_start_value_O)
	);
	SplitFifo_17 REG_T2_SOUTH_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T2_SOUTH_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T2_SOUTH_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T2_SOUTH_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T2_SOUTH_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst9_out[0]),
		.end_fifo(REG_T2_SOUTH_B17_end_value_O[0]),
		.valid0(MUX_SB_T2_SOUTH_SB_OUT_B17_valid_out),
		.valid1(REG_T2_SOUTH_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T2_SOUTH_B17_ready_out),
		.fifo_en(REG_T2_SOUTH_B17_fifo_value_O[0])
	);
	SliceWrapper_32_30_31 REG_T2_SOUTH_B17_end_value(
		.I(config_reg_0_O),
		.O(REG_T2_SOUTH_B17_end_value_O)
	);
	SliceWrapper_32_31_32 REG_T2_SOUTH_B17_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T2_SOUTH_B17_fifo_value_O)
	);
	SliceWrapper_32_0_1 REG_T2_SOUTH_B17_start_value(
		.I(config_reg_1_O),
		.O(REG_T2_SOUTH_B17_start_value_O)
	);
	SplitFifo_17 REG_T2_WEST_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T2_WEST_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T2_WEST_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T2_WEST_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T2_WEST_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst11_out[0]),
		.end_fifo(REG_T2_WEST_B17_end_value_O[0]),
		.valid0(MUX_SB_T2_WEST_SB_OUT_B17_valid_out),
		.valid1(REG_T2_WEST_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T2_WEST_B17_ready_out),
		.fifo_en(REG_T2_WEST_B17_fifo_value_O[0])
	);
	SliceWrapper_32_1_2 REG_T2_WEST_B17_end_value(
		.I(config_reg_1_O),
		.O(REG_T2_WEST_B17_end_value_O)
	);
	SliceWrapper_32_2_3 REG_T2_WEST_B17_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T2_WEST_B17_fifo_value_O)
	);
	SliceWrapper_32_3_4 REG_T2_WEST_B17_start_value(
		.I(config_reg_1_O),
		.O(REG_T2_WEST_B17_start_value_O)
	);
	SplitFifo_17 REG_T3_EAST_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T3_EAST_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T3_EAST_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T3_EAST_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T3_EAST_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst14_out[0]),
		.end_fifo(REG_T3_EAST_B17_end_value_O[0]),
		.valid0(MUX_SB_T3_EAST_SB_OUT_B17_valid_out),
		.valid1(REG_T3_EAST_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T3_EAST_B17_ready_out),
		.fifo_en(REG_T3_EAST_B17_fifo_value_O[0])
	);
	SliceWrapper_32_4_5 REG_T3_EAST_B17_end_value(
		.I(config_reg_1_O),
		.O(REG_T3_EAST_B17_end_value_O)
	);
	SliceWrapper_32_5_6 REG_T3_EAST_B17_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T3_EAST_B17_fifo_value_O)
	);
	SliceWrapper_32_6_7 REG_T3_EAST_B17_start_value(
		.I(config_reg_1_O),
		.O(REG_T3_EAST_B17_start_value_O)
	);
	SplitFifo_17 REG_T3_NORTH_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T3_NORTH_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T3_NORTH_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T3_NORTH_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T3_NORTH_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst12_out[0]),
		.end_fifo(REG_T3_NORTH_B17_end_value_O[0]),
		.valid0(MUX_SB_T3_NORTH_SB_OUT_B17_valid_out),
		.valid1(REG_T3_NORTH_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T3_NORTH_B17_ready_out),
		.fifo_en(REG_T3_NORTH_B17_fifo_value_O[0])
	);
	SliceWrapper_32_7_8 REG_T3_NORTH_B17_end_value(
		.I(config_reg_1_O),
		.O(REG_T3_NORTH_B17_end_value_O)
	);
	SliceWrapper_32_8_9 REG_T3_NORTH_B17_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T3_NORTH_B17_fifo_value_O)
	);
	SliceWrapper_32_9_10 REG_T3_NORTH_B17_start_value(
		.I(config_reg_1_O),
		.O(REG_T3_NORTH_B17_start_value_O)
	);
	SplitFifo_17 REG_T3_SOUTH_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T3_SOUTH_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T3_SOUTH_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T3_SOUTH_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T3_SOUTH_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst13_out[0]),
		.end_fifo(REG_T3_SOUTH_B17_end_value_O[0]),
		.valid0(MUX_SB_T3_SOUTH_SB_OUT_B17_valid_out),
		.valid1(REG_T3_SOUTH_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T3_SOUTH_B17_ready_out),
		.fifo_en(REG_T3_SOUTH_B17_fifo_value_O[0])
	);
	SliceWrapper_32_10_11 REG_T3_SOUTH_B17_end_value(
		.I(config_reg_1_O),
		.O(REG_T3_SOUTH_B17_end_value_O)
	);
	SliceWrapper_32_11_12 REG_T3_SOUTH_B17_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T3_SOUTH_B17_fifo_value_O)
	);
	SliceWrapper_32_12_13 REG_T3_SOUTH_B17_start_value(
		.I(config_reg_1_O),
		.O(REG_T3_SOUTH_B17_start_value_O)
	);
	SplitFifo_17 REG_T3_WEST_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T3_WEST_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T3_WEST_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T3_WEST_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T3_WEST_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst15_out[0]),
		.end_fifo(REG_T3_WEST_B17_end_value_O[0]),
		.valid0(MUX_SB_T3_WEST_SB_OUT_B17_valid_out),
		.valid1(REG_T3_WEST_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T3_WEST_B17_ready_out),
		.fifo_en(REG_T3_WEST_B17_fifo_value_O[0])
	);
	SliceWrapper_32_13_14 REG_T3_WEST_B17_end_value(
		.I(config_reg_1_O),
		.O(REG_T3_WEST_B17_end_value_O)
	);
	SliceWrapper_32_14_15 REG_T3_WEST_B17_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T3_WEST_B17_fifo_value_O)
	);
	SliceWrapper_32_15_16 REG_T3_WEST_B17_start_value(
		.I(config_reg_1_O),
		.O(REG_T3_WEST_B17_start_value_O)
	);
	SplitFifo_17 REG_T4_EAST_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T4_EAST_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T4_EAST_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T4_EAST_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T4_EAST_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst18_out[0]),
		.end_fifo(REG_T4_EAST_B17_end_value_O[0]),
		.valid0(MUX_SB_T4_EAST_SB_OUT_B17_valid_out),
		.valid1(REG_T4_EAST_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T4_EAST_B17_ready_out),
		.fifo_en(REG_T4_EAST_B17_fifo_value_O[0])
	);
	SliceWrapper_32_16_17 REG_T4_EAST_B17_end_value(
		.I(config_reg_1_O),
		.O(REG_T4_EAST_B17_end_value_O)
	);
	SliceWrapper_32_17_18 REG_T4_EAST_B17_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T4_EAST_B17_fifo_value_O)
	);
	SliceWrapper_32_18_19 REG_T4_EAST_B17_start_value(
		.I(config_reg_1_O),
		.O(REG_T4_EAST_B17_start_value_O)
	);
	SplitFifo_17 REG_T4_NORTH_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T4_NORTH_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T4_NORTH_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T4_NORTH_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T4_NORTH_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst16_out[0]),
		.end_fifo(REG_T4_NORTH_B17_end_value_O[0]),
		.valid0(MUX_SB_T4_NORTH_SB_OUT_B17_valid_out),
		.valid1(REG_T4_NORTH_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T4_NORTH_B17_ready_out),
		.fifo_en(REG_T4_NORTH_B17_fifo_value_O[0])
	);
	SliceWrapper_32_19_20 REG_T4_NORTH_B17_end_value(
		.I(config_reg_1_O),
		.O(REG_T4_NORTH_B17_end_value_O)
	);
	SliceWrapper_32_20_21 REG_T4_NORTH_B17_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T4_NORTH_B17_fifo_value_O)
	);
	SliceWrapper_32_21_22 REG_T4_NORTH_B17_start_value(
		.I(config_reg_1_O),
		.O(REG_T4_NORTH_B17_start_value_O)
	);
	SplitFifo_17 REG_T4_SOUTH_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T4_SOUTH_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T4_SOUTH_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T4_SOUTH_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T4_SOUTH_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst17_out[0]),
		.end_fifo(REG_T4_SOUTH_B17_end_value_O[0]),
		.valid0(MUX_SB_T4_SOUTH_SB_OUT_B17_valid_out),
		.valid1(REG_T4_SOUTH_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T4_SOUTH_B17_ready_out),
		.fifo_en(REG_T4_SOUTH_B17_fifo_value_O[0])
	);
	SliceWrapper_32_22_23 REG_T4_SOUTH_B17_end_value(
		.I(config_reg_1_O),
		.O(REG_T4_SOUTH_B17_end_value_O)
	);
	SliceWrapper_32_23_24 REG_T4_SOUTH_B17_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T4_SOUTH_B17_fifo_value_O)
	);
	SliceWrapper_32_24_25 REG_T4_SOUTH_B17_start_value(
		.I(config_reg_1_O),
		.O(REG_T4_SOUTH_B17_start_value_O)
	);
	SplitFifo_17 REG_T4_WEST_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T4_WEST_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T4_WEST_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T4_WEST_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T4_WEST_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst19_out[0]),
		.end_fifo(REG_T4_WEST_B17_end_value_O[0]),
		.valid0(MUX_SB_T4_WEST_SB_OUT_B17_valid_out),
		.valid1(REG_T4_WEST_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T4_WEST_B17_ready_out),
		.fifo_en(REG_T4_WEST_B17_fifo_value_O[0])
	);
	SliceWrapper_32_25_26 REG_T4_WEST_B17_end_value(
		.I(config_reg_1_O),
		.O(REG_T4_WEST_B17_end_value_O)
	);
	SliceWrapper_32_26_27 REG_T4_WEST_B17_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T4_WEST_B17_fifo_value_O)
	);
	SliceWrapper_32_27_28 REG_T4_WEST_B17_start_value(
		.I(config_reg_1_O),
		.O(REG_T4_WEST_B17_start_value_O)
	);
	wire [33:0] RMUX_T0_EAST_B17_I;
	assign RMUX_T0_EAST_B17_I[17+:17] = REG_T0_EAST_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T0_EAST_B17_I[0+:17] = MUX_SB_T0_EAST_SB_OUT_B17_O;
	wire [1:0] RMUX_T0_EAST_B17_valid_in;
	assign RMUX_T0_EAST_B17_valid_in = {REG_T0_EAST_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T0_EAST_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T0_EAST_B17(
		.I(RMUX_T0_EAST_B17_I),
		.O(RMUX_T0_EAST_B17_O),
		.ready_in(SB_T0_EAST_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T0_EAST_B17_ready_out),
		.valid_in(RMUX_T0_EAST_B17_valid_in),
		.valid_out(RMUX_T0_EAST_B17_valid_out),
		.S(RMUX_T0_EAST_B17_sel_value_O),
		.out_sel(RMUX_T0_EAST_B17_out_sel)
	);
	SliceWrapper_32_28_29 RMUX_T0_EAST_B17_sel_value(
		.I(config_reg_1_O),
		.O(RMUX_T0_EAST_B17_sel_value_O)
	);
	wire [33:0] RMUX_T0_NORTH_B17_I;
	assign RMUX_T0_NORTH_B17_I[17+:17] = REG_T0_NORTH_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T0_NORTH_B17_I[0+:17] = MUX_SB_T0_NORTH_SB_OUT_B17_O;
	wire [1:0] RMUX_T0_NORTH_B17_valid_in;
	assign RMUX_T0_NORTH_B17_valid_in = {REG_T0_NORTH_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T0_NORTH_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T0_NORTH_B17(
		.I(RMUX_T0_NORTH_B17_I),
		.O(RMUX_T0_NORTH_B17_O),
		.ready_in(SB_T0_NORTH_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T0_NORTH_B17_ready_out),
		.valid_in(RMUX_T0_NORTH_B17_valid_in),
		.valid_out(RMUX_T0_NORTH_B17_valid_out),
		.S(RMUX_T0_NORTH_B17_sel_value_O),
		.out_sel(RMUX_T0_NORTH_B17_out_sel)
	);
	SliceWrapper_32_29_30 RMUX_T0_NORTH_B17_sel_value(
		.I(config_reg_1_O),
		.O(RMUX_T0_NORTH_B17_sel_value_O)
	);
	wire [33:0] RMUX_T0_SOUTH_B17_I;
	assign RMUX_T0_SOUTH_B17_I[17+:17] = REG_T0_SOUTH_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T0_SOUTH_B17_I[0+:17] = MUX_SB_T0_SOUTH_SB_OUT_B17_O;
	wire [1:0] RMUX_T0_SOUTH_B17_valid_in;
	assign RMUX_T0_SOUTH_B17_valid_in = {REG_T0_SOUTH_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T0_SOUTH_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T0_SOUTH_B17(
		.I(RMUX_T0_SOUTH_B17_I),
		.O(RMUX_T0_SOUTH_B17_O),
		.ready_in(SB_T0_SOUTH_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T0_SOUTH_B17_ready_out),
		.valid_in(RMUX_T0_SOUTH_B17_valid_in),
		.valid_out(RMUX_T0_SOUTH_B17_valid_out),
		.S(RMUX_T0_SOUTH_B17_sel_value_O),
		.out_sel(RMUX_T0_SOUTH_B17_out_sel)
	);
	SliceWrapper_32_30_31 RMUX_T0_SOUTH_B17_sel_value(
		.I(config_reg_1_O),
		.O(RMUX_T0_SOUTH_B17_sel_value_O)
	);
	wire [33:0] RMUX_T0_WEST_B17_I;
	assign RMUX_T0_WEST_B17_I[17+:17] = REG_T0_WEST_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T0_WEST_B17_I[0+:17] = MUX_SB_T0_WEST_SB_OUT_B17_O;
	wire [1:0] RMUX_T0_WEST_B17_valid_in;
	assign RMUX_T0_WEST_B17_valid_in = {REG_T0_WEST_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T0_WEST_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T0_WEST_B17(
		.I(RMUX_T0_WEST_B17_I),
		.O(RMUX_T0_WEST_B17_O),
		.ready_in(SB_T0_WEST_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T0_WEST_B17_ready_out),
		.valid_in(RMUX_T0_WEST_B17_valid_in),
		.valid_out(RMUX_T0_WEST_B17_valid_out),
		.S(RMUX_T0_WEST_B17_sel_value_O),
		.out_sel(RMUX_T0_WEST_B17_out_sel)
	);
	SliceWrapper_32_31_32 RMUX_T0_WEST_B17_sel_value(
		.I(config_reg_1_O),
		.O(RMUX_T0_WEST_B17_sel_value_O)
	);
	wire [33:0] RMUX_T1_EAST_B17_I;
	assign RMUX_T1_EAST_B17_I[17+:17] = REG_T1_EAST_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T1_EAST_B17_I[0+:17] = MUX_SB_T1_EAST_SB_OUT_B17_O;
	wire [1:0] RMUX_T1_EAST_B17_valid_in;
	assign RMUX_T1_EAST_B17_valid_in = {REG_T1_EAST_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T1_EAST_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T1_EAST_B17(
		.I(RMUX_T1_EAST_B17_I),
		.O(RMUX_T1_EAST_B17_O),
		.ready_in(SB_T1_EAST_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T1_EAST_B17_ready_out),
		.valid_in(RMUX_T1_EAST_B17_valid_in),
		.valid_out(RMUX_T1_EAST_B17_valid_out),
		.S(RMUX_T1_EAST_B17_sel_value_O),
		.out_sel(RMUX_T1_EAST_B17_out_sel)
	);
	SliceWrapper_32_0_1 RMUX_T1_EAST_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T1_EAST_B17_sel_value_O)
	);
	wire [33:0] RMUX_T1_NORTH_B17_I;
	assign RMUX_T1_NORTH_B17_I[17+:17] = REG_T1_NORTH_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T1_NORTH_B17_I[0+:17] = MUX_SB_T1_NORTH_SB_OUT_B17_O;
	wire [1:0] RMUX_T1_NORTH_B17_valid_in;
	assign RMUX_T1_NORTH_B17_valid_in = {REG_T1_NORTH_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T1_NORTH_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T1_NORTH_B17(
		.I(RMUX_T1_NORTH_B17_I),
		.O(RMUX_T1_NORTH_B17_O),
		.ready_in(SB_T1_NORTH_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T1_NORTH_B17_ready_out),
		.valid_in(RMUX_T1_NORTH_B17_valid_in),
		.valid_out(RMUX_T1_NORTH_B17_valid_out),
		.S(RMUX_T1_NORTH_B17_sel_value_O),
		.out_sel(RMUX_T1_NORTH_B17_out_sel)
	);
	SliceWrapper_32_1_2 RMUX_T1_NORTH_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T1_NORTH_B17_sel_value_O)
	);
	wire [33:0] RMUX_T1_SOUTH_B17_I;
	assign RMUX_T1_SOUTH_B17_I[17+:17] = REG_T1_SOUTH_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T1_SOUTH_B17_I[0+:17] = MUX_SB_T1_SOUTH_SB_OUT_B17_O;
	wire [1:0] RMUX_T1_SOUTH_B17_valid_in;
	assign RMUX_T1_SOUTH_B17_valid_in = {REG_T1_SOUTH_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T1_SOUTH_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T1_SOUTH_B17(
		.I(RMUX_T1_SOUTH_B17_I),
		.O(RMUX_T1_SOUTH_B17_O),
		.ready_in(SB_T1_SOUTH_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T1_SOUTH_B17_ready_out),
		.valid_in(RMUX_T1_SOUTH_B17_valid_in),
		.valid_out(RMUX_T1_SOUTH_B17_valid_out),
		.S(RMUX_T1_SOUTH_B17_sel_value_O),
		.out_sel(RMUX_T1_SOUTH_B17_out_sel)
	);
	SliceWrapper_32_2_3 RMUX_T1_SOUTH_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T1_SOUTH_B17_sel_value_O)
	);
	wire [33:0] RMUX_T1_WEST_B17_I;
	assign RMUX_T1_WEST_B17_I[17+:17] = REG_T1_WEST_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T1_WEST_B17_I[0+:17] = MUX_SB_T1_WEST_SB_OUT_B17_O;
	wire [1:0] RMUX_T1_WEST_B17_valid_in;
	assign RMUX_T1_WEST_B17_valid_in = {REG_T1_WEST_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T1_WEST_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T1_WEST_B17(
		.I(RMUX_T1_WEST_B17_I),
		.O(RMUX_T1_WEST_B17_O),
		.ready_in(SB_T1_WEST_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T1_WEST_B17_ready_out),
		.valid_in(RMUX_T1_WEST_B17_valid_in),
		.valid_out(RMUX_T1_WEST_B17_valid_out),
		.S(RMUX_T1_WEST_B17_sel_value_O),
		.out_sel(RMUX_T1_WEST_B17_out_sel)
	);
	SliceWrapper_32_3_4 RMUX_T1_WEST_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T1_WEST_B17_sel_value_O)
	);
	wire [33:0] RMUX_T2_EAST_B17_I;
	assign RMUX_T2_EAST_B17_I[17+:17] = REG_T2_EAST_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T2_EAST_B17_I[0+:17] = MUX_SB_T2_EAST_SB_OUT_B17_O;
	wire [1:0] RMUX_T2_EAST_B17_valid_in;
	assign RMUX_T2_EAST_B17_valid_in = {REG_T2_EAST_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T2_EAST_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T2_EAST_B17(
		.I(RMUX_T2_EAST_B17_I),
		.O(RMUX_T2_EAST_B17_O),
		.ready_in(SB_T2_EAST_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T2_EAST_B17_ready_out),
		.valid_in(RMUX_T2_EAST_B17_valid_in),
		.valid_out(RMUX_T2_EAST_B17_valid_out),
		.S(RMUX_T2_EAST_B17_sel_value_O),
		.out_sel(RMUX_T2_EAST_B17_out_sel)
	);
	SliceWrapper_32_4_5 RMUX_T2_EAST_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T2_EAST_B17_sel_value_O)
	);
	wire [33:0] RMUX_T2_NORTH_B17_I;
	assign RMUX_T2_NORTH_B17_I[17+:17] = REG_T2_NORTH_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T2_NORTH_B17_I[0+:17] = MUX_SB_T2_NORTH_SB_OUT_B17_O;
	wire [1:0] RMUX_T2_NORTH_B17_valid_in;
	assign RMUX_T2_NORTH_B17_valid_in = {REG_T2_NORTH_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T2_NORTH_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T2_NORTH_B17(
		.I(RMUX_T2_NORTH_B17_I),
		.O(RMUX_T2_NORTH_B17_O),
		.ready_in(SB_T2_NORTH_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T2_NORTH_B17_ready_out),
		.valid_in(RMUX_T2_NORTH_B17_valid_in),
		.valid_out(RMUX_T2_NORTH_B17_valid_out),
		.S(RMUX_T2_NORTH_B17_sel_value_O),
		.out_sel(RMUX_T2_NORTH_B17_out_sel)
	);
	SliceWrapper_32_5_6 RMUX_T2_NORTH_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T2_NORTH_B17_sel_value_O)
	);
	wire [33:0] RMUX_T2_SOUTH_B17_I;
	assign RMUX_T2_SOUTH_B17_I[17+:17] = REG_T2_SOUTH_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T2_SOUTH_B17_I[0+:17] = MUX_SB_T2_SOUTH_SB_OUT_B17_O;
	wire [1:0] RMUX_T2_SOUTH_B17_valid_in;
	assign RMUX_T2_SOUTH_B17_valid_in = {REG_T2_SOUTH_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T2_SOUTH_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T2_SOUTH_B17(
		.I(RMUX_T2_SOUTH_B17_I),
		.O(RMUX_T2_SOUTH_B17_O),
		.ready_in(SB_T2_SOUTH_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T2_SOUTH_B17_ready_out),
		.valid_in(RMUX_T2_SOUTH_B17_valid_in),
		.valid_out(RMUX_T2_SOUTH_B17_valid_out),
		.S(RMUX_T2_SOUTH_B17_sel_value_O),
		.out_sel(RMUX_T2_SOUTH_B17_out_sel)
	);
	SliceWrapper_32_6_7 RMUX_T2_SOUTH_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T2_SOUTH_B17_sel_value_O)
	);
	wire [33:0] RMUX_T2_WEST_B17_I;
	assign RMUX_T2_WEST_B17_I[17+:17] = REG_T2_WEST_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T2_WEST_B17_I[0+:17] = MUX_SB_T2_WEST_SB_OUT_B17_O;
	wire [1:0] RMUX_T2_WEST_B17_valid_in;
	assign RMUX_T2_WEST_B17_valid_in = {REG_T2_WEST_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T2_WEST_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T2_WEST_B17(
		.I(RMUX_T2_WEST_B17_I),
		.O(RMUX_T2_WEST_B17_O),
		.ready_in(SB_T2_WEST_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T2_WEST_B17_ready_out),
		.valid_in(RMUX_T2_WEST_B17_valid_in),
		.valid_out(RMUX_T2_WEST_B17_valid_out),
		.S(RMUX_T2_WEST_B17_sel_value_O),
		.out_sel(RMUX_T2_WEST_B17_out_sel)
	);
	SliceWrapper_32_7_8 RMUX_T2_WEST_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T2_WEST_B17_sel_value_O)
	);
	wire [33:0] RMUX_T3_EAST_B17_I;
	assign RMUX_T3_EAST_B17_I[17+:17] = REG_T3_EAST_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T3_EAST_B17_I[0+:17] = MUX_SB_T3_EAST_SB_OUT_B17_O;
	wire [1:0] RMUX_T3_EAST_B17_valid_in;
	assign RMUX_T3_EAST_B17_valid_in = {REG_T3_EAST_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T3_EAST_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T3_EAST_B17(
		.I(RMUX_T3_EAST_B17_I),
		.O(RMUX_T3_EAST_B17_O),
		.ready_in(SB_T3_EAST_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T3_EAST_B17_ready_out),
		.valid_in(RMUX_T3_EAST_B17_valid_in),
		.valid_out(RMUX_T3_EAST_B17_valid_out),
		.S(RMUX_T3_EAST_B17_sel_value_O),
		.out_sel(RMUX_T3_EAST_B17_out_sel)
	);
	SliceWrapper_32_8_9 RMUX_T3_EAST_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T3_EAST_B17_sel_value_O)
	);
	wire [33:0] RMUX_T3_NORTH_B17_I;
	assign RMUX_T3_NORTH_B17_I[17+:17] = REG_T3_NORTH_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T3_NORTH_B17_I[0+:17] = MUX_SB_T3_NORTH_SB_OUT_B17_O;
	wire [1:0] RMUX_T3_NORTH_B17_valid_in;
	assign RMUX_T3_NORTH_B17_valid_in = {REG_T3_NORTH_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T3_NORTH_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T3_NORTH_B17(
		.I(RMUX_T3_NORTH_B17_I),
		.O(RMUX_T3_NORTH_B17_O),
		.ready_in(SB_T3_NORTH_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T3_NORTH_B17_ready_out),
		.valid_in(RMUX_T3_NORTH_B17_valid_in),
		.valid_out(RMUX_T3_NORTH_B17_valid_out),
		.S(RMUX_T3_NORTH_B17_sel_value_O),
		.out_sel(RMUX_T3_NORTH_B17_out_sel)
	);
	SliceWrapper_32_9_10 RMUX_T3_NORTH_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T3_NORTH_B17_sel_value_O)
	);
	wire [33:0] RMUX_T3_SOUTH_B17_I;
	assign RMUX_T3_SOUTH_B17_I[17+:17] = REG_T3_SOUTH_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T3_SOUTH_B17_I[0+:17] = MUX_SB_T3_SOUTH_SB_OUT_B17_O;
	wire [1:0] RMUX_T3_SOUTH_B17_valid_in;
	assign RMUX_T3_SOUTH_B17_valid_in = {REG_T3_SOUTH_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T3_SOUTH_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T3_SOUTH_B17(
		.I(RMUX_T3_SOUTH_B17_I),
		.O(RMUX_T3_SOUTH_B17_O),
		.ready_in(SB_T3_SOUTH_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T3_SOUTH_B17_ready_out),
		.valid_in(RMUX_T3_SOUTH_B17_valid_in),
		.valid_out(RMUX_T3_SOUTH_B17_valid_out),
		.S(RMUX_T3_SOUTH_B17_sel_value_O),
		.out_sel(RMUX_T3_SOUTH_B17_out_sel)
	);
	SliceWrapper_32_10_11 RMUX_T3_SOUTH_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T3_SOUTH_B17_sel_value_O)
	);
	wire [33:0] RMUX_T3_WEST_B17_I;
	assign RMUX_T3_WEST_B17_I[17+:17] = REG_T3_WEST_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T3_WEST_B17_I[0+:17] = MUX_SB_T3_WEST_SB_OUT_B17_O;
	wire [1:0] RMUX_T3_WEST_B17_valid_in;
	assign RMUX_T3_WEST_B17_valid_in = {REG_T3_WEST_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T3_WEST_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T3_WEST_B17(
		.I(RMUX_T3_WEST_B17_I),
		.O(RMUX_T3_WEST_B17_O),
		.ready_in(SB_T3_WEST_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T3_WEST_B17_ready_out),
		.valid_in(RMUX_T3_WEST_B17_valid_in),
		.valid_out(RMUX_T3_WEST_B17_valid_out),
		.S(RMUX_T3_WEST_B17_sel_value_O),
		.out_sel(RMUX_T3_WEST_B17_out_sel)
	);
	SliceWrapper_32_11_12 RMUX_T3_WEST_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T3_WEST_B17_sel_value_O)
	);
	wire [33:0] RMUX_T4_EAST_B17_I;
	assign RMUX_T4_EAST_B17_I[17+:17] = REG_T4_EAST_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T4_EAST_B17_I[0+:17] = MUX_SB_T4_EAST_SB_OUT_B17_O;
	wire [1:0] RMUX_T4_EAST_B17_valid_in;
	assign RMUX_T4_EAST_B17_valid_in = {REG_T4_EAST_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T4_EAST_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T4_EAST_B17(
		.I(RMUX_T4_EAST_B17_I),
		.O(RMUX_T4_EAST_B17_O),
		.ready_in(SB_T4_EAST_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T4_EAST_B17_ready_out),
		.valid_in(RMUX_T4_EAST_B17_valid_in),
		.valid_out(RMUX_T4_EAST_B17_valid_out),
		.S(RMUX_T4_EAST_B17_sel_value_O),
		.out_sel(RMUX_T4_EAST_B17_out_sel)
	);
	SliceWrapper_32_12_13 RMUX_T4_EAST_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T4_EAST_B17_sel_value_O)
	);
	wire [33:0] RMUX_T4_NORTH_B17_I;
	assign RMUX_T4_NORTH_B17_I[17+:17] = REG_T4_NORTH_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T4_NORTH_B17_I[0+:17] = MUX_SB_T4_NORTH_SB_OUT_B17_O;
	wire [1:0] RMUX_T4_NORTH_B17_valid_in;
	assign RMUX_T4_NORTH_B17_valid_in = {REG_T4_NORTH_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T4_NORTH_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T4_NORTH_B17(
		.I(RMUX_T4_NORTH_B17_I),
		.O(RMUX_T4_NORTH_B17_O),
		.ready_in(SB_T4_NORTH_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T4_NORTH_B17_ready_out),
		.valid_in(RMUX_T4_NORTH_B17_valid_in),
		.valid_out(RMUX_T4_NORTH_B17_valid_out),
		.S(RMUX_T4_NORTH_B17_sel_value_O),
		.out_sel(RMUX_T4_NORTH_B17_out_sel)
	);
	SliceWrapper_32_13_14 RMUX_T4_NORTH_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T4_NORTH_B17_sel_value_O)
	);
	wire [33:0] RMUX_T4_SOUTH_B17_I;
	assign RMUX_T4_SOUTH_B17_I[17+:17] = REG_T4_SOUTH_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T4_SOUTH_B17_I[0+:17] = MUX_SB_T4_SOUTH_SB_OUT_B17_O;
	wire [1:0] RMUX_T4_SOUTH_B17_valid_in;
	assign RMUX_T4_SOUTH_B17_valid_in = {REG_T4_SOUTH_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T4_SOUTH_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T4_SOUTH_B17(
		.I(RMUX_T4_SOUTH_B17_I),
		.O(RMUX_T4_SOUTH_B17_O),
		.ready_in(SB_T4_SOUTH_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T4_SOUTH_B17_ready_out),
		.valid_in(RMUX_T4_SOUTH_B17_valid_in),
		.valid_out(RMUX_T4_SOUTH_B17_valid_out),
		.S(RMUX_T4_SOUTH_B17_sel_value_O),
		.out_sel(RMUX_T4_SOUTH_B17_out_sel)
	);
	SliceWrapper_32_14_15 RMUX_T4_SOUTH_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T4_SOUTH_B17_sel_value_O)
	);
	wire [33:0] RMUX_T4_WEST_B17_I;
	assign RMUX_T4_WEST_B17_I[17+:17] = REG_T4_WEST_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T4_WEST_B17_I[0+:17] = MUX_SB_T4_WEST_SB_OUT_B17_O;
	wire [1:0] RMUX_T4_WEST_B17_valid_in;
	assign RMUX_T4_WEST_B17_valid_in = {REG_T4_WEST_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T4_WEST_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T4_WEST_B17(
		.I(RMUX_T4_WEST_B17_I),
		.O(RMUX_T4_WEST_B17_O),
		.ready_in(SB_T4_WEST_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T4_WEST_B17_ready_out),
		.valid_in(RMUX_T4_WEST_B17_valid_in),
		.valid_out(RMUX_T4_WEST_B17_valid_out),
		.S(RMUX_T4_WEST_B17_sel_value_O),
		.out_sel(RMUX_T4_WEST_B17_out_sel)
	);
	SliceWrapper_32_15_16 RMUX_T4_WEST_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T4_WEST_B17_sel_value_O)
	);
	SliceWrapper_32_16_17 SB_T0_EAST_SB_IN_B17_enable_value(
		.I(config_reg_2_O),
		.O(SB_T0_EAST_SB_IN_B17_enable_value_O)
	);
	FanoutHash_55B00FA90A0098BB SB_T0_EAST_SB_IN_B17_fan_in(
		.E8(PondTop_input_width_17_num_1_enable),
		.E6(PE_input_width_17_num_3_enable),
		.E3(PE_input_width_17_num_0_enable),
		.I5(PE_input_width_17_num_2_ready),
		.S6(PE_input_width_17_num_3_out_sel),
		.E0(SB_T0_WEST_SB_OUT_B17_enable_value_O),
		.S5(PE_input_width_17_num_2_out_sel),
		.I6(PE_input_width_17_num_3_ready),
		.I8(PondTop_input_width_17_num_1_ready),
		.S3(PE_input_width_17_num_0_out_sel),
		.S4(PE_input_width_17_num_1_out_sel),
		.I3(PE_input_width_17_num_0_ready),
		.I4(PE_input_width_17_num_1_ready),
		.S1(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T0_WEST_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel),
		.S8(PondTop_input_width_17_num_1_out_sel),
		.E2(SB_T4_NORTH_SB_OUT_B17_enable_value_O),
		.E5(PE_input_width_17_num_2_enable),
		.E4(PE_input_width_17_num_1_enable),
		.I2(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
		.O(SB_T0_EAST_SB_IN_B17_fan_in_O),
		.S7(PondTop_input_width_17_num_0_out_sel),
		.E1(SB_T3_SOUTH_SB_OUT_B17_enable_value_O),
		.I7(PondTop_input_width_17_num_0_ready),
		.I0(MUX_SB_T0_WEST_SB_OUT_B17_ready_out),
		.E7(PondTop_input_width_17_num_0_enable)
	);
	wire [1:0] SB_T0_EAST_SB_OUT_B17_FANOUT_I;
	assign SB_T0_EAST_SB_OUT_B17_FANOUT_I = {REG_T0_EAST_B17$SplitFifo_17_inst0_ready0[0], RMUX_T0_EAST_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T0_EAST_SB_OUT_B17_FANOUT(
		.O(SB_T0_EAST_SB_OUT_B17_FANOUT_O),
		.I(SB_T0_EAST_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T0_EAST_B17_out_sel)
	);
	SliceWrapper_32_17_18 SB_T0_EAST_SB_OUT_B17_enable_value(
		.I(config_reg_2_O),
		.O(SB_T0_EAST_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_32_18_21 SB_T0_EAST_SB_OUT_B17_sel_value(
		.I(config_reg_2_O),
		.O(SB_T0_EAST_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_32_21_22 SB_T0_NORTH_SB_IN_B17_enable_value(
		.I(config_reg_2_O),
		.O(SB_T0_NORTH_SB_IN_B17_enable_value_O)
	);
	FanoutHash_3A6A5822E84DCC71 SB_T0_NORTH_SB_IN_B17_fan_in(
		.E8(PondTop_input_width_17_num_1_enable),
		.E6(PE_input_width_17_num_3_enable),
		.E3(PE_input_width_17_num_0_enable),
		.I5(PE_input_width_17_num_2_ready),
		.S6(PE_input_width_17_num_3_out_sel),
		.E0(SB_T0_WEST_SB_OUT_B17_enable_value_O),
		.S5(PE_input_width_17_num_2_out_sel),
		.I6(PE_input_width_17_num_3_ready),
		.I8(PondTop_input_width_17_num_1_ready),
		.S3(PE_input_width_17_num_0_out_sel),
		.S4(PE_input_width_17_num_1_out_sel),
		.I3(PE_input_width_17_num_0_ready),
		.I4(PE_input_width_17_num_1_ready),
		.S1(MUX_SB_T1_EAST_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T0_WEST_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel),
		.S8(PondTop_input_width_17_num_1_out_sel),
		.E2(SB_T0_SOUTH_SB_OUT_B17_enable_value_O),
		.E5(PE_input_width_17_num_2_enable),
		.E4(PE_input_width_17_num_1_enable),
		.I2(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
		.O(SB_T0_NORTH_SB_IN_B17_fan_in_O),
		.S7(PondTop_input_width_17_num_0_out_sel),
		.E1(SB_T1_EAST_SB_OUT_B17_enable_value_O),
		.I7(PondTop_input_width_17_num_0_ready),
		.I0(MUX_SB_T0_WEST_SB_OUT_B17_ready_out),
		.E7(PondTop_input_width_17_num_0_enable)
	);
	wire [1:0] SB_T0_NORTH_SB_OUT_B17_FANOUT_I;
	assign SB_T0_NORTH_SB_OUT_B17_FANOUT_I = {REG_T0_NORTH_B17$SplitFifo_17_inst0_ready0[0], RMUX_T0_NORTH_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T0_NORTH_SB_OUT_B17_FANOUT(
		.O(SB_T0_NORTH_SB_OUT_B17_FANOUT_O),
		.I(SB_T0_NORTH_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T0_NORTH_B17_out_sel)
	);
	SliceWrapper_32_22_23 SB_T0_NORTH_SB_OUT_B17_enable_value(
		.I(config_reg_2_O),
		.O(SB_T0_NORTH_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_32_23_26 SB_T0_NORTH_SB_OUT_B17_sel_value(
		.I(config_reg_2_O),
		.O(SB_T0_NORTH_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_32_26_27 SB_T0_SOUTH_SB_IN_B17_enable_value(
		.I(config_reg_2_O),
		.O(SB_T0_SOUTH_SB_IN_B17_enable_value_O)
	);
	FanoutHash_3E05574A9CE9CA8A SB_T0_SOUTH_SB_IN_B17_fan_in(
		.E8(PondTop_input_width_17_num_1_enable),
		.E6(PE_input_width_17_num_3_enable),
		.E3(PE_input_width_17_num_0_enable),
		.I5(PE_input_width_17_num_2_ready),
		.S6(PE_input_width_17_num_3_out_sel),
		.E0(SB_T3_EAST_SB_OUT_B17_enable_value_O),
		.S5(PE_input_width_17_num_2_out_sel),
		.I6(PE_input_width_17_num_3_ready),
		.I8(PondTop_input_width_17_num_1_ready),
		.S3(PE_input_width_17_num_0_out_sel),
		.S4(PE_input_width_17_num_1_out_sel),
		.I3(PE_input_width_17_num_0_ready),
		.I4(PE_input_width_17_num_1_ready),
		.S1(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T3_EAST_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T1_WEST_SB_OUT_B17_out_sel),
		.S8(PondTop_input_width_17_num_1_out_sel),
		.E2(SB_T1_WEST_SB_OUT_B17_enable_value_O),
		.E5(PE_input_width_17_num_2_enable),
		.E4(PE_input_width_17_num_1_enable),
		.I2(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out),
		.O(SB_T0_SOUTH_SB_IN_B17_fan_in_O),
		.S7(PondTop_input_width_17_num_0_out_sel),
		.E1(SB_T0_NORTH_SB_OUT_B17_enable_value_O),
		.I7(PondTop_input_width_17_num_0_ready),
		.I0(MUX_SB_T3_EAST_SB_OUT_B17_ready_out),
		.E7(PondTop_input_width_17_num_0_enable)
	);
	wire [1:0] SB_T0_SOUTH_SB_OUT_B17_FANOUT_I;
	assign SB_T0_SOUTH_SB_OUT_B17_FANOUT_I = {REG_T0_SOUTH_B17$SplitFifo_17_inst0_ready0[0], RMUX_T0_SOUTH_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T0_SOUTH_SB_OUT_B17_FANOUT(
		.O(SB_T0_SOUTH_SB_OUT_B17_FANOUT_O),
		.I(SB_T0_SOUTH_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T0_SOUTH_B17_out_sel)
	);
	SliceWrapper_32_27_28 SB_T0_SOUTH_SB_OUT_B17_enable_value(
		.I(config_reg_2_O),
		.O(SB_T0_SOUTH_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_32_28_31 SB_T0_SOUTH_SB_OUT_B17_sel_value(
		.I(config_reg_2_O),
		.O(SB_T0_SOUTH_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_32_31_32 SB_T0_WEST_SB_IN_B17_enable_value(
		.I(config_reg_2_O),
		.O(SB_T0_WEST_SB_IN_B17_enable_value_O)
	);
	FanoutHash_87642A353688B49 SB_T0_WEST_SB_IN_B17_fan_in(
		.E8(PondTop_input_width_17_num_1_enable),
		.E6(PE_input_width_17_num_3_enable),
		.E3(PE_input_width_17_num_0_enable),
		.I5(PE_input_width_17_num_2_ready),
		.S6(PE_input_width_17_num_3_out_sel),
		.E0(SB_T0_NORTH_SB_OUT_B17_enable_value_O),
		.S5(PE_input_width_17_num_2_out_sel),
		.I6(PE_input_width_17_num_3_ready),
		.I8(PondTop_input_width_17_num_1_ready),
		.S3(PE_input_width_17_num_0_out_sel),
		.S4(PE_input_width_17_num_1_out_sel),
		.I3(PE_input_width_17_num_0_ready),
		.I4(PE_input_width_17_num_1_ready),
		.S1(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T0_EAST_SB_OUT_B17_out_sel),
		.S8(PondTop_input_width_17_num_1_out_sel),
		.E2(SB_T0_EAST_SB_OUT_B17_enable_value_O),
		.E5(PE_input_width_17_num_2_enable),
		.E4(PE_input_width_17_num_1_enable),
		.I2(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
		.O(SB_T0_WEST_SB_IN_B17_fan_in_O),
		.S7(PondTop_input_width_17_num_0_out_sel),
		.E1(SB_T4_SOUTH_SB_OUT_B17_enable_value_O),
		.I7(PondTop_input_width_17_num_0_ready),
		.I0(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out),
		.E7(PondTop_input_width_17_num_0_enable)
	);
	wire [1:0] SB_T0_WEST_SB_OUT_B17_FANOUT_I;
	assign SB_T0_WEST_SB_OUT_B17_FANOUT_I = {REG_T0_WEST_B17$SplitFifo_17_inst0_ready0[0], RMUX_T0_WEST_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T0_WEST_SB_OUT_B17_FANOUT(
		.O(SB_T0_WEST_SB_OUT_B17_FANOUT_O),
		.I(SB_T0_WEST_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T0_WEST_B17_out_sel)
	);
	SliceWrapper_31_0_1 SB_T0_WEST_SB_OUT_B17_enable_value(
		.I(config_reg_3_O),
		.O(SB_T0_WEST_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_31_1_4 SB_T0_WEST_SB_OUT_B17_sel_value(
		.I(config_reg_3_O),
		.O(SB_T0_WEST_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_31_4_5 SB_T1_EAST_SB_IN_B17_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_EAST_SB_IN_B17_enable_value_O)
	);
	FanoutHash_245560850976C879 SB_T1_EAST_SB_IN_B17_fan_in(
		.E8(PondTop_input_width_17_num_1_enable),
		.E6(PE_input_width_17_num_3_enable),
		.E3(PE_input_width_17_num_0_enable),
		.I5(PE_input_width_17_num_2_ready),
		.S6(PE_input_width_17_num_3_out_sel),
		.E0(SB_T0_NORTH_SB_OUT_B17_enable_value_O),
		.S5(PE_input_width_17_num_2_out_sel),
		.I6(PE_input_width_17_num_3_ready),
		.I8(PondTop_input_width_17_num_1_ready),
		.S3(PE_input_width_17_num_0_out_sel),
		.S4(PE_input_width_17_num_1_out_sel),
		.I3(PE_input_width_17_num_0_ready),
		.I4(PE_input_width_17_num_1_ready),
		.S1(MUX_SB_T1_WEST_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel),
		.S8(PondTop_input_width_17_num_1_out_sel),
		.E2(SB_T2_SOUTH_SB_OUT_B17_enable_value_O),
		.E5(PE_input_width_17_num_2_enable),
		.E4(PE_input_width_17_num_1_enable),
		.I2(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
		.O(SB_T1_EAST_SB_IN_B17_fan_in_O),
		.S7(PondTop_input_width_17_num_0_out_sel),
		.E1(SB_T1_WEST_SB_OUT_B17_enable_value_O),
		.I7(PondTop_input_width_17_num_0_ready),
		.I0(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out),
		.E7(PondTop_input_width_17_num_0_enable)
	);
	wire [1:0] SB_T1_EAST_SB_OUT_B17_FANOUT_I;
	assign SB_T1_EAST_SB_OUT_B17_FANOUT_I = {REG_T1_EAST_B17$SplitFifo_17_inst0_ready0[0], RMUX_T1_EAST_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T1_EAST_SB_OUT_B17_FANOUT(
		.O(SB_T1_EAST_SB_OUT_B17_FANOUT_O),
		.I(SB_T1_EAST_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T1_EAST_B17_out_sel)
	);
	SliceWrapper_31_5_6 SB_T1_EAST_SB_OUT_B17_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_EAST_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_31_6_9 SB_T1_EAST_SB_OUT_B17_sel_value(
		.I(config_reg_3_O),
		.O(SB_T1_EAST_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_31_9_10 SB_T1_NORTH_SB_IN_B17_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_NORTH_SB_IN_B17_enable_value_O)
	);
	FanoutHash_37E9FE88073C5BAC SB_T1_NORTH_SB_IN_B17_fan_in(
		.E8(PondTop_input_width_17_num_1_enable),
		.E6(PE_input_width_17_num_3_enable),
		.E3(PE_input_width_17_num_0_enable),
		.I5(PE_input_width_17_num_2_ready),
		.S6(PE_input_width_17_num_3_out_sel),
		.E0(SB_T2_EAST_SB_OUT_B17_enable_value_O),
		.S5(PE_input_width_17_num_2_out_sel),
		.I6(PE_input_width_17_num_3_ready),
		.I8(PondTop_input_width_17_num_1_ready),
		.S3(PE_input_width_17_num_0_out_sel),
		.S4(PE_input_width_17_num_1_out_sel),
		.I3(PE_input_width_17_num_0_ready),
		.I4(PE_input_width_17_num_1_ready),
		.S1(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T2_EAST_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T4_WEST_SB_OUT_B17_out_sel),
		.S8(PondTop_input_width_17_num_1_out_sel),
		.E2(SB_T4_WEST_SB_OUT_B17_enable_value_O),
		.E5(PE_input_width_17_num_2_enable),
		.E4(PE_input_width_17_num_1_enable),
		.I2(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
		.O(SB_T1_NORTH_SB_IN_B17_fan_in_O),
		.S7(PondTop_input_width_17_num_0_out_sel),
		.E1(SB_T1_SOUTH_SB_OUT_B17_enable_value_O),
		.I7(PondTop_input_width_17_num_0_ready),
		.I0(MUX_SB_T2_EAST_SB_OUT_B17_ready_out),
		.E7(PondTop_input_width_17_num_0_enable)
	);
	wire [1:0] SB_T1_NORTH_SB_OUT_B17_FANOUT_I;
	assign SB_T1_NORTH_SB_OUT_B17_FANOUT_I = {REG_T1_NORTH_B17$SplitFifo_17_inst0_ready0[0], RMUX_T1_NORTH_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T1_NORTH_SB_OUT_B17_FANOUT(
		.O(SB_T1_NORTH_SB_OUT_B17_FANOUT_O),
		.I(SB_T1_NORTH_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T1_NORTH_B17_out_sel)
	);
	SliceWrapper_31_10_11 SB_T1_NORTH_SB_OUT_B17_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_NORTH_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_31_11_14 SB_T1_NORTH_SB_OUT_B17_sel_value(
		.I(config_reg_3_O),
		.O(SB_T1_NORTH_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_31_14_15 SB_T1_SOUTH_SB_IN_B17_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_SOUTH_SB_IN_B17_enable_value_O)
	);
	FanoutHash_2F92967E9F56D548 SB_T1_SOUTH_SB_IN_B17_fan_in(
		.E8(PondTop_input_width_17_num_1_enable),
		.E6(PE_input_width_17_num_3_enable),
		.E3(PE_input_width_17_num_0_enable),
		.I5(PE_input_width_17_num_2_ready),
		.S6(PE_input_width_17_num_3_out_sel),
		.E0(SB_T2_EAST_SB_OUT_B17_enable_value_O),
		.S5(PE_input_width_17_num_2_out_sel),
		.I6(PE_input_width_17_num_3_ready),
		.I8(PondTop_input_width_17_num_1_ready),
		.S3(PE_input_width_17_num_0_out_sel),
		.S4(PE_input_width_17_num_1_out_sel),
		.I3(PE_input_width_17_num_0_ready),
		.I4(PE_input_width_17_num_1_ready),
		.S1(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T2_EAST_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T2_WEST_SB_OUT_B17_out_sel),
		.S8(PondTop_input_width_17_num_1_out_sel),
		.E2(SB_T2_WEST_SB_OUT_B17_enable_value_O),
		.E5(PE_input_width_17_num_2_enable),
		.E4(PE_input_width_17_num_1_enable),
		.I2(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out),
		.O(SB_T1_SOUTH_SB_IN_B17_fan_in_O),
		.S7(PondTop_input_width_17_num_0_out_sel),
		.E1(SB_T1_NORTH_SB_OUT_B17_enable_value_O),
		.I7(PondTop_input_width_17_num_0_ready),
		.I0(MUX_SB_T2_EAST_SB_OUT_B17_ready_out),
		.E7(PondTop_input_width_17_num_0_enable)
	);
	wire [1:0] SB_T1_SOUTH_SB_OUT_B17_FANOUT_I;
	assign SB_T1_SOUTH_SB_OUT_B17_FANOUT_I = {REG_T1_SOUTH_B17$SplitFifo_17_inst0_ready0[0], RMUX_T1_SOUTH_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T1_SOUTH_SB_OUT_B17_FANOUT(
		.O(SB_T1_SOUTH_SB_OUT_B17_FANOUT_O),
		.I(SB_T1_SOUTH_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T1_SOUTH_B17_out_sel)
	);
	SliceWrapper_31_15_16 SB_T1_SOUTH_SB_OUT_B17_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_SOUTH_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_31_16_19 SB_T1_SOUTH_SB_OUT_B17_sel_value(
		.I(config_reg_3_O),
		.O(SB_T1_SOUTH_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_31_19_20 SB_T1_WEST_SB_IN_B17_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_WEST_SB_IN_B17_enable_value_O)
	);
	FanoutHash_653384C8EF52B5E3 SB_T1_WEST_SB_IN_B17_fan_in(
		.E8(PondTop_input_width_17_num_1_enable),
		.E6(PE_input_width_17_num_3_enable),
		.E3(PE_input_width_17_num_0_enable),
		.I5(PE_input_width_17_num_2_ready),
		.S6(PE_input_width_17_num_3_out_sel),
		.E0(SB_T4_NORTH_SB_OUT_B17_enable_value_O),
		.S5(PE_input_width_17_num_2_out_sel),
		.I6(PE_input_width_17_num_3_ready),
		.I8(PondTop_input_width_17_num_1_ready),
		.S3(PE_input_width_17_num_0_out_sel),
		.S4(PE_input_width_17_num_1_out_sel),
		.I3(PE_input_width_17_num_0_ready),
		.I4(PE_input_width_17_num_1_ready),
		.S1(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T1_EAST_SB_OUT_B17_out_sel),
		.S8(PondTop_input_width_17_num_1_out_sel),
		.E2(SB_T1_EAST_SB_OUT_B17_enable_value_O),
		.E5(PE_input_width_17_num_2_enable),
		.E4(PE_input_width_17_num_1_enable),
		.I2(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
		.O(SB_T1_WEST_SB_IN_B17_fan_in_O),
		.S7(PondTop_input_width_17_num_0_out_sel),
		.E1(SB_T0_SOUTH_SB_OUT_B17_enable_value_O),
		.I7(PondTop_input_width_17_num_0_ready),
		.I0(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
		.E7(PondTop_input_width_17_num_0_enable)
	);
	wire [1:0] SB_T1_WEST_SB_OUT_B17_FANOUT_I;
	assign SB_T1_WEST_SB_OUT_B17_FANOUT_I = {REG_T1_WEST_B17$SplitFifo_17_inst0_ready0[0], RMUX_T1_WEST_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T1_WEST_SB_OUT_B17_FANOUT(
		.O(SB_T1_WEST_SB_OUT_B17_FANOUT_O),
		.I(SB_T1_WEST_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T1_WEST_B17_out_sel)
	);
	SliceWrapper_31_20_21 SB_T1_WEST_SB_OUT_B17_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_WEST_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_31_21_24 SB_T1_WEST_SB_OUT_B17_sel_value(
		.I(config_reg_3_O),
		.O(SB_T1_WEST_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_31_24_25 SB_T2_EAST_SB_IN_B17_enable_value(
		.I(config_reg_3_O),
		.O(SB_T2_EAST_SB_IN_B17_enable_value_O)
	);
	FanoutHash_5CD8077D054B887B SB_T2_EAST_SB_IN_B17_fan_in(
		.E8(PondTop_input_width_17_num_1_enable),
		.E6(PE_input_width_17_num_3_enable),
		.E3(PE_input_width_17_num_0_enable),
		.I5(PE_input_width_17_num_2_ready),
		.S6(PE_input_width_17_num_3_out_sel),
		.E0(SB_T1_NORTH_SB_OUT_B17_enable_value_O),
		.S5(PE_input_width_17_num_2_out_sel),
		.I6(PE_input_width_17_num_3_ready),
		.I8(PondTop_input_width_17_num_1_ready),
		.S3(PE_input_width_17_num_0_out_sel),
		.S4(PE_input_width_17_num_1_out_sel),
		.I3(PE_input_width_17_num_0_ready),
		.I4(PE_input_width_17_num_1_ready),
		.S1(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T2_WEST_SB_OUT_B17_out_sel),
		.S8(PondTop_input_width_17_num_1_out_sel),
		.E2(SB_T2_WEST_SB_OUT_B17_enable_value_O),
		.E5(PE_input_width_17_num_2_enable),
		.E4(PE_input_width_17_num_1_enable),
		.I2(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
		.O(SB_T2_EAST_SB_IN_B17_fan_in_O),
		.S7(PondTop_input_width_17_num_0_out_sel),
		.E1(SB_T1_SOUTH_SB_OUT_B17_enable_value_O),
		.I7(PondTop_input_width_17_num_0_ready),
		.I0(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out),
		.E7(PondTop_input_width_17_num_0_enable)
	);
	wire [1:0] SB_T2_EAST_SB_OUT_B17_FANOUT_I;
	assign SB_T2_EAST_SB_OUT_B17_FANOUT_I = {REG_T2_EAST_B17$SplitFifo_17_inst0_ready0[0], RMUX_T2_EAST_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T2_EAST_SB_OUT_B17_FANOUT(
		.O(SB_T2_EAST_SB_OUT_B17_FANOUT_O),
		.I(SB_T2_EAST_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T2_EAST_B17_out_sel)
	);
	SliceWrapper_31_25_26 SB_T2_EAST_SB_OUT_B17_enable_value(
		.I(config_reg_3_O),
		.O(SB_T2_EAST_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_31_26_29 SB_T2_EAST_SB_OUT_B17_sel_value(
		.I(config_reg_3_O),
		.O(SB_T2_EAST_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_31_29_30 SB_T2_NORTH_SB_IN_B17_enable_value(
		.I(config_reg_3_O),
		.O(SB_T2_NORTH_SB_IN_B17_enable_value_O)
	);
	FanoutHash_74A3E41836ECED62 SB_T2_NORTH_SB_IN_B17_fan_in(
		.E8(PondTop_input_width_17_num_1_enable),
		.E6(PE_input_width_17_num_3_enable),
		.E3(PE_input_width_17_num_0_enable),
		.I5(PE_input_width_17_num_2_ready),
		.S6(PE_input_width_17_num_3_out_sel),
		.E0(SB_T3_EAST_SB_OUT_B17_enable_value_O),
		.S5(PE_input_width_17_num_2_out_sel),
		.I6(PE_input_width_17_num_3_ready),
		.I8(PondTop_input_width_17_num_1_ready),
		.S3(PE_input_width_17_num_0_out_sel),
		.S4(PE_input_width_17_num_1_out_sel),
		.I3(PE_input_width_17_num_0_ready),
		.I4(PE_input_width_17_num_1_ready),
		.S1(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T3_EAST_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T3_WEST_SB_OUT_B17_out_sel),
		.S8(PondTop_input_width_17_num_1_out_sel),
		.E2(SB_T3_WEST_SB_OUT_B17_enable_value_O),
		.E5(PE_input_width_17_num_2_enable),
		.E4(PE_input_width_17_num_1_enable),
		.I2(MUX_SB_T3_WEST_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
		.O(SB_T2_NORTH_SB_IN_B17_fan_in_O),
		.S7(PondTop_input_width_17_num_0_out_sel),
		.E1(SB_T2_SOUTH_SB_OUT_B17_enable_value_O),
		.I7(PondTop_input_width_17_num_0_ready),
		.I0(MUX_SB_T3_EAST_SB_OUT_B17_ready_out),
		.E7(PondTop_input_width_17_num_0_enable)
	);
	wire [1:0] SB_T2_NORTH_SB_OUT_B17_FANOUT_I;
	assign SB_T2_NORTH_SB_OUT_B17_FANOUT_I = {REG_T2_NORTH_B17$SplitFifo_17_inst0_ready0[0], RMUX_T2_NORTH_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T2_NORTH_SB_OUT_B17_FANOUT(
		.O(SB_T2_NORTH_SB_OUT_B17_FANOUT_O),
		.I(SB_T2_NORTH_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T2_NORTH_B17_out_sel)
	);
	SliceWrapper_31_30_31 SB_T2_NORTH_SB_OUT_B17_enable_value(
		.I(config_reg_3_O),
		.O(SB_T2_NORTH_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_30_0_3 SB_T2_NORTH_SB_OUT_B17_sel_value(
		.I(config_reg_4_O),
		.O(SB_T2_NORTH_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_30_3_4 SB_T2_SOUTH_SB_IN_B17_enable_value(
		.I(config_reg_4_O),
		.O(SB_T2_SOUTH_SB_IN_B17_enable_value_O)
	);
	FanoutHash_2CE3041FDDDDEC1A SB_T2_SOUTH_SB_IN_B17_fan_in(
		.E8(PondTop_input_width_17_num_1_enable),
		.E6(PE_input_width_17_num_3_enable),
		.E3(PE_input_width_17_num_0_enable),
		.I5(PE_input_width_17_num_2_ready),
		.S6(PE_input_width_17_num_3_out_sel),
		.E0(SB_T1_EAST_SB_OUT_B17_enable_value_O),
		.S5(PE_input_width_17_num_2_out_sel),
		.I6(PE_input_width_17_num_3_ready),
		.I8(PondTop_input_width_17_num_1_ready),
		.S3(PE_input_width_17_num_0_out_sel),
		.S4(PE_input_width_17_num_1_out_sel),
		.I3(PE_input_width_17_num_0_ready),
		.I4(PE_input_width_17_num_1_ready),
		.S1(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T1_EAST_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T3_WEST_SB_OUT_B17_out_sel),
		.S8(PondTop_input_width_17_num_1_out_sel),
		.E2(SB_T3_WEST_SB_OUT_B17_enable_value_O),
		.E5(PE_input_width_17_num_2_enable),
		.E4(PE_input_width_17_num_1_enable),
		.I2(MUX_SB_T3_WEST_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
		.O(SB_T2_SOUTH_SB_IN_B17_fan_in_O),
		.S7(PondTop_input_width_17_num_0_out_sel),
		.E1(SB_T2_NORTH_SB_OUT_B17_enable_value_O),
		.I7(PondTop_input_width_17_num_0_ready),
		.I0(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
		.E7(PondTop_input_width_17_num_0_enable)
	);
	wire [1:0] SB_T2_SOUTH_SB_OUT_B17_FANOUT_I;
	assign SB_T2_SOUTH_SB_OUT_B17_FANOUT_I = {REG_T2_SOUTH_B17$SplitFifo_17_inst0_ready0[0], RMUX_T2_SOUTH_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T2_SOUTH_SB_OUT_B17_FANOUT(
		.O(SB_T2_SOUTH_SB_OUT_B17_FANOUT_O),
		.I(SB_T2_SOUTH_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T2_SOUTH_B17_out_sel)
	);
	SliceWrapper_30_4_5 SB_T2_SOUTH_SB_OUT_B17_enable_value(
		.I(config_reg_4_O),
		.O(SB_T2_SOUTH_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_30_5_8 SB_T2_SOUTH_SB_OUT_B17_sel_value(
		.I(config_reg_4_O),
		.O(SB_T2_SOUTH_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_30_8_9 SB_T2_WEST_SB_IN_B17_enable_value(
		.I(config_reg_4_O),
		.O(SB_T2_WEST_SB_IN_B17_enable_value_O)
	);
	FanoutHash_4A74B16B611BA7E4 SB_T2_WEST_SB_IN_B17_fan_in(
		.E8(PondTop_input_width_17_num_1_enable),
		.E6(PE_input_width_17_num_3_enable),
		.E3(PE_input_width_17_num_0_enable),
		.I5(PE_input_width_17_num_2_ready),
		.S6(PE_input_width_17_num_3_out_sel),
		.E0(SB_T3_NORTH_SB_OUT_B17_enable_value_O),
		.S5(PE_input_width_17_num_2_out_sel),
		.I6(PE_input_width_17_num_3_ready),
		.I8(PondTop_input_width_17_num_1_ready),
		.S3(PE_input_width_17_num_0_out_sel),
		.S4(PE_input_width_17_num_1_out_sel),
		.I3(PE_input_width_17_num_0_ready),
		.I4(PE_input_width_17_num_1_ready),
		.S1(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T2_EAST_SB_OUT_B17_out_sel),
		.S8(PondTop_input_width_17_num_1_out_sel),
		.E2(SB_T2_EAST_SB_OUT_B17_enable_value_O),
		.E5(PE_input_width_17_num_2_enable),
		.E4(PE_input_width_17_num_1_enable),
		.I2(MUX_SB_T2_EAST_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
		.O(SB_T2_WEST_SB_IN_B17_fan_in_O),
		.S7(PondTop_input_width_17_num_0_out_sel),
		.E1(SB_T1_SOUTH_SB_OUT_B17_enable_value_O),
		.I7(PondTop_input_width_17_num_0_ready),
		.I0(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out),
		.E7(PondTop_input_width_17_num_0_enable)
	);
	wire [1:0] SB_T2_WEST_SB_OUT_B17_FANOUT_I;
	assign SB_T2_WEST_SB_OUT_B17_FANOUT_I = {REG_T2_WEST_B17$SplitFifo_17_inst0_ready0[0], RMUX_T2_WEST_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T2_WEST_SB_OUT_B17_FANOUT(
		.O(SB_T2_WEST_SB_OUT_B17_FANOUT_O),
		.I(SB_T2_WEST_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T2_WEST_B17_out_sel)
	);
	SliceWrapper_30_9_10 SB_T2_WEST_SB_OUT_B17_enable_value(
		.I(config_reg_4_O),
		.O(SB_T2_WEST_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_30_10_13 SB_T2_WEST_SB_OUT_B17_sel_value(
		.I(config_reg_4_O),
		.O(SB_T2_WEST_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_30_13_14 SB_T3_EAST_SB_IN_B17_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_EAST_SB_IN_B17_enable_value_O)
	);
	FanoutHash_276F8381CE025648 SB_T3_EAST_SB_IN_B17_fan_in(
		.E8(PondTop_input_width_17_num_1_enable),
		.E6(PE_input_width_17_num_3_enable),
		.E3(PE_input_width_17_num_0_enable),
		.I5(PE_input_width_17_num_2_ready),
		.S6(PE_input_width_17_num_3_out_sel),
		.E0(SB_T0_SOUTH_SB_OUT_B17_enable_value_O),
		.S5(PE_input_width_17_num_2_out_sel),
		.I6(PE_input_width_17_num_3_ready),
		.I8(PondTop_input_width_17_num_1_ready),
		.S3(PE_input_width_17_num_0_out_sel),
		.S4(PE_input_width_17_num_1_out_sel),
		.I3(PE_input_width_17_num_0_ready),
		.I4(PE_input_width_17_num_1_ready),
		.S1(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T3_WEST_SB_OUT_B17_out_sel),
		.S8(PondTop_input_width_17_num_1_out_sel),
		.E2(SB_T3_WEST_SB_OUT_B17_enable_value_O),
		.E5(PE_input_width_17_num_2_enable),
		.E4(PE_input_width_17_num_1_enable),
		.I2(MUX_SB_T3_WEST_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
		.O(SB_T3_EAST_SB_IN_B17_fan_in_O),
		.S7(PondTop_input_width_17_num_0_out_sel),
		.E1(SB_T2_NORTH_SB_OUT_B17_enable_value_O),
		.I7(PondTop_input_width_17_num_0_ready),
		.I0(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
		.E7(PondTop_input_width_17_num_0_enable)
	);
	wire [1:0] SB_T3_EAST_SB_OUT_B17_FANOUT_I;
	assign SB_T3_EAST_SB_OUT_B17_FANOUT_I = {REG_T3_EAST_B17$SplitFifo_17_inst0_ready0[0], RMUX_T3_EAST_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T3_EAST_SB_OUT_B17_FANOUT(
		.O(SB_T3_EAST_SB_OUT_B17_FANOUT_O),
		.I(SB_T3_EAST_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T3_EAST_B17_out_sel)
	);
	SliceWrapper_30_14_15 SB_T3_EAST_SB_OUT_B17_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_EAST_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_30_15_18 SB_T3_EAST_SB_OUT_B17_sel_value(
		.I(config_reg_4_O),
		.O(SB_T3_EAST_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_30_18_19 SB_T3_NORTH_SB_IN_B17_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_NORTH_SB_IN_B17_enable_value_O)
	);
	FanoutHash_7E22D83B42537D1D SB_T3_NORTH_SB_IN_B17_fan_in(
		.E8(PondTop_input_width_17_num_1_enable),
		.E6(PE_input_width_17_num_3_enable),
		.E3(PE_input_width_17_num_0_enable),
		.I5(PE_input_width_17_num_2_ready),
		.S6(PE_input_width_17_num_3_out_sel),
		.E0(SB_T2_WEST_SB_OUT_B17_enable_value_O),
		.S5(PE_input_width_17_num_2_out_sel),
		.I6(PE_input_width_17_num_3_ready),
		.I8(PondTop_input_width_17_num_1_ready),
		.S3(PE_input_width_17_num_0_out_sel),
		.S4(PE_input_width_17_num_1_out_sel),
		.I3(PE_input_width_17_num_0_ready),
		.I4(PE_input_width_17_num_1_ready),
		.S1(MUX_SB_T4_EAST_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T2_WEST_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel),
		.S8(PondTop_input_width_17_num_1_out_sel),
		.E2(SB_T3_SOUTH_SB_OUT_B17_enable_value_O),
		.E5(PE_input_width_17_num_2_enable),
		.E4(PE_input_width_17_num_1_enable),
		.I2(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T4_EAST_SB_OUT_B17_ready_out),
		.O(SB_T3_NORTH_SB_IN_B17_fan_in_O),
		.S7(PondTop_input_width_17_num_0_out_sel),
		.E1(SB_T4_EAST_SB_OUT_B17_enable_value_O),
		.I7(PondTop_input_width_17_num_0_ready),
		.I0(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
		.E7(PondTop_input_width_17_num_0_enable)
	);
	wire [1:0] SB_T3_NORTH_SB_OUT_B17_FANOUT_I;
	assign SB_T3_NORTH_SB_OUT_B17_FANOUT_I = {REG_T3_NORTH_B17$SplitFifo_17_inst0_ready0[0], RMUX_T3_NORTH_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T3_NORTH_SB_OUT_B17_FANOUT(
		.O(SB_T3_NORTH_SB_OUT_B17_FANOUT_O),
		.I(SB_T3_NORTH_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T3_NORTH_B17_out_sel)
	);
	SliceWrapper_30_19_20 SB_T3_NORTH_SB_OUT_B17_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_NORTH_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_30_20_23 SB_T3_NORTH_SB_OUT_B17_sel_value(
		.I(config_reg_4_O),
		.O(SB_T3_NORTH_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_30_23_24 SB_T3_SOUTH_SB_IN_B17_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_SOUTH_SB_IN_B17_enable_value_O)
	);
	FanoutHash_59B7E37DAE2221E3 SB_T3_SOUTH_SB_IN_B17_fan_in(
		.E8(PondTop_input_width_17_num_1_enable),
		.E6(PE_input_width_17_num_3_enable),
		.E3(PE_input_width_17_num_0_enable),
		.I5(PE_input_width_17_num_2_ready),
		.S6(PE_input_width_17_num_3_out_sel),
		.E0(SB_T0_EAST_SB_OUT_B17_enable_value_O),
		.S5(PE_input_width_17_num_2_out_sel),
		.I6(PE_input_width_17_num_3_ready),
		.I8(PondTop_input_width_17_num_1_ready),
		.S3(PE_input_width_17_num_0_out_sel),
		.S4(PE_input_width_17_num_1_out_sel),
		.I3(PE_input_width_17_num_0_ready),
		.I4(PE_input_width_17_num_1_ready),
		.S1(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T0_EAST_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T4_WEST_SB_OUT_B17_out_sel),
		.S8(PondTop_input_width_17_num_1_out_sel),
		.E2(SB_T4_WEST_SB_OUT_B17_enable_value_O),
		.E5(PE_input_width_17_num_2_enable),
		.E4(PE_input_width_17_num_1_enable),
		.I2(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out),
		.O(SB_T3_SOUTH_SB_IN_B17_fan_in_O),
		.S7(PondTop_input_width_17_num_0_out_sel),
		.E1(SB_T3_NORTH_SB_OUT_B17_enable_value_O),
		.I7(PondTop_input_width_17_num_0_ready),
		.I0(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
		.E7(PondTop_input_width_17_num_0_enable)
	);
	wire [1:0] SB_T3_SOUTH_SB_OUT_B17_FANOUT_I;
	assign SB_T3_SOUTH_SB_OUT_B17_FANOUT_I = {REG_T3_SOUTH_B17$SplitFifo_17_inst0_ready0[0], RMUX_T3_SOUTH_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T3_SOUTH_SB_OUT_B17_FANOUT(
		.O(SB_T3_SOUTH_SB_OUT_B17_FANOUT_O),
		.I(SB_T3_SOUTH_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T3_SOUTH_B17_out_sel)
	);
	SliceWrapper_30_24_25 SB_T3_SOUTH_SB_OUT_B17_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_SOUTH_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_30_25_28 SB_T3_SOUTH_SB_OUT_B17_sel_value(
		.I(config_reg_4_O),
		.O(SB_T3_SOUTH_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_30_28_29 SB_T3_WEST_SB_IN_B17_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_WEST_SB_IN_B17_enable_value_O)
	);
	FanoutHash_41D739158D58E184 SB_T3_WEST_SB_IN_B17_fan_in(
		.E8(PondTop_input_width_17_num_1_enable),
		.E6(PE_input_width_17_num_3_enable),
		.E3(PE_input_width_17_num_0_enable),
		.I5(PE_input_width_17_num_2_ready),
		.S6(PE_input_width_17_num_3_out_sel),
		.E0(SB_T2_NORTH_SB_OUT_B17_enable_value_O),
		.S5(PE_input_width_17_num_2_out_sel),
		.I6(PE_input_width_17_num_3_ready),
		.I8(PondTop_input_width_17_num_1_ready),
		.S3(PE_input_width_17_num_0_out_sel),
		.S4(PE_input_width_17_num_1_out_sel),
		.I3(PE_input_width_17_num_0_ready),
		.I4(PE_input_width_17_num_1_ready),
		.S1(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T3_EAST_SB_OUT_B17_out_sel),
		.S8(PondTop_input_width_17_num_1_out_sel),
		.E2(SB_T3_EAST_SB_OUT_B17_enable_value_O),
		.E5(PE_input_width_17_num_2_enable),
		.E4(PE_input_width_17_num_1_enable),
		.I2(MUX_SB_T3_EAST_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
		.O(SB_T3_WEST_SB_IN_B17_fan_in_O),
		.S7(PondTop_input_width_17_num_0_out_sel),
		.E1(SB_T2_SOUTH_SB_OUT_B17_enable_value_O),
		.I7(PondTop_input_width_17_num_0_ready),
		.I0(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
		.E7(PondTop_input_width_17_num_0_enable)
	);
	wire [1:0] SB_T3_WEST_SB_OUT_B17_FANOUT_I;
	assign SB_T3_WEST_SB_OUT_B17_FANOUT_I = {REG_T3_WEST_B17$SplitFifo_17_inst0_ready0[0], RMUX_T3_WEST_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T3_WEST_SB_OUT_B17_FANOUT(
		.O(SB_T3_WEST_SB_OUT_B17_FANOUT_O),
		.I(SB_T3_WEST_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T3_WEST_B17_out_sel)
	);
	SliceWrapper_30_29_30 SB_T3_WEST_SB_OUT_B17_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_WEST_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_23_0_3 SB_T3_WEST_SB_OUT_B17_sel_value(
		.I(config_reg_5_O),
		.O(SB_T3_WEST_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_23_3_4 SB_T4_EAST_SB_IN_B17_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_EAST_SB_IN_B17_enable_value_O)
	);
	FanoutHash_55169EB19E10AA09 SB_T4_EAST_SB_IN_B17_fan_in(
		.E8(PondTop_input_width_17_num_1_enable),
		.E6(PE_input_width_17_num_3_enable),
		.E3(PE_input_width_17_num_0_enable),
		.I5(PE_input_width_17_num_2_ready),
		.S6(PE_input_width_17_num_3_out_sel),
		.E0(SB_T3_NORTH_SB_OUT_B17_enable_value_O),
		.S5(PE_input_width_17_num_2_out_sel),
		.I6(PE_input_width_17_num_3_ready),
		.I8(PondTop_input_width_17_num_1_ready),
		.S3(PE_input_width_17_num_0_out_sel),
		.S4(PE_input_width_17_num_1_out_sel),
		.I3(PE_input_width_17_num_0_ready),
		.I4(PE_input_width_17_num_1_ready),
		.S1(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T4_WEST_SB_OUT_B17_out_sel),
		.S8(PondTop_input_width_17_num_1_out_sel),
		.E2(SB_T4_WEST_SB_OUT_B17_enable_value_O),
		.E5(PE_input_width_17_num_2_enable),
		.E4(PE_input_width_17_num_1_enable),
		.I2(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
		.O(SB_T4_EAST_SB_IN_B17_fan_in_O),
		.S7(PondTop_input_width_17_num_0_out_sel),
		.E1(SB_T4_SOUTH_SB_OUT_B17_enable_value_O),
		.I7(PondTop_input_width_17_num_0_ready),
		.I0(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out),
		.E7(PondTop_input_width_17_num_0_enable)
	);
	wire [1:0] SB_T4_EAST_SB_OUT_B17_FANOUT_I;
	assign SB_T4_EAST_SB_OUT_B17_FANOUT_I = {REG_T4_EAST_B17$SplitFifo_17_inst0_ready0[0], RMUX_T4_EAST_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T4_EAST_SB_OUT_B17_FANOUT(
		.O(SB_T4_EAST_SB_OUT_B17_FANOUT_O),
		.I(SB_T4_EAST_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T4_EAST_B17_out_sel)
	);
	SliceWrapper_23_4_5 SB_T4_EAST_SB_OUT_B17_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_EAST_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_23_5_8 SB_T4_EAST_SB_OUT_B17_sel_value(
		.I(config_reg_5_O),
		.O(SB_T4_EAST_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_23_8_9 SB_T4_NORTH_SB_IN_B17_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_NORTH_SB_IN_B17_enable_value_O)
	);
	FanoutHash_244497FCED8BEB80 SB_T4_NORTH_SB_IN_B17_fan_in(
		.E8(PondTop_input_width_17_num_1_enable),
		.E6(PE_input_width_17_num_3_enable),
		.E3(PE_input_width_17_num_0_enable),
		.I5(PE_input_width_17_num_2_ready),
		.S6(PE_input_width_17_num_3_out_sel),
		.E0(SB_T1_WEST_SB_OUT_B17_enable_value_O),
		.S5(PE_input_width_17_num_2_out_sel),
		.I6(PE_input_width_17_num_3_ready),
		.I8(PondTop_input_width_17_num_1_ready),
		.S3(PE_input_width_17_num_0_out_sel),
		.S4(PE_input_width_17_num_1_out_sel),
		.I3(PE_input_width_17_num_0_ready),
		.I4(PE_input_width_17_num_1_ready),
		.S1(MUX_SB_T0_EAST_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T1_WEST_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel),
		.S8(PondTop_input_width_17_num_1_out_sel),
		.E2(SB_T4_SOUTH_SB_OUT_B17_enable_value_O),
		.E5(PE_input_width_17_num_2_enable),
		.E4(PE_input_width_17_num_1_enable),
		.I2(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
		.O(SB_T4_NORTH_SB_IN_B17_fan_in_O),
		.S7(PondTop_input_width_17_num_0_out_sel),
		.E1(SB_T0_EAST_SB_OUT_B17_enable_value_O),
		.I7(PondTop_input_width_17_num_0_ready),
		.I0(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
		.E7(PondTop_input_width_17_num_0_enable)
	);
	wire [1:0] SB_T4_NORTH_SB_OUT_B17_FANOUT_I;
	assign SB_T4_NORTH_SB_OUT_B17_FANOUT_I = {REG_T4_NORTH_B17$SplitFifo_17_inst0_ready0[0], RMUX_T4_NORTH_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T4_NORTH_SB_OUT_B17_FANOUT(
		.O(SB_T4_NORTH_SB_OUT_B17_FANOUT_O),
		.I(SB_T4_NORTH_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T4_NORTH_B17_out_sel)
	);
	SliceWrapper_23_9_10 SB_T4_NORTH_SB_OUT_B17_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_NORTH_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_23_10_13 SB_T4_NORTH_SB_OUT_B17_sel_value(
		.I(config_reg_5_O),
		.O(SB_T4_NORTH_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_23_13_14 SB_T4_SOUTH_SB_IN_B17_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_SOUTH_SB_IN_B17_enable_value_O)
	);
	FanoutHash_AE7392256DF8B0F SB_T4_SOUTH_SB_IN_B17_fan_in(
		.E8(PondTop_input_width_17_num_1_enable),
		.E6(PE_input_width_17_num_3_enable),
		.E3(PE_input_width_17_num_0_enable),
		.I5(PE_input_width_17_num_2_ready),
		.S6(PE_input_width_17_num_3_out_sel),
		.E0(SB_T0_WEST_SB_OUT_B17_enable_value_O),
		.S5(PE_input_width_17_num_2_out_sel),
		.I6(PE_input_width_17_num_3_ready),
		.I8(PondTop_input_width_17_num_1_ready),
		.S3(PE_input_width_17_num_0_out_sel),
		.S4(PE_input_width_17_num_1_out_sel),
		.I3(PE_input_width_17_num_0_ready),
		.I4(PE_input_width_17_num_1_ready),
		.S1(MUX_SB_T4_EAST_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T0_WEST_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel),
		.S8(PondTop_input_width_17_num_1_out_sel),
		.E2(SB_T4_NORTH_SB_OUT_B17_enable_value_O),
		.E5(PE_input_width_17_num_2_enable),
		.E4(PE_input_width_17_num_1_enable),
		.I2(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T4_EAST_SB_OUT_B17_ready_out),
		.O(SB_T4_SOUTH_SB_IN_B17_fan_in_O),
		.S7(PondTop_input_width_17_num_0_out_sel),
		.E1(SB_T4_EAST_SB_OUT_B17_enable_value_O),
		.I7(PondTop_input_width_17_num_0_ready),
		.I0(MUX_SB_T0_WEST_SB_OUT_B17_ready_out),
		.E7(PondTop_input_width_17_num_0_enable)
	);
	wire [1:0] SB_T4_SOUTH_SB_OUT_B17_FANOUT_I;
	assign SB_T4_SOUTH_SB_OUT_B17_FANOUT_I = {REG_T4_SOUTH_B17$SplitFifo_17_inst0_ready0[0], RMUX_T4_SOUTH_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T4_SOUTH_SB_OUT_B17_FANOUT(
		.O(SB_T4_SOUTH_SB_OUT_B17_FANOUT_O),
		.I(SB_T4_SOUTH_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T4_SOUTH_B17_out_sel)
	);
	SliceWrapper_23_14_15 SB_T4_SOUTH_SB_OUT_B17_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_SOUTH_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_23_15_18 SB_T4_SOUTH_SB_OUT_B17_sel_value(
		.I(config_reg_5_O),
		.O(SB_T4_SOUTH_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_23_18_19 SB_T4_WEST_SB_IN_B17_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_WEST_SB_IN_B17_enable_value_O)
	);
	FanoutHash_6E1094CE0D0F6DFA SB_T4_WEST_SB_IN_B17_fan_in(
		.E8(PondTop_input_width_17_num_1_enable),
		.E6(PE_input_width_17_num_3_enable),
		.E3(PE_input_width_17_num_0_enable),
		.I5(PE_input_width_17_num_2_ready),
		.S6(PE_input_width_17_num_3_out_sel),
		.E0(SB_T1_NORTH_SB_OUT_B17_enable_value_O),
		.S5(PE_input_width_17_num_2_out_sel),
		.I6(PE_input_width_17_num_3_ready),
		.I8(PondTop_input_width_17_num_1_ready),
		.S3(PE_input_width_17_num_0_out_sel),
		.S4(PE_input_width_17_num_1_out_sel),
		.I3(PE_input_width_17_num_0_ready),
		.I4(PE_input_width_17_num_1_ready),
		.S1(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T4_EAST_SB_OUT_B17_out_sel),
		.S8(PondTop_input_width_17_num_1_out_sel),
		.E2(SB_T4_EAST_SB_OUT_B17_enable_value_O),
		.E5(PE_input_width_17_num_2_enable),
		.E4(PE_input_width_17_num_1_enable),
		.I2(MUX_SB_T4_EAST_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
		.O(SB_T4_WEST_SB_IN_B17_fan_in_O),
		.S7(PondTop_input_width_17_num_0_out_sel),
		.E1(SB_T3_SOUTH_SB_OUT_B17_enable_value_O),
		.I7(PondTop_input_width_17_num_0_ready),
		.I0(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out),
		.E7(PondTop_input_width_17_num_0_enable)
	);
	wire [1:0] SB_T4_WEST_SB_OUT_B17_FANOUT_I;
	assign SB_T4_WEST_SB_OUT_B17_FANOUT_I = {REG_T4_WEST_B17$SplitFifo_17_inst0_ready0[0], RMUX_T4_WEST_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T4_WEST_SB_OUT_B17_FANOUT(
		.O(SB_T4_WEST_SB_OUT_B17_FANOUT_O),
		.I(SB_T4_WEST_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T4_WEST_B17_out_sel)
	);
	SliceWrapper_23_19_20 SB_T4_WEST_SB_OUT_B17_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_WEST_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_23_20_23 SB_T4_WEST_SB_OUT_B17_sel_value(
		.I(config_reg_5_O),
		.O(SB_T4_WEST_SB_OUT_B17_sel_value_O)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T0_EAST_SB_IN_B17(
		.I(SB_T0_EAST_SB_IN_B17),
		.O(WIRE_SB_T0_EAST_SB_IN_B17_O),
		.ready_in(SB_T0_EAST_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T0_EAST_SB_IN_B17_ready_out),
		.valid_in(SB_T0_EAST_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T0_EAST_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T0_NORTH_SB_IN_B17(
		.I(SB_T0_NORTH_SB_IN_B17),
		.O(WIRE_SB_T0_NORTH_SB_IN_B17_O),
		.ready_in(SB_T0_NORTH_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T0_NORTH_SB_IN_B17_ready_out),
		.valid_in(SB_T0_NORTH_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T0_NORTH_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T0_SOUTH_SB_IN_B17(
		.I(SB_T0_SOUTH_SB_IN_B17),
		.O(WIRE_SB_T0_SOUTH_SB_IN_B17_O),
		.ready_in(SB_T0_SOUTH_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T0_SOUTH_SB_IN_B17_ready_out),
		.valid_in(SB_T0_SOUTH_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T0_SOUTH_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T0_WEST_SB_IN_B17(
		.I(SB_T0_WEST_SB_IN_B17),
		.O(WIRE_SB_T0_WEST_SB_IN_B17_O),
		.ready_in(SB_T0_WEST_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T0_WEST_SB_IN_B17_ready_out),
		.valid_in(SB_T0_WEST_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T0_WEST_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T1_EAST_SB_IN_B17(
		.I(SB_T1_EAST_SB_IN_B17),
		.O(WIRE_SB_T1_EAST_SB_IN_B17_O),
		.ready_in(SB_T1_EAST_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T1_EAST_SB_IN_B17_ready_out),
		.valid_in(SB_T1_EAST_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T1_EAST_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T1_NORTH_SB_IN_B17(
		.I(SB_T1_NORTH_SB_IN_B17),
		.O(WIRE_SB_T1_NORTH_SB_IN_B17_O),
		.ready_in(SB_T1_NORTH_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T1_NORTH_SB_IN_B17_ready_out),
		.valid_in(SB_T1_NORTH_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T1_NORTH_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T1_SOUTH_SB_IN_B17(
		.I(SB_T1_SOUTH_SB_IN_B17),
		.O(WIRE_SB_T1_SOUTH_SB_IN_B17_O),
		.ready_in(SB_T1_SOUTH_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T1_SOUTH_SB_IN_B17_ready_out),
		.valid_in(SB_T1_SOUTH_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T1_SOUTH_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T1_WEST_SB_IN_B17(
		.I(SB_T1_WEST_SB_IN_B17),
		.O(WIRE_SB_T1_WEST_SB_IN_B17_O),
		.ready_in(SB_T1_WEST_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T1_WEST_SB_IN_B17_ready_out),
		.valid_in(SB_T1_WEST_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T1_WEST_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T2_EAST_SB_IN_B17(
		.I(SB_T2_EAST_SB_IN_B17),
		.O(WIRE_SB_T2_EAST_SB_IN_B17_O),
		.ready_in(SB_T2_EAST_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T2_EAST_SB_IN_B17_ready_out),
		.valid_in(SB_T2_EAST_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T2_EAST_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T2_NORTH_SB_IN_B17(
		.I(SB_T2_NORTH_SB_IN_B17),
		.O(WIRE_SB_T2_NORTH_SB_IN_B17_O),
		.ready_in(SB_T2_NORTH_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T2_NORTH_SB_IN_B17_ready_out),
		.valid_in(SB_T2_NORTH_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T2_NORTH_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T2_SOUTH_SB_IN_B17(
		.I(SB_T2_SOUTH_SB_IN_B17),
		.O(WIRE_SB_T2_SOUTH_SB_IN_B17_O),
		.ready_in(SB_T2_SOUTH_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T2_SOUTH_SB_IN_B17_ready_out),
		.valid_in(SB_T2_SOUTH_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T2_SOUTH_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T2_WEST_SB_IN_B17(
		.I(SB_T2_WEST_SB_IN_B17),
		.O(WIRE_SB_T2_WEST_SB_IN_B17_O),
		.ready_in(SB_T2_WEST_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T2_WEST_SB_IN_B17_ready_out),
		.valid_in(SB_T2_WEST_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T2_WEST_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T3_EAST_SB_IN_B17(
		.I(SB_T3_EAST_SB_IN_B17),
		.O(WIRE_SB_T3_EAST_SB_IN_B17_O),
		.ready_in(SB_T3_EAST_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T3_EAST_SB_IN_B17_ready_out),
		.valid_in(SB_T3_EAST_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T3_EAST_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T3_NORTH_SB_IN_B17(
		.I(SB_T3_NORTH_SB_IN_B17),
		.O(WIRE_SB_T3_NORTH_SB_IN_B17_O),
		.ready_in(SB_T3_NORTH_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T3_NORTH_SB_IN_B17_ready_out),
		.valid_in(SB_T3_NORTH_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T3_NORTH_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T3_SOUTH_SB_IN_B17(
		.I(SB_T3_SOUTH_SB_IN_B17),
		.O(WIRE_SB_T3_SOUTH_SB_IN_B17_O),
		.ready_in(SB_T3_SOUTH_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T3_SOUTH_SB_IN_B17_ready_out),
		.valid_in(SB_T3_SOUTH_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T3_SOUTH_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T3_WEST_SB_IN_B17(
		.I(SB_T3_WEST_SB_IN_B17),
		.O(WIRE_SB_T3_WEST_SB_IN_B17_O),
		.ready_in(SB_T3_WEST_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T3_WEST_SB_IN_B17_ready_out),
		.valid_in(SB_T3_WEST_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T3_WEST_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T4_EAST_SB_IN_B17(
		.I(SB_T4_EAST_SB_IN_B17),
		.O(WIRE_SB_T4_EAST_SB_IN_B17_O),
		.ready_in(SB_T4_EAST_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T4_EAST_SB_IN_B17_ready_out),
		.valid_in(SB_T4_EAST_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T4_EAST_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T4_NORTH_SB_IN_B17(
		.I(SB_T4_NORTH_SB_IN_B17),
		.O(WIRE_SB_T4_NORTH_SB_IN_B17_O),
		.ready_in(SB_T4_NORTH_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T4_NORTH_SB_IN_B17_ready_out),
		.valid_in(SB_T4_NORTH_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T4_NORTH_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T4_SOUTH_SB_IN_B17(
		.I(SB_T4_SOUTH_SB_IN_B17),
		.O(WIRE_SB_T4_SOUTH_SB_IN_B17_O),
		.ready_in(SB_T4_SOUTH_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T4_SOUTH_SB_IN_B17_ready_out),
		.valid_in(SB_T4_SOUTH_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T4_SOUTH_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T4_WEST_SB_IN_B17(
		.I(SB_T4_WEST_SB_IN_B17),
		.O(WIRE_SB_T4_WEST_SB_IN_B17_O),
		.ready_in(SB_T4_WEST_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T4_WEST_SB_IN_B17_ready_out),
		.valid_in(SB_T4_WEST_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T4_WEST_SB_IN_B17_valid_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_23_32_inst0$bit_const_0_None(.out(ZextWrapper_23_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_23_32_inst0$self_O_out;
	assign ZextWrapper_23_32_inst0$self_O_out = {ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, config_reg_5_O};
	mantle_wire__typeBitIn32 ZextWrapper_23_32_inst0$self_O(
		.in(ZextWrapper_23_32_inst0$self_O_in),
		.out(ZextWrapper_23_32_inst0$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_30_32_inst0$bit_const_0_None(.out(ZextWrapper_30_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_30_32_inst0$self_O_out;
	assign ZextWrapper_30_32_inst0$self_O_out = {ZextWrapper_30_32_inst0$bit_const_0_None_out, ZextWrapper_30_32_inst0$bit_const_0_None_out, config_reg_4_O};
	mantle_wire__typeBitIn32 ZextWrapper_30_32_inst0$self_O(
		.in(ZextWrapper_30_32_inst0$self_O_in),
		.out(ZextWrapper_30_32_inst0$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_31_32_inst0$bit_const_0_None(.out(ZextWrapper_31_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_31_32_inst0$self_O_out;
	assign ZextWrapper_31_32_inst0$self_O_out = {ZextWrapper_31_32_inst0$bit_const_0_None_out, config_reg_3_O};
	mantle_wire__typeBitIn32 ZextWrapper_31_32_inst0$self_O(
		.in(ZextWrapper_31_32_inst0$self_O_in),
		.out(ZextWrapper_31_32_inst0$self_O_out)
	);
	coreir_and #(.width(1)) and1_inst0(
		.in0(coreir_eq_1_inst0_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst0_out)
	);
	coreir_and #(.width(1)) and1_inst1(
		.in0(coreir_eq_1_inst1_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst1_out)
	);
	coreir_and #(.width(1)) and1_inst10(
		.in0(coreir_eq_1_inst10_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst10_out)
	);
	coreir_and #(.width(1)) and1_inst11(
		.in0(coreir_eq_1_inst11_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst11_out)
	);
	coreir_and #(.width(1)) and1_inst12(
		.in0(coreir_eq_1_inst12_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst12_out)
	);
	coreir_and #(.width(1)) and1_inst13(
		.in0(coreir_eq_1_inst13_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst13_out)
	);
	coreir_and #(.width(1)) and1_inst14(
		.in0(coreir_eq_1_inst14_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst14_out)
	);
	coreir_and #(.width(1)) and1_inst15(
		.in0(coreir_eq_1_inst15_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst15_out)
	);
	coreir_and #(.width(1)) and1_inst16(
		.in0(coreir_eq_1_inst16_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst16_out)
	);
	coreir_and #(.width(1)) and1_inst17(
		.in0(coreir_eq_1_inst17_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst17_out)
	);
	coreir_and #(.width(1)) and1_inst18(
		.in0(coreir_eq_1_inst18_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst18_out)
	);
	coreir_and #(.width(1)) and1_inst19(
		.in0(coreir_eq_1_inst19_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst19_out)
	);
	coreir_and #(.width(1)) and1_inst2(
		.in0(coreir_eq_1_inst2_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst2_out)
	);
	coreir_and #(.width(1)) and1_inst3(
		.in0(coreir_eq_1_inst3_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst3_out)
	);
	coreir_and #(.width(1)) and1_inst4(
		.in0(coreir_eq_1_inst4_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst4_out)
	);
	coreir_and #(.width(1)) and1_inst5(
		.in0(coreir_eq_1_inst5_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst5_out)
	);
	coreir_and #(.width(1)) and1_inst6(
		.in0(coreir_eq_1_inst6_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst6_out)
	);
	coreir_and #(.width(1)) and1_inst7(
		.in0(coreir_eq_1_inst7_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst7_out)
	);
	coreir_and #(.width(1)) and1_inst8(
		.in0(coreir_eq_1_inst8_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst8_out)
	);
	coreir_and #(.width(1)) and1_inst9(
		.in0(coreir_eq_1_inst9_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst9_out)
	);
	wire [7:0] config_reg_0_config_addr;
	assign config_reg_0_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4], self_config_config_addr_out[3], self_config_config_addr_out[2:0]};
	ConfigRegister_32_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_reg_0_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_1_config_addr;
	assign config_reg_1_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4], self_config_config_addr_out[3], self_config_config_addr_out[2:0]};
	ConfigRegister_32_8_32_1 config_reg_1(
		.clk(clk),
		.reset(reset),
		.O(config_reg_1_O),
		.config_addr(config_reg_1_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_2_config_addr;
	assign config_reg_2_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4], self_config_config_addr_out[3], self_config_config_addr_out[2:0]};
	ConfigRegister_32_8_32_2 config_reg_2(
		.clk(clk),
		.reset(reset),
		.O(config_reg_2_O),
		.config_addr(config_reg_2_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_3_config_addr;
	assign config_reg_3_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4], self_config_config_addr_out[3], self_config_config_addr_out[2:0]};
	ConfigRegister_31_8_32_3 config_reg_3(
		.clk(clk),
		.reset(reset),
		.O(config_reg_3_O),
		.config_addr(config_reg_3_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_4_config_addr;
	assign config_reg_4_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4], self_config_config_addr_out[3], self_config_config_addr_out[2:0]};
	ConfigRegister_30_8_32_4 config_reg_4(
		.clk(clk),
		.reset(reset),
		.O(config_reg_4_O),
		.config_addr(config_reg_4_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_5_config_addr;
	assign config_reg_5_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4], self_config_config_addr_out[3], self_config_config_addr_out[2:0]};
	ConfigRegister_23_8_32_5 config_reg_5(
		.clk(clk),
		.reset(reset),
		.O(config_reg_5_O),
		.config_addr(config_reg_5_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	coreir_const #(
		.value(1'h1),
		.width(1)
	) const_1_1(.out(const_1_1_out));
	coreir_eq #(.width(1)) coreir_eq_1_inst0(
		.in0(const_1_1_out),
		.in1(RMUX_T0_NORTH_B17_sel_value_O),
		.out(coreir_eq_1_inst0_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst1(
		.in0(const_1_1_out),
		.in1(RMUX_T0_SOUTH_B17_sel_value_O),
		.out(coreir_eq_1_inst1_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst10(
		.in0(const_1_1_out),
		.in1(RMUX_T2_EAST_B17_sel_value_O),
		.out(coreir_eq_1_inst10_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst11(
		.in0(const_1_1_out),
		.in1(RMUX_T2_WEST_B17_sel_value_O),
		.out(coreir_eq_1_inst11_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst12(
		.in0(const_1_1_out),
		.in1(RMUX_T3_NORTH_B17_sel_value_O),
		.out(coreir_eq_1_inst12_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst13(
		.in0(const_1_1_out),
		.in1(RMUX_T3_SOUTH_B17_sel_value_O),
		.out(coreir_eq_1_inst13_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst14(
		.in0(const_1_1_out),
		.in1(RMUX_T3_EAST_B17_sel_value_O),
		.out(coreir_eq_1_inst14_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst15(
		.in0(const_1_1_out),
		.in1(RMUX_T3_WEST_B17_sel_value_O),
		.out(coreir_eq_1_inst15_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst16(
		.in0(const_1_1_out),
		.in1(RMUX_T4_NORTH_B17_sel_value_O),
		.out(coreir_eq_1_inst16_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst17(
		.in0(const_1_1_out),
		.in1(RMUX_T4_SOUTH_B17_sel_value_O),
		.out(coreir_eq_1_inst17_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst18(
		.in0(const_1_1_out),
		.in1(RMUX_T4_EAST_B17_sel_value_O),
		.out(coreir_eq_1_inst18_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst19(
		.in0(const_1_1_out),
		.in1(RMUX_T4_WEST_B17_sel_value_O),
		.out(coreir_eq_1_inst19_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst2(
		.in0(const_1_1_out),
		.in1(RMUX_T0_EAST_B17_sel_value_O),
		.out(coreir_eq_1_inst2_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst3(
		.in0(const_1_1_out),
		.in1(RMUX_T0_WEST_B17_sel_value_O),
		.out(coreir_eq_1_inst3_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst4(
		.in0(const_1_1_out),
		.in1(RMUX_T1_NORTH_B17_sel_value_O),
		.out(coreir_eq_1_inst4_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst5(
		.in0(const_1_1_out),
		.in1(RMUX_T1_SOUTH_B17_sel_value_O),
		.out(coreir_eq_1_inst5_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst6(
		.in0(const_1_1_out),
		.in1(RMUX_T1_EAST_B17_sel_value_O),
		.out(coreir_eq_1_inst6_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst7(
		.in0(const_1_1_out),
		.in1(RMUX_T1_WEST_B17_sel_value_O),
		.out(coreir_eq_1_inst7_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst8(
		.in0(const_1_1_out),
		.in1(RMUX_T2_NORTH_B17_sel_value_O),
		.out(coreir_eq_1_inst8_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst9(
		.in0(const_1_1_out),
		.in1(RMUX_T2_SOUTH_B17_sel_value_O),
		.out(coreir_eq_1_inst9_out)
	);
	wire [191:0] mux_aoi_6_32_inst0_I;
	assign mux_aoi_6_32_inst0_I[160+:32] = ZextWrapper_23_32_inst0$self_O_in;
	assign mux_aoi_6_32_inst0_I[128+:32] = ZextWrapper_30_32_inst0$self_O_in;
	assign mux_aoi_6_32_inst0_I[96+:32] = ZextWrapper_31_32_inst0$self_O_in;
	assign mux_aoi_6_32_inst0_I[64+:32] = config_reg_2_O;
	assign mux_aoi_6_32_inst0_I[32+:32] = config_reg_1_O;
	assign mux_aoi_6_32_inst0_I[0+:32] = config_reg_0_O;
	mux_aoi_6_32 mux_aoi_6_32_inst0(
		.I(mux_aoi_6_32_inst0_I),
		.O(mux_aoi_6_32_inst0_O),
		.S(self_config_config_addr_out[2:0]),
		.out_sel(mux_aoi_6_32_inst0_out_sel)
	);
	mantle_wire__typeBit8 self_config_config_addr(
		.in(config_config_addr),
		.out(self_config_config_addr_out)
	);
	assign PE_output_width_17_num_0_ready_out = CB_PE_output_width_17_num_0_fan_in_O[0];
	assign PE_output_width_17_num_1_ready_out = CB_PE_output_width_17_num_1_fan_in_O[0];
	assign PE_output_width_17_num_2_ready_out = CB_PE_output_width_17_num_2_fan_in_O[0];
	assign PondTop_output_width_17_num_0_ready_out = CB_PondTop_output_width_17_num_0_fan_in_O[0];
	assign PondTop_output_width_17_num_1_ready_out = CB_PondTop_output_width_17_num_1_fan_in_O[0];
	assign SB_T0_EAST_SB_IN_B17_enable = SB_T0_EAST_SB_IN_B17_enable_value_O[0];
	assign SB_T0_EAST_SB_IN_B17_ready_out = WIRE_SB_T0_EAST_SB_IN_B17_ready_out;
	assign SB_T0_EAST_SB_OUT_B17 = RMUX_T0_EAST_B17_O;
	assign SB_T0_EAST_SB_OUT_B17_enable = SB_T0_EAST_SB_OUT_B17_enable_value_O[0];
	assign SB_T0_EAST_SB_OUT_B17_valid_out = RMUX_T0_EAST_B17_valid_out;
	assign SB_T0_NORTH_SB_IN_B17_enable = SB_T0_NORTH_SB_IN_B17_enable_value_O[0];
	assign SB_T0_NORTH_SB_IN_B17_ready_out = WIRE_SB_T0_NORTH_SB_IN_B17_ready_out;
	assign SB_T0_NORTH_SB_OUT_B17 = RMUX_T0_NORTH_B17_O;
	assign SB_T0_NORTH_SB_OUT_B17_enable = SB_T0_NORTH_SB_OUT_B17_enable_value_O[0];
	assign SB_T0_NORTH_SB_OUT_B17_valid_out = RMUX_T0_NORTH_B17_valid_out;
	assign SB_T0_SOUTH_SB_IN_B17_enable = SB_T0_SOUTH_SB_IN_B17_enable_value_O[0];
	assign SB_T0_SOUTH_SB_IN_B17_ready_out = WIRE_SB_T0_SOUTH_SB_IN_B17_ready_out;
	assign SB_T0_SOUTH_SB_OUT_B17 = RMUX_T0_SOUTH_B17_O;
	assign SB_T0_SOUTH_SB_OUT_B17_enable = SB_T0_SOUTH_SB_OUT_B17_enable_value_O[0];
	assign SB_T0_SOUTH_SB_OUT_B17_valid_out = RMUX_T0_SOUTH_B17_valid_out;
	assign SB_T0_WEST_SB_IN_B17_enable = SB_T0_WEST_SB_IN_B17_enable_value_O[0];
	assign SB_T0_WEST_SB_IN_B17_ready_out = WIRE_SB_T0_WEST_SB_IN_B17_ready_out;
	assign SB_T0_WEST_SB_OUT_B17 = RMUX_T0_WEST_B17_O;
	assign SB_T0_WEST_SB_OUT_B17_enable = SB_T0_WEST_SB_OUT_B17_enable_value_O[0];
	assign SB_T0_WEST_SB_OUT_B17_valid_out = RMUX_T0_WEST_B17_valid_out;
	assign SB_T1_EAST_SB_IN_B17_enable = SB_T1_EAST_SB_IN_B17_enable_value_O[0];
	assign SB_T1_EAST_SB_IN_B17_ready_out = WIRE_SB_T1_EAST_SB_IN_B17_ready_out;
	assign SB_T1_EAST_SB_OUT_B17 = RMUX_T1_EAST_B17_O;
	assign SB_T1_EAST_SB_OUT_B17_enable = SB_T1_EAST_SB_OUT_B17_enable_value_O[0];
	assign SB_T1_EAST_SB_OUT_B17_valid_out = RMUX_T1_EAST_B17_valid_out;
	assign SB_T1_NORTH_SB_IN_B17_enable = SB_T1_NORTH_SB_IN_B17_enable_value_O[0];
	assign SB_T1_NORTH_SB_IN_B17_ready_out = WIRE_SB_T1_NORTH_SB_IN_B17_ready_out;
	assign SB_T1_NORTH_SB_OUT_B17 = RMUX_T1_NORTH_B17_O;
	assign SB_T1_NORTH_SB_OUT_B17_enable = SB_T1_NORTH_SB_OUT_B17_enable_value_O[0];
	assign SB_T1_NORTH_SB_OUT_B17_valid_out = RMUX_T1_NORTH_B17_valid_out;
	assign SB_T1_SOUTH_SB_IN_B17_enable = SB_T1_SOUTH_SB_IN_B17_enable_value_O[0];
	assign SB_T1_SOUTH_SB_IN_B17_ready_out = WIRE_SB_T1_SOUTH_SB_IN_B17_ready_out;
	assign SB_T1_SOUTH_SB_OUT_B17 = RMUX_T1_SOUTH_B17_O;
	assign SB_T1_SOUTH_SB_OUT_B17_enable = SB_T1_SOUTH_SB_OUT_B17_enable_value_O[0];
	assign SB_T1_SOUTH_SB_OUT_B17_valid_out = RMUX_T1_SOUTH_B17_valid_out;
	assign SB_T1_WEST_SB_IN_B17_enable = SB_T1_WEST_SB_IN_B17_enable_value_O[0];
	assign SB_T1_WEST_SB_IN_B17_ready_out = WIRE_SB_T1_WEST_SB_IN_B17_ready_out;
	assign SB_T1_WEST_SB_OUT_B17 = RMUX_T1_WEST_B17_O;
	assign SB_T1_WEST_SB_OUT_B17_enable = SB_T1_WEST_SB_OUT_B17_enable_value_O[0];
	assign SB_T1_WEST_SB_OUT_B17_valid_out = RMUX_T1_WEST_B17_valid_out;
	assign SB_T2_EAST_SB_IN_B17_enable = SB_T2_EAST_SB_IN_B17_enable_value_O[0];
	assign SB_T2_EAST_SB_IN_B17_ready_out = WIRE_SB_T2_EAST_SB_IN_B17_ready_out;
	assign SB_T2_EAST_SB_OUT_B17 = RMUX_T2_EAST_B17_O;
	assign SB_T2_EAST_SB_OUT_B17_enable = SB_T2_EAST_SB_OUT_B17_enable_value_O[0];
	assign SB_T2_EAST_SB_OUT_B17_valid_out = RMUX_T2_EAST_B17_valid_out;
	assign SB_T2_NORTH_SB_IN_B17_enable = SB_T2_NORTH_SB_IN_B17_enable_value_O[0];
	assign SB_T2_NORTH_SB_IN_B17_ready_out = WIRE_SB_T2_NORTH_SB_IN_B17_ready_out;
	assign SB_T2_NORTH_SB_OUT_B17 = RMUX_T2_NORTH_B17_O;
	assign SB_T2_NORTH_SB_OUT_B17_enable = SB_T2_NORTH_SB_OUT_B17_enable_value_O[0];
	assign SB_T2_NORTH_SB_OUT_B17_valid_out = RMUX_T2_NORTH_B17_valid_out;
	assign SB_T2_SOUTH_SB_IN_B17_enable = SB_T2_SOUTH_SB_IN_B17_enable_value_O[0];
	assign SB_T2_SOUTH_SB_IN_B17_ready_out = WIRE_SB_T2_SOUTH_SB_IN_B17_ready_out;
	assign SB_T2_SOUTH_SB_OUT_B17 = RMUX_T2_SOUTH_B17_O;
	assign SB_T2_SOUTH_SB_OUT_B17_enable = SB_T2_SOUTH_SB_OUT_B17_enable_value_O[0];
	assign SB_T2_SOUTH_SB_OUT_B17_valid_out = RMUX_T2_SOUTH_B17_valid_out;
	assign SB_T2_WEST_SB_IN_B17_enable = SB_T2_WEST_SB_IN_B17_enable_value_O[0];
	assign SB_T2_WEST_SB_IN_B17_ready_out = WIRE_SB_T2_WEST_SB_IN_B17_ready_out;
	assign SB_T2_WEST_SB_OUT_B17 = RMUX_T2_WEST_B17_O;
	assign SB_T2_WEST_SB_OUT_B17_enable = SB_T2_WEST_SB_OUT_B17_enable_value_O[0];
	assign SB_T2_WEST_SB_OUT_B17_valid_out = RMUX_T2_WEST_B17_valid_out;
	assign SB_T3_EAST_SB_IN_B17_enable = SB_T3_EAST_SB_IN_B17_enable_value_O[0];
	assign SB_T3_EAST_SB_IN_B17_ready_out = WIRE_SB_T3_EAST_SB_IN_B17_ready_out;
	assign SB_T3_EAST_SB_OUT_B17 = RMUX_T3_EAST_B17_O;
	assign SB_T3_EAST_SB_OUT_B17_enable = SB_T3_EAST_SB_OUT_B17_enable_value_O[0];
	assign SB_T3_EAST_SB_OUT_B17_valid_out = RMUX_T3_EAST_B17_valid_out;
	assign SB_T3_NORTH_SB_IN_B17_enable = SB_T3_NORTH_SB_IN_B17_enable_value_O[0];
	assign SB_T3_NORTH_SB_IN_B17_ready_out = WIRE_SB_T3_NORTH_SB_IN_B17_ready_out;
	assign SB_T3_NORTH_SB_OUT_B17 = RMUX_T3_NORTH_B17_O;
	assign SB_T3_NORTH_SB_OUT_B17_enable = SB_T3_NORTH_SB_OUT_B17_enable_value_O[0];
	assign SB_T3_NORTH_SB_OUT_B17_valid_out = RMUX_T3_NORTH_B17_valid_out;
	assign SB_T3_SOUTH_SB_IN_B17_enable = SB_T3_SOUTH_SB_IN_B17_enable_value_O[0];
	assign SB_T3_SOUTH_SB_IN_B17_ready_out = WIRE_SB_T3_SOUTH_SB_IN_B17_ready_out;
	assign SB_T3_SOUTH_SB_OUT_B17 = RMUX_T3_SOUTH_B17_O;
	assign SB_T3_SOUTH_SB_OUT_B17_enable = SB_T3_SOUTH_SB_OUT_B17_enable_value_O[0];
	assign SB_T3_SOUTH_SB_OUT_B17_valid_out = RMUX_T3_SOUTH_B17_valid_out;
	assign SB_T3_WEST_SB_IN_B17_enable = SB_T3_WEST_SB_IN_B17_enable_value_O[0];
	assign SB_T3_WEST_SB_IN_B17_ready_out = WIRE_SB_T3_WEST_SB_IN_B17_ready_out;
	assign SB_T3_WEST_SB_OUT_B17 = RMUX_T3_WEST_B17_O;
	assign SB_T3_WEST_SB_OUT_B17_enable = SB_T3_WEST_SB_OUT_B17_enable_value_O[0];
	assign SB_T3_WEST_SB_OUT_B17_valid_out = RMUX_T3_WEST_B17_valid_out;
	assign SB_T4_EAST_SB_IN_B17_enable = SB_T4_EAST_SB_IN_B17_enable_value_O[0];
	assign SB_T4_EAST_SB_IN_B17_ready_out = WIRE_SB_T4_EAST_SB_IN_B17_ready_out;
	assign SB_T4_EAST_SB_OUT_B17 = RMUX_T4_EAST_B17_O;
	assign SB_T4_EAST_SB_OUT_B17_enable = SB_T4_EAST_SB_OUT_B17_enable_value_O[0];
	assign SB_T4_EAST_SB_OUT_B17_valid_out = RMUX_T4_EAST_B17_valid_out;
	assign SB_T4_NORTH_SB_IN_B17_enable = SB_T4_NORTH_SB_IN_B17_enable_value_O[0];
	assign SB_T4_NORTH_SB_IN_B17_ready_out = WIRE_SB_T4_NORTH_SB_IN_B17_ready_out;
	assign SB_T4_NORTH_SB_OUT_B17 = RMUX_T4_NORTH_B17_O;
	assign SB_T4_NORTH_SB_OUT_B17_enable = SB_T4_NORTH_SB_OUT_B17_enable_value_O[0];
	assign SB_T4_NORTH_SB_OUT_B17_valid_out = RMUX_T4_NORTH_B17_valid_out;
	assign SB_T4_SOUTH_SB_IN_B17_enable = SB_T4_SOUTH_SB_IN_B17_enable_value_O[0];
	assign SB_T4_SOUTH_SB_IN_B17_ready_out = WIRE_SB_T4_SOUTH_SB_IN_B17_ready_out;
	assign SB_T4_SOUTH_SB_OUT_B17 = RMUX_T4_SOUTH_B17_O;
	assign SB_T4_SOUTH_SB_OUT_B17_enable = SB_T4_SOUTH_SB_OUT_B17_enable_value_O[0];
	assign SB_T4_SOUTH_SB_OUT_B17_valid_out = RMUX_T4_SOUTH_B17_valid_out;
	assign SB_T4_WEST_SB_IN_B17_enable = SB_T4_WEST_SB_IN_B17_enable_value_O[0];
	assign SB_T4_WEST_SB_IN_B17_ready_out = WIRE_SB_T4_WEST_SB_IN_B17_ready_out;
	assign SB_T4_WEST_SB_OUT_B17 = RMUX_T4_WEST_B17_O;
	assign SB_T4_WEST_SB_OUT_B17_enable = SB_T4_WEST_SB_OUT_B17_enable_value_O[0];
	assign SB_T4_WEST_SB_OUT_B17_valid_out = RMUX_T4_WEST_B17_valid_out;
	assign read_config_data = mux_aoi_6_32_inst0_O;
endmodule
module SB_ID0_5TRACKS_B17_MemCore (
	MEM_input_width_17_num_0_enable,
	MEM_input_width_17_num_0_out_sel,
	MEM_input_width_17_num_0_ready,
	MEM_input_width_17_num_1_enable,
	MEM_input_width_17_num_1_out_sel,
	MEM_input_width_17_num_1_ready,
	MEM_input_width_17_num_2_enable,
	MEM_input_width_17_num_2_out_sel,
	MEM_input_width_17_num_2_ready,
	MEM_input_width_17_num_3_enable,
	MEM_input_width_17_num_3_out_sel,
	MEM_input_width_17_num_3_ready,
	MEM_output_width_17_num_0,
	MEM_output_width_17_num_0_ready_out,
	MEM_output_width_17_num_0_valid,
	MEM_output_width_17_num_1,
	MEM_output_width_17_num_1_ready_out,
	MEM_output_width_17_num_1_valid,
	MEM_output_width_17_num_2,
	MEM_output_width_17_num_2_ready_out,
	MEM_output_width_17_num_2_valid,
	SB_T0_EAST_SB_IN_B17,
	SB_T0_EAST_SB_IN_B17_enable,
	SB_T0_EAST_SB_IN_B17_ready_out,
	SB_T0_EAST_SB_IN_B17_valid_in,
	SB_T0_EAST_SB_OUT_B17,
	SB_T0_EAST_SB_OUT_B17_enable,
	SB_T0_EAST_SB_OUT_B17_ready_in,
	SB_T0_EAST_SB_OUT_B17_valid_out,
	SB_T0_NORTH_SB_IN_B17,
	SB_T0_NORTH_SB_IN_B17_enable,
	SB_T0_NORTH_SB_IN_B17_ready_out,
	SB_T0_NORTH_SB_IN_B17_valid_in,
	SB_T0_NORTH_SB_OUT_B17,
	SB_T0_NORTH_SB_OUT_B17_enable,
	SB_T0_NORTH_SB_OUT_B17_ready_in,
	SB_T0_NORTH_SB_OUT_B17_valid_out,
	SB_T0_SOUTH_SB_IN_B17,
	SB_T0_SOUTH_SB_IN_B17_enable,
	SB_T0_SOUTH_SB_IN_B17_ready_out,
	SB_T0_SOUTH_SB_IN_B17_valid_in,
	SB_T0_SOUTH_SB_OUT_B17,
	SB_T0_SOUTH_SB_OUT_B17_enable,
	SB_T0_SOUTH_SB_OUT_B17_ready_in,
	SB_T0_SOUTH_SB_OUT_B17_valid_out,
	SB_T0_WEST_SB_IN_B17,
	SB_T0_WEST_SB_IN_B17_enable,
	SB_T0_WEST_SB_IN_B17_ready_out,
	SB_T0_WEST_SB_IN_B17_valid_in,
	SB_T0_WEST_SB_OUT_B17,
	SB_T0_WEST_SB_OUT_B17_enable,
	SB_T0_WEST_SB_OUT_B17_ready_in,
	SB_T0_WEST_SB_OUT_B17_valid_out,
	SB_T1_EAST_SB_IN_B17,
	SB_T1_EAST_SB_IN_B17_enable,
	SB_T1_EAST_SB_IN_B17_ready_out,
	SB_T1_EAST_SB_IN_B17_valid_in,
	SB_T1_EAST_SB_OUT_B17,
	SB_T1_EAST_SB_OUT_B17_enable,
	SB_T1_EAST_SB_OUT_B17_ready_in,
	SB_T1_EAST_SB_OUT_B17_valid_out,
	SB_T1_NORTH_SB_IN_B17,
	SB_T1_NORTH_SB_IN_B17_enable,
	SB_T1_NORTH_SB_IN_B17_ready_out,
	SB_T1_NORTH_SB_IN_B17_valid_in,
	SB_T1_NORTH_SB_OUT_B17,
	SB_T1_NORTH_SB_OUT_B17_enable,
	SB_T1_NORTH_SB_OUT_B17_ready_in,
	SB_T1_NORTH_SB_OUT_B17_valid_out,
	SB_T1_SOUTH_SB_IN_B17,
	SB_T1_SOUTH_SB_IN_B17_enable,
	SB_T1_SOUTH_SB_IN_B17_ready_out,
	SB_T1_SOUTH_SB_IN_B17_valid_in,
	SB_T1_SOUTH_SB_OUT_B17,
	SB_T1_SOUTH_SB_OUT_B17_enable,
	SB_T1_SOUTH_SB_OUT_B17_ready_in,
	SB_T1_SOUTH_SB_OUT_B17_valid_out,
	SB_T1_WEST_SB_IN_B17,
	SB_T1_WEST_SB_IN_B17_enable,
	SB_T1_WEST_SB_IN_B17_ready_out,
	SB_T1_WEST_SB_IN_B17_valid_in,
	SB_T1_WEST_SB_OUT_B17,
	SB_T1_WEST_SB_OUT_B17_enable,
	SB_T1_WEST_SB_OUT_B17_ready_in,
	SB_T1_WEST_SB_OUT_B17_valid_out,
	SB_T2_EAST_SB_IN_B17,
	SB_T2_EAST_SB_IN_B17_enable,
	SB_T2_EAST_SB_IN_B17_ready_out,
	SB_T2_EAST_SB_IN_B17_valid_in,
	SB_T2_EAST_SB_OUT_B17,
	SB_T2_EAST_SB_OUT_B17_enable,
	SB_T2_EAST_SB_OUT_B17_ready_in,
	SB_T2_EAST_SB_OUT_B17_valid_out,
	SB_T2_NORTH_SB_IN_B17,
	SB_T2_NORTH_SB_IN_B17_enable,
	SB_T2_NORTH_SB_IN_B17_ready_out,
	SB_T2_NORTH_SB_IN_B17_valid_in,
	SB_T2_NORTH_SB_OUT_B17,
	SB_T2_NORTH_SB_OUT_B17_enable,
	SB_T2_NORTH_SB_OUT_B17_ready_in,
	SB_T2_NORTH_SB_OUT_B17_valid_out,
	SB_T2_SOUTH_SB_IN_B17,
	SB_T2_SOUTH_SB_IN_B17_enable,
	SB_T2_SOUTH_SB_IN_B17_ready_out,
	SB_T2_SOUTH_SB_IN_B17_valid_in,
	SB_T2_SOUTH_SB_OUT_B17,
	SB_T2_SOUTH_SB_OUT_B17_enable,
	SB_T2_SOUTH_SB_OUT_B17_ready_in,
	SB_T2_SOUTH_SB_OUT_B17_valid_out,
	SB_T2_WEST_SB_IN_B17,
	SB_T2_WEST_SB_IN_B17_enable,
	SB_T2_WEST_SB_IN_B17_ready_out,
	SB_T2_WEST_SB_IN_B17_valid_in,
	SB_T2_WEST_SB_OUT_B17,
	SB_T2_WEST_SB_OUT_B17_enable,
	SB_T2_WEST_SB_OUT_B17_ready_in,
	SB_T2_WEST_SB_OUT_B17_valid_out,
	SB_T3_EAST_SB_IN_B17,
	SB_T3_EAST_SB_IN_B17_enable,
	SB_T3_EAST_SB_IN_B17_ready_out,
	SB_T3_EAST_SB_IN_B17_valid_in,
	SB_T3_EAST_SB_OUT_B17,
	SB_T3_EAST_SB_OUT_B17_enable,
	SB_T3_EAST_SB_OUT_B17_ready_in,
	SB_T3_EAST_SB_OUT_B17_valid_out,
	SB_T3_NORTH_SB_IN_B17,
	SB_T3_NORTH_SB_IN_B17_enable,
	SB_T3_NORTH_SB_IN_B17_ready_out,
	SB_T3_NORTH_SB_IN_B17_valid_in,
	SB_T3_NORTH_SB_OUT_B17,
	SB_T3_NORTH_SB_OUT_B17_enable,
	SB_T3_NORTH_SB_OUT_B17_ready_in,
	SB_T3_NORTH_SB_OUT_B17_valid_out,
	SB_T3_SOUTH_SB_IN_B17,
	SB_T3_SOUTH_SB_IN_B17_enable,
	SB_T3_SOUTH_SB_IN_B17_ready_out,
	SB_T3_SOUTH_SB_IN_B17_valid_in,
	SB_T3_SOUTH_SB_OUT_B17,
	SB_T3_SOUTH_SB_OUT_B17_enable,
	SB_T3_SOUTH_SB_OUT_B17_ready_in,
	SB_T3_SOUTH_SB_OUT_B17_valid_out,
	SB_T3_WEST_SB_IN_B17,
	SB_T3_WEST_SB_IN_B17_enable,
	SB_T3_WEST_SB_IN_B17_ready_out,
	SB_T3_WEST_SB_IN_B17_valid_in,
	SB_T3_WEST_SB_OUT_B17,
	SB_T3_WEST_SB_OUT_B17_enable,
	SB_T3_WEST_SB_OUT_B17_ready_in,
	SB_T3_WEST_SB_OUT_B17_valid_out,
	SB_T4_EAST_SB_IN_B17,
	SB_T4_EAST_SB_IN_B17_enable,
	SB_T4_EAST_SB_IN_B17_ready_out,
	SB_T4_EAST_SB_IN_B17_valid_in,
	SB_T4_EAST_SB_OUT_B17,
	SB_T4_EAST_SB_OUT_B17_enable,
	SB_T4_EAST_SB_OUT_B17_ready_in,
	SB_T4_EAST_SB_OUT_B17_valid_out,
	SB_T4_NORTH_SB_IN_B17,
	SB_T4_NORTH_SB_IN_B17_enable,
	SB_T4_NORTH_SB_IN_B17_ready_out,
	SB_T4_NORTH_SB_IN_B17_valid_in,
	SB_T4_NORTH_SB_OUT_B17,
	SB_T4_NORTH_SB_OUT_B17_enable,
	SB_T4_NORTH_SB_OUT_B17_ready_in,
	SB_T4_NORTH_SB_OUT_B17_valid_out,
	SB_T4_SOUTH_SB_IN_B17,
	SB_T4_SOUTH_SB_IN_B17_enable,
	SB_T4_SOUTH_SB_IN_B17_ready_out,
	SB_T4_SOUTH_SB_IN_B17_valid_in,
	SB_T4_SOUTH_SB_OUT_B17,
	SB_T4_SOUTH_SB_OUT_B17_enable,
	SB_T4_SOUTH_SB_OUT_B17_ready_in,
	SB_T4_SOUTH_SB_OUT_B17_valid_out,
	SB_T4_WEST_SB_IN_B17,
	SB_T4_WEST_SB_IN_B17_enable,
	SB_T4_WEST_SB_IN_B17_ready_out,
	SB_T4_WEST_SB_IN_B17_valid_in,
	SB_T4_WEST_SB_OUT_B17,
	SB_T4_WEST_SB_OUT_B17_enable,
	SB_T4_WEST_SB_OUT_B17_ready_in,
	SB_T4_WEST_SB_OUT_B17_valid_out,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	read_config_data,
	reset,
	stall
);
	input [0:0] MEM_input_width_17_num_0_enable;
	input [31:0] MEM_input_width_17_num_0_out_sel;
	input MEM_input_width_17_num_0_ready;
	input [0:0] MEM_input_width_17_num_1_enable;
	input [31:0] MEM_input_width_17_num_1_out_sel;
	input MEM_input_width_17_num_1_ready;
	input [0:0] MEM_input_width_17_num_2_enable;
	input [31:0] MEM_input_width_17_num_2_out_sel;
	input MEM_input_width_17_num_2_ready;
	input [0:0] MEM_input_width_17_num_3_enable;
	input [31:0] MEM_input_width_17_num_3_out_sel;
	input MEM_input_width_17_num_3_ready;
	input [16:0] MEM_output_width_17_num_0;
	output wire MEM_output_width_17_num_0_ready_out;
	input MEM_output_width_17_num_0_valid;
	input [16:0] MEM_output_width_17_num_1;
	output wire MEM_output_width_17_num_1_ready_out;
	input MEM_output_width_17_num_1_valid;
	input [16:0] MEM_output_width_17_num_2;
	output wire MEM_output_width_17_num_2_ready_out;
	input MEM_output_width_17_num_2_valid;
	input [16:0] SB_T0_EAST_SB_IN_B17;
	output wire SB_T0_EAST_SB_IN_B17_enable;
	output wire SB_T0_EAST_SB_IN_B17_ready_out;
	input SB_T0_EAST_SB_IN_B17_valid_in;
	output wire [16:0] SB_T0_EAST_SB_OUT_B17;
	output wire SB_T0_EAST_SB_OUT_B17_enable;
	input SB_T0_EAST_SB_OUT_B17_ready_in;
	output wire SB_T0_EAST_SB_OUT_B17_valid_out;
	input [16:0] SB_T0_NORTH_SB_IN_B17;
	output wire SB_T0_NORTH_SB_IN_B17_enable;
	output wire SB_T0_NORTH_SB_IN_B17_ready_out;
	input SB_T0_NORTH_SB_IN_B17_valid_in;
	output wire [16:0] SB_T0_NORTH_SB_OUT_B17;
	output wire SB_T0_NORTH_SB_OUT_B17_enable;
	input SB_T0_NORTH_SB_OUT_B17_ready_in;
	output wire SB_T0_NORTH_SB_OUT_B17_valid_out;
	input [16:0] SB_T0_SOUTH_SB_IN_B17;
	output wire SB_T0_SOUTH_SB_IN_B17_enable;
	output wire SB_T0_SOUTH_SB_IN_B17_ready_out;
	input SB_T0_SOUTH_SB_IN_B17_valid_in;
	output wire [16:0] SB_T0_SOUTH_SB_OUT_B17;
	output wire SB_T0_SOUTH_SB_OUT_B17_enable;
	input SB_T0_SOUTH_SB_OUT_B17_ready_in;
	output wire SB_T0_SOUTH_SB_OUT_B17_valid_out;
	input [16:0] SB_T0_WEST_SB_IN_B17;
	output wire SB_T0_WEST_SB_IN_B17_enable;
	output wire SB_T0_WEST_SB_IN_B17_ready_out;
	input SB_T0_WEST_SB_IN_B17_valid_in;
	output wire [16:0] SB_T0_WEST_SB_OUT_B17;
	output wire SB_T0_WEST_SB_OUT_B17_enable;
	input SB_T0_WEST_SB_OUT_B17_ready_in;
	output wire SB_T0_WEST_SB_OUT_B17_valid_out;
	input [16:0] SB_T1_EAST_SB_IN_B17;
	output wire SB_T1_EAST_SB_IN_B17_enable;
	output wire SB_T1_EAST_SB_IN_B17_ready_out;
	input SB_T1_EAST_SB_IN_B17_valid_in;
	output wire [16:0] SB_T1_EAST_SB_OUT_B17;
	output wire SB_T1_EAST_SB_OUT_B17_enable;
	input SB_T1_EAST_SB_OUT_B17_ready_in;
	output wire SB_T1_EAST_SB_OUT_B17_valid_out;
	input [16:0] SB_T1_NORTH_SB_IN_B17;
	output wire SB_T1_NORTH_SB_IN_B17_enable;
	output wire SB_T1_NORTH_SB_IN_B17_ready_out;
	input SB_T1_NORTH_SB_IN_B17_valid_in;
	output wire [16:0] SB_T1_NORTH_SB_OUT_B17;
	output wire SB_T1_NORTH_SB_OUT_B17_enable;
	input SB_T1_NORTH_SB_OUT_B17_ready_in;
	output wire SB_T1_NORTH_SB_OUT_B17_valid_out;
	input [16:0] SB_T1_SOUTH_SB_IN_B17;
	output wire SB_T1_SOUTH_SB_IN_B17_enable;
	output wire SB_T1_SOUTH_SB_IN_B17_ready_out;
	input SB_T1_SOUTH_SB_IN_B17_valid_in;
	output wire [16:0] SB_T1_SOUTH_SB_OUT_B17;
	output wire SB_T1_SOUTH_SB_OUT_B17_enable;
	input SB_T1_SOUTH_SB_OUT_B17_ready_in;
	output wire SB_T1_SOUTH_SB_OUT_B17_valid_out;
	input [16:0] SB_T1_WEST_SB_IN_B17;
	output wire SB_T1_WEST_SB_IN_B17_enable;
	output wire SB_T1_WEST_SB_IN_B17_ready_out;
	input SB_T1_WEST_SB_IN_B17_valid_in;
	output wire [16:0] SB_T1_WEST_SB_OUT_B17;
	output wire SB_T1_WEST_SB_OUT_B17_enable;
	input SB_T1_WEST_SB_OUT_B17_ready_in;
	output wire SB_T1_WEST_SB_OUT_B17_valid_out;
	input [16:0] SB_T2_EAST_SB_IN_B17;
	output wire SB_T2_EAST_SB_IN_B17_enable;
	output wire SB_T2_EAST_SB_IN_B17_ready_out;
	input SB_T2_EAST_SB_IN_B17_valid_in;
	output wire [16:0] SB_T2_EAST_SB_OUT_B17;
	output wire SB_T2_EAST_SB_OUT_B17_enable;
	input SB_T2_EAST_SB_OUT_B17_ready_in;
	output wire SB_T2_EAST_SB_OUT_B17_valid_out;
	input [16:0] SB_T2_NORTH_SB_IN_B17;
	output wire SB_T2_NORTH_SB_IN_B17_enable;
	output wire SB_T2_NORTH_SB_IN_B17_ready_out;
	input SB_T2_NORTH_SB_IN_B17_valid_in;
	output wire [16:0] SB_T2_NORTH_SB_OUT_B17;
	output wire SB_T2_NORTH_SB_OUT_B17_enable;
	input SB_T2_NORTH_SB_OUT_B17_ready_in;
	output wire SB_T2_NORTH_SB_OUT_B17_valid_out;
	input [16:0] SB_T2_SOUTH_SB_IN_B17;
	output wire SB_T2_SOUTH_SB_IN_B17_enable;
	output wire SB_T2_SOUTH_SB_IN_B17_ready_out;
	input SB_T2_SOUTH_SB_IN_B17_valid_in;
	output wire [16:0] SB_T2_SOUTH_SB_OUT_B17;
	output wire SB_T2_SOUTH_SB_OUT_B17_enable;
	input SB_T2_SOUTH_SB_OUT_B17_ready_in;
	output wire SB_T2_SOUTH_SB_OUT_B17_valid_out;
	input [16:0] SB_T2_WEST_SB_IN_B17;
	output wire SB_T2_WEST_SB_IN_B17_enable;
	output wire SB_T2_WEST_SB_IN_B17_ready_out;
	input SB_T2_WEST_SB_IN_B17_valid_in;
	output wire [16:0] SB_T2_WEST_SB_OUT_B17;
	output wire SB_T2_WEST_SB_OUT_B17_enable;
	input SB_T2_WEST_SB_OUT_B17_ready_in;
	output wire SB_T2_WEST_SB_OUT_B17_valid_out;
	input [16:0] SB_T3_EAST_SB_IN_B17;
	output wire SB_T3_EAST_SB_IN_B17_enable;
	output wire SB_T3_EAST_SB_IN_B17_ready_out;
	input SB_T3_EAST_SB_IN_B17_valid_in;
	output wire [16:0] SB_T3_EAST_SB_OUT_B17;
	output wire SB_T3_EAST_SB_OUT_B17_enable;
	input SB_T3_EAST_SB_OUT_B17_ready_in;
	output wire SB_T3_EAST_SB_OUT_B17_valid_out;
	input [16:0] SB_T3_NORTH_SB_IN_B17;
	output wire SB_T3_NORTH_SB_IN_B17_enable;
	output wire SB_T3_NORTH_SB_IN_B17_ready_out;
	input SB_T3_NORTH_SB_IN_B17_valid_in;
	output wire [16:0] SB_T3_NORTH_SB_OUT_B17;
	output wire SB_T3_NORTH_SB_OUT_B17_enable;
	input SB_T3_NORTH_SB_OUT_B17_ready_in;
	output wire SB_T3_NORTH_SB_OUT_B17_valid_out;
	input [16:0] SB_T3_SOUTH_SB_IN_B17;
	output wire SB_T3_SOUTH_SB_IN_B17_enable;
	output wire SB_T3_SOUTH_SB_IN_B17_ready_out;
	input SB_T3_SOUTH_SB_IN_B17_valid_in;
	output wire [16:0] SB_T3_SOUTH_SB_OUT_B17;
	output wire SB_T3_SOUTH_SB_OUT_B17_enable;
	input SB_T3_SOUTH_SB_OUT_B17_ready_in;
	output wire SB_T3_SOUTH_SB_OUT_B17_valid_out;
	input [16:0] SB_T3_WEST_SB_IN_B17;
	output wire SB_T3_WEST_SB_IN_B17_enable;
	output wire SB_T3_WEST_SB_IN_B17_ready_out;
	input SB_T3_WEST_SB_IN_B17_valid_in;
	output wire [16:0] SB_T3_WEST_SB_OUT_B17;
	output wire SB_T3_WEST_SB_OUT_B17_enable;
	input SB_T3_WEST_SB_OUT_B17_ready_in;
	output wire SB_T3_WEST_SB_OUT_B17_valid_out;
	input [16:0] SB_T4_EAST_SB_IN_B17;
	output wire SB_T4_EAST_SB_IN_B17_enable;
	output wire SB_T4_EAST_SB_IN_B17_ready_out;
	input SB_T4_EAST_SB_IN_B17_valid_in;
	output wire [16:0] SB_T4_EAST_SB_OUT_B17;
	output wire SB_T4_EAST_SB_OUT_B17_enable;
	input SB_T4_EAST_SB_OUT_B17_ready_in;
	output wire SB_T4_EAST_SB_OUT_B17_valid_out;
	input [16:0] SB_T4_NORTH_SB_IN_B17;
	output wire SB_T4_NORTH_SB_IN_B17_enable;
	output wire SB_T4_NORTH_SB_IN_B17_ready_out;
	input SB_T4_NORTH_SB_IN_B17_valid_in;
	output wire [16:0] SB_T4_NORTH_SB_OUT_B17;
	output wire SB_T4_NORTH_SB_OUT_B17_enable;
	input SB_T4_NORTH_SB_OUT_B17_ready_in;
	output wire SB_T4_NORTH_SB_OUT_B17_valid_out;
	input [16:0] SB_T4_SOUTH_SB_IN_B17;
	output wire SB_T4_SOUTH_SB_IN_B17_enable;
	output wire SB_T4_SOUTH_SB_IN_B17_ready_out;
	input SB_T4_SOUTH_SB_IN_B17_valid_in;
	output wire [16:0] SB_T4_SOUTH_SB_OUT_B17;
	output wire SB_T4_SOUTH_SB_OUT_B17_enable;
	input SB_T4_SOUTH_SB_OUT_B17_ready_in;
	output wire SB_T4_SOUTH_SB_OUT_B17_valid_out;
	input [16:0] SB_T4_WEST_SB_IN_B17;
	output wire SB_T4_WEST_SB_IN_B17_enable;
	output wire SB_T4_WEST_SB_IN_B17_ready_out;
	input SB_T4_WEST_SB_IN_B17_valid_in;
	output wire [16:0] SB_T4_WEST_SB_OUT_B17;
	output wire SB_T4_WEST_SB_OUT_B17_enable;
	input SB_T4_WEST_SB_OUT_B17_ready_in;
	output wire SB_T4_WEST_SB_OUT_B17_valid_out;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output wire [31:0] read_config_data;
	input reset;
	input [0:0] stall;
	wire [0:0] CB_MEM_output_width_17_num_0_fan_in_O;
	wire [0:0] CB_MEM_output_width_17_num_1_fan_in_O;
	wire [0:0] CB_MEM_output_width_17_num_2_fan_in_O;
	wire [0:0] Invert1_inst0_out;
	wire [16:0] MUX_SB_T0_EAST_SB_OUT_B17_O;
	wire MUX_SB_T0_EAST_SB_OUT_B17_ready_out;
	wire MUX_SB_T0_EAST_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T0_EAST_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T0_NORTH_SB_OUT_B17_O;
	wire MUX_SB_T0_NORTH_SB_OUT_B17_ready_out;
	wire MUX_SB_T0_NORTH_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T0_NORTH_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T0_SOUTH_SB_OUT_B17_O;
	wire MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out;
	wire MUX_SB_T0_SOUTH_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T0_WEST_SB_OUT_B17_O;
	wire MUX_SB_T0_WEST_SB_OUT_B17_ready_out;
	wire MUX_SB_T0_WEST_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T0_WEST_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T1_EAST_SB_OUT_B17_O;
	wire MUX_SB_T1_EAST_SB_OUT_B17_ready_out;
	wire MUX_SB_T1_EAST_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T1_EAST_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T1_NORTH_SB_OUT_B17_O;
	wire MUX_SB_T1_NORTH_SB_OUT_B17_ready_out;
	wire MUX_SB_T1_NORTH_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T1_NORTH_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T1_SOUTH_SB_OUT_B17_O;
	wire MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out;
	wire MUX_SB_T1_SOUTH_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T1_WEST_SB_OUT_B17_O;
	wire MUX_SB_T1_WEST_SB_OUT_B17_ready_out;
	wire MUX_SB_T1_WEST_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T1_WEST_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T2_EAST_SB_OUT_B17_O;
	wire MUX_SB_T2_EAST_SB_OUT_B17_ready_out;
	wire MUX_SB_T2_EAST_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T2_EAST_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T2_NORTH_SB_OUT_B17_O;
	wire MUX_SB_T2_NORTH_SB_OUT_B17_ready_out;
	wire MUX_SB_T2_NORTH_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T2_NORTH_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T2_SOUTH_SB_OUT_B17_O;
	wire MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out;
	wire MUX_SB_T2_SOUTH_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T2_WEST_SB_OUT_B17_O;
	wire MUX_SB_T2_WEST_SB_OUT_B17_ready_out;
	wire MUX_SB_T2_WEST_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T2_WEST_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T3_EAST_SB_OUT_B17_O;
	wire MUX_SB_T3_EAST_SB_OUT_B17_ready_out;
	wire MUX_SB_T3_EAST_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T3_EAST_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T3_NORTH_SB_OUT_B17_O;
	wire MUX_SB_T3_NORTH_SB_OUT_B17_ready_out;
	wire MUX_SB_T3_NORTH_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T3_NORTH_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T3_SOUTH_SB_OUT_B17_O;
	wire MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out;
	wire MUX_SB_T3_SOUTH_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T3_WEST_SB_OUT_B17_O;
	wire MUX_SB_T3_WEST_SB_OUT_B17_ready_out;
	wire MUX_SB_T3_WEST_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T3_WEST_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T4_EAST_SB_OUT_B17_O;
	wire MUX_SB_T4_EAST_SB_OUT_B17_ready_out;
	wire MUX_SB_T4_EAST_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T4_EAST_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T4_NORTH_SB_OUT_B17_O;
	wire MUX_SB_T4_NORTH_SB_OUT_B17_ready_out;
	wire MUX_SB_T4_NORTH_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T4_NORTH_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T4_SOUTH_SB_OUT_B17_O;
	wire MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out;
	wire MUX_SB_T4_SOUTH_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel;
	wire [16:0] MUX_SB_T4_WEST_SB_OUT_B17_O;
	wire MUX_SB_T4_WEST_SB_OUT_B17_ready_out;
	wire MUX_SB_T4_WEST_SB_OUT_B17_valid_out;
	wire [7:0] MUX_SB_T4_WEST_SB_OUT_B17_out_sel;
	wire [0:0] REG_T0_EAST_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T0_EAST_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T0_EAST_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T0_EAST_B17_end_value_O;
	wire [0:0] REG_T0_EAST_B17_fifo_value_O;
	wire [0:0] REG_T0_EAST_B17_start_value_O;
	wire [0:0] REG_T0_NORTH_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T0_NORTH_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T0_NORTH_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T0_NORTH_B17_end_value_O;
	wire [0:0] REG_T0_NORTH_B17_fifo_value_O;
	wire [0:0] REG_T0_NORTH_B17_start_value_O;
	wire [0:0] REG_T0_SOUTH_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T0_SOUTH_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T0_SOUTH_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T0_SOUTH_B17_end_value_O;
	wire [0:0] REG_T0_SOUTH_B17_fifo_value_O;
	wire [0:0] REG_T0_SOUTH_B17_start_value_O;
	wire [0:0] REG_T0_WEST_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T0_WEST_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T0_WEST_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T0_WEST_B17_end_value_O;
	wire [0:0] REG_T0_WEST_B17_fifo_value_O;
	wire [0:0] REG_T0_WEST_B17_start_value_O;
	wire [0:0] REG_T1_EAST_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T1_EAST_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T1_EAST_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T1_EAST_B17_end_value_O;
	wire [0:0] REG_T1_EAST_B17_fifo_value_O;
	wire [0:0] REG_T1_EAST_B17_start_value_O;
	wire [0:0] REG_T1_NORTH_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T1_NORTH_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T1_NORTH_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T1_NORTH_B17_end_value_O;
	wire [0:0] REG_T1_NORTH_B17_fifo_value_O;
	wire [0:0] REG_T1_NORTH_B17_start_value_O;
	wire [0:0] REG_T1_SOUTH_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T1_SOUTH_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T1_SOUTH_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T1_SOUTH_B17_end_value_O;
	wire [0:0] REG_T1_SOUTH_B17_fifo_value_O;
	wire [0:0] REG_T1_SOUTH_B17_start_value_O;
	wire [0:0] REG_T1_WEST_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T1_WEST_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T1_WEST_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T1_WEST_B17_end_value_O;
	wire [0:0] REG_T1_WEST_B17_fifo_value_O;
	wire [0:0] REG_T1_WEST_B17_start_value_O;
	wire [0:0] REG_T2_EAST_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T2_EAST_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T2_EAST_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T2_EAST_B17_end_value_O;
	wire [0:0] REG_T2_EAST_B17_fifo_value_O;
	wire [0:0] REG_T2_EAST_B17_start_value_O;
	wire [0:0] REG_T2_NORTH_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T2_NORTH_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T2_NORTH_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T2_NORTH_B17_end_value_O;
	wire [0:0] REG_T2_NORTH_B17_fifo_value_O;
	wire [0:0] REG_T2_NORTH_B17_start_value_O;
	wire [0:0] REG_T2_SOUTH_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T2_SOUTH_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T2_SOUTH_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T2_SOUTH_B17_end_value_O;
	wire [0:0] REG_T2_SOUTH_B17_fifo_value_O;
	wire [0:0] REG_T2_SOUTH_B17_start_value_O;
	wire [0:0] REG_T2_WEST_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T2_WEST_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T2_WEST_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T2_WEST_B17_end_value_O;
	wire [0:0] REG_T2_WEST_B17_fifo_value_O;
	wire [0:0] REG_T2_WEST_B17_start_value_O;
	wire [0:0] REG_T3_EAST_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T3_EAST_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T3_EAST_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T3_EAST_B17_end_value_O;
	wire [0:0] REG_T3_EAST_B17_fifo_value_O;
	wire [0:0] REG_T3_EAST_B17_start_value_O;
	wire [0:0] REG_T3_NORTH_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T3_NORTH_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T3_NORTH_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T3_NORTH_B17_end_value_O;
	wire [0:0] REG_T3_NORTH_B17_fifo_value_O;
	wire [0:0] REG_T3_NORTH_B17_start_value_O;
	wire [0:0] REG_T3_SOUTH_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T3_SOUTH_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T3_SOUTH_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T3_SOUTH_B17_end_value_O;
	wire [0:0] REG_T3_SOUTH_B17_fifo_value_O;
	wire [0:0] REG_T3_SOUTH_B17_start_value_O;
	wire [0:0] REG_T3_WEST_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T3_WEST_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T3_WEST_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T3_WEST_B17_end_value_O;
	wire [0:0] REG_T3_WEST_B17_fifo_value_O;
	wire [0:0] REG_T3_WEST_B17_start_value_O;
	wire [0:0] REG_T4_EAST_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T4_EAST_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T4_EAST_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T4_EAST_B17_end_value_O;
	wire [0:0] REG_T4_EAST_B17_fifo_value_O;
	wire [0:0] REG_T4_EAST_B17_start_value_O;
	wire [0:0] REG_T4_NORTH_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T4_NORTH_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T4_NORTH_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T4_NORTH_B17_end_value_O;
	wire [0:0] REG_T4_NORTH_B17_fifo_value_O;
	wire [0:0] REG_T4_NORTH_B17_start_value_O;
	wire [0:0] REG_T4_SOUTH_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T4_SOUTH_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T4_SOUTH_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T4_SOUTH_B17_end_value_O;
	wire [0:0] REG_T4_SOUTH_B17_fifo_value_O;
	wire [0:0] REG_T4_SOUTH_B17_start_value_O;
	wire [0:0] REG_T4_WEST_B17$SplitFifo_17_inst0_ready0;
	wire [16:0] REG_T4_WEST_B17$SplitFifo_17_inst0_data_out;
	wire [0:0] REG_T4_WEST_B17$SplitFifo_17_inst0_valid1;
	wire [0:0] REG_T4_WEST_B17_end_value_O;
	wire [0:0] REG_T4_WEST_B17_fifo_value_O;
	wire [0:0] REG_T4_WEST_B17_start_value_O;
	wire [16:0] RMUX_T0_EAST_B17_O;
	wire RMUX_T0_EAST_B17_ready_out;
	wire RMUX_T0_EAST_B17_valid_out;
	wire [1:0] RMUX_T0_EAST_B17_out_sel;
	wire [0:0] RMUX_T0_EAST_B17_sel_value_O;
	wire [16:0] RMUX_T0_NORTH_B17_O;
	wire RMUX_T0_NORTH_B17_ready_out;
	wire RMUX_T0_NORTH_B17_valid_out;
	wire [1:0] RMUX_T0_NORTH_B17_out_sel;
	wire [0:0] RMUX_T0_NORTH_B17_sel_value_O;
	wire [16:0] RMUX_T0_SOUTH_B17_O;
	wire RMUX_T0_SOUTH_B17_ready_out;
	wire RMUX_T0_SOUTH_B17_valid_out;
	wire [1:0] RMUX_T0_SOUTH_B17_out_sel;
	wire [0:0] RMUX_T0_SOUTH_B17_sel_value_O;
	wire [16:0] RMUX_T0_WEST_B17_O;
	wire RMUX_T0_WEST_B17_ready_out;
	wire RMUX_T0_WEST_B17_valid_out;
	wire [1:0] RMUX_T0_WEST_B17_out_sel;
	wire [0:0] RMUX_T0_WEST_B17_sel_value_O;
	wire [16:0] RMUX_T1_EAST_B17_O;
	wire RMUX_T1_EAST_B17_ready_out;
	wire RMUX_T1_EAST_B17_valid_out;
	wire [1:0] RMUX_T1_EAST_B17_out_sel;
	wire [0:0] RMUX_T1_EAST_B17_sel_value_O;
	wire [16:0] RMUX_T1_NORTH_B17_O;
	wire RMUX_T1_NORTH_B17_ready_out;
	wire RMUX_T1_NORTH_B17_valid_out;
	wire [1:0] RMUX_T1_NORTH_B17_out_sel;
	wire [0:0] RMUX_T1_NORTH_B17_sel_value_O;
	wire [16:0] RMUX_T1_SOUTH_B17_O;
	wire RMUX_T1_SOUTH_B17_ready_out;
	wire RMUX_T1_SOUTH_B17_valid_out;
	wire [1:0] RMUX_T1_SOUTH_B17_out_sel;
	wire [0:0] RMUX_T1_SOUTH_B17_sel_value_O;
	wire [16:0] RMUX_T1_WEST_B17_O;
	wire RMUX_T1_WEST_B17_ready_out;
	wire RMUX_T1_WEST_B17_valid_out;
	wire [1:0] RMUX_T1_WEST_B17_out_sel;
	wire [0:0] RMUX_T1_WEST_B17_sel_value_O;
	wire [16:0] RMUX_T2_EAST_B17_O;
	wire RMUX_T2_EAST_B17_ready_out;
	wire RMUX_T2_EAST_B17_valid_out;
	wire [1:0] RMUX_T2_EAST_B17_out_sel;
	wire [0:0] RMUX_T2_EAST_B17_sel_value_O;
	wire [16:0] RMUX_T2_NORTH_B17_O;
	wire RMUX_T2_NORTH_B17_ready_out;
	wire RMUX_T2_NORTH_B17_valid_out;
	wire [1:0] RMUX_T2_NORTH_B17_out_sel;
	wire [0:0] RMUX_T2_NORTH_B17_sel_value_O;
	wire [16:0] RMUX_T2_SOUTH_B17_O;
	wire RMUX_T2_SOUTH_B17_ready_out;
	wire RMUX_T2_SOUTH_B17_valid_out;
	wire [1:0] RMUX_T2_SOUTH_B17_out_sel;
	wire [0:0] RMUX_T2_SOUTH_B17_sel_value_O;
	wire [16:0] RMUX_T2_WEST_B17_O;
	wire RMUX_T2_WEST_B17_ready_out;
	wire RMUX_T2_WEST_B17_valid_out;
	wire [1:0] RMUX_T2_WEST_B17_out_sel;
	wire [0:0] RMUX_T2_WEST_B17_sel_value_O;
	wire [16:0] RMUX_T3_EAST_B17_O;
	wire RMUX_T3_EAST_B17_ready_out;
	wire RMUX_T3_EAST_B17_valid_out;
	wire [1:0] RMUX_T3_EAST_B17_out_sel;
	wire [0:0] RMUX_T3_EAST_B17_sel_value_O;
	wire [16:0] RMUX_T3_NORTH_B17_O;
	wire RMUX_T3_NORTH_B17_ready_out;
	wire RMUX_T3_NORTH_B17_valid_out;
	wire [1:0] RMUX_T3_NORTH_B17_out_sel;
	wire [0:0] RMUX_T3_NORTH_B17_sel_value_O;
	wire [16:0] RMUX_T3_SOUTH_B17_O;
	wire RMUX_T3_SOUTH_B17_ready_out;
	wire RMUX_T3_SOUTH_B17_valid_out;
	wire [1:0] RMUX_T3_SOUTH_B17_out_sel;
	wire [0:0] RMUX_T3_SOUTH_B17_sel_value_O;
	wire [16:0] RMUX_T3_WEST_B17_O;
	wire RMUX_T3_WEST_B17_ready_out;
	wire RMUX_T3_WEST_B17_valid_out;
	wire [1:0] RMUX_T3_WEST_B17_out_sel;
	wire [0:0] RMUX_T3_WEST_B17_sel_value_O;
	wire [16:0] RMUX_T4_EAST_B17_O;
	wire RMUX_T4_EAST_B17_ready_out;
	wire RMUX_T4_EAST_B17_valid_out;
	wire [1:0] RMUX_T4_EAST_B17_out_sel;
	wire [0:0] RMUX_T4_EAST_B17_sel_value_O;
	wire [16:0] RMUX_T4_NORTH_B17_O;
	wire RMUX_T4_NORTH_B17_ready_out;
	wire RMUX_T4_NORTH_B17_valid_out;
	wire [1:0] RMUX_T4_NORTH_B17_out_sel;
	wire [0:0] RMUX_T4_NORTH_B17_sel_value_O;
	wire [16:0] RMUX_T4_SOUTH_B17_O;
	wire RMUX_T4_SOUTH_B17_ready_out;
	wire RMUX_T4_SOUTH_B17_valid_out;
	wire [1:0] RMUX_T4_SOUTH_B17_out_sel;
	wire [0:0] RMUX_T4_SOUTH_B17_sel_value_O;
	wire [16:0] RMUX_T4_WEST_B17_O;
	wire RMUX_T4_WEST_B17_ready_out;
	wire RMUX_T4_WEST_B17_valid_out;
	wire [1:0] RMUX_T4_WEST_B17_out_sel;
	wire [0:0] RMUX_T4_WEST_B17_sel_value_O;
	wire [0:0] SB_T0_EAST_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T0_EAST_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T0_EAST_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T0_EAST_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T0_EAST_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T0_NORTH_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T0_NORTH_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T0_NORTH_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T0_NORTH_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T0_NORTH_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T0_SOUTH_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T0_SOUTH_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T0_SOUTH_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T0_SOUTH_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T0_SOUTH_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T0_WEST_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T0_WEST_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T0_WEST_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T0_WEST_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T0_WEST_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T1_EAST_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T1_EAST_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T1_EAST_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T1_EAST_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T1_EAST_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T1_NORTH_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T1_NORTH_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T1_NORTH_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T1_NORTH_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T1_NORTH_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T1_SOUTH_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T1_SOUTH_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T1_SOUTH_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T1_SOUTH_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T1_SOUTH_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T1_WEST_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T1_WEST_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T1_WEST_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T1_WEST_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T1_WEST_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T2_EAST_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T2_EAST_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T2_EAST_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T2_EAST_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T2_EAST_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T2_NORTH_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T2_NORTH_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T2_NORTH_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T2_NORTH_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T2_NORTH_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T2_SOUTH_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T2_SOUTH_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T2_SOUTH_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T2_SOUTH_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T2_SOUTH_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T2_WEST_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T2_WEST_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T2_WEST_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T2_WEST_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T2_WEST_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T3_EAST_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T3_EAST_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T3_EAST_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T3_EAST_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T3_EAST_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T3_NORTH_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T3_NORTH_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T3_NORTH_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T3_NORTH_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T3_NORTH_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T3_SOUTH_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T3_SOUTH_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T3_SOUTH_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T3_SOUTH_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T3_SOUTH_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T3_WEST_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T3_WEST_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T3_WEST_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T3_WEST_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T3_WEST_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T4_EAST_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T4_EAST_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T4_EAST_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T4_EAST_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T4_EAST_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T4_NORTH_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T4_NORTH_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T4_NORTH_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T4_NORTH_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T4_NORTH_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T4_SOUTH_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T4_SOUTH_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T4_SOUTH_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T4_SOUTH_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T4_SOUTH_SB_OUT_B17_sel_value_O;
	wire [0:0] SB_T4_WEST_SB_IN_B17_enable_value_O;
	wire [0:0] SB_T4_WEST_SB_IN_B17_fan_in_O;
	wire [0:0] SB_T4_WEST_SB_OUT_B17_FANOUT_O;
	wire [0:0] SB_T4_WEST_SB_OUT_B17_enable_value_O;
	wire [2:0] SB_T4_WEST_SB_OUT_B17_sel_value_O;
	wire [16:0] WIRE_SB_T0_EAST_SB_IN_B17_O;
	wire WIRE_SB_T0_EAST_SB_IN_B17_ready_out;
	wire WIRE_SB_T0_EAST_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T0_NORTH_SB_IN_B17_O;
	wire WIRE_SB_T0_NORTH_SB_IN_B17_ready_out;
	wire WIRE_SB_T0_NORTH_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T0_SOUTH_SB_IN_B17_O;
	wire WIRE_SB_T0_SOUTH_SB_IN_B17_ready_out;
	wire WIRE_SB_T0_SOUTH_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T0_WEST_SB_IN_B17_O;
	wire WIRE_SB_T0_WEST_SB_IN_B17_ready_out;
	wire WIRE_SB_T0_WEST_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T1_EAST_SB_IN_B17_O;
	wire WIRE_SB_T1_EAST_SB_IN_B17_ready_out;
	wire WIRE_SB_T1_EAST_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T1_NORTH_SB_IN_B17_O;
	wire WIRE_SB_T1_NORTH_SB_IN_B17_ready_out;
	wire WIRE_SB_T1_NORTH_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T1_SOUTH_SB_IN_B17_O;
	wire WIRE_SB_T1_SOUTH_SB_IN_B17_ready_out;
	wire WIRE_SB_T1_SOUTH_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T1_WEST_SB_IN_B17_O;
	wire WIRE_SB_T1_WEST_SB_IN_B17_ready_out;
	wire WIRE_SB_T1_WEST_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T2_EAST_SB_IN_B17_O;
	wire WIRE_SB_T2_EAST_SB_IN_B17_ready_out;
	wire WIRE_SB_T2_EAST_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T2_NORTH_SB_IN_B17_O;
	wire WIRE_SB_T2_NORTH_SB_IN_B17_ready_out;
	wire WIRE_SB_T2_NORTH_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T2_SOUTH_SB_IN_B17_O;
	wire WIRE_SB_T2_SOUTH_SB_IN_B17_ready_out;
	wire WIRE_SB_T2_SOUTH_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T2_WEST_SB_IN_B17_O;
	wire WIRE_SB_T2_WEST_SB_IN_B17_ready_out;
	wire WIRE_SB_T2_WEST_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T3_EAST_SB_IN_B17_O;
	wire WIRE_SB_T3_EAST_SB_IN_B17_ready_out;
	wire WIRE_SB_T3_EAST_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T3_NORTH_SB_IN_B17_O;
	wire WIRE_SB_T3_NORTH_SB_IN_B17_ready_out;
	wire WIRE_SB_T3_NORTH_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T3_SOUTH_SB_IN_B17_O;
	wire WIRE_SB_T3_SOUTH_SB_IN_B17_ready_out;
	wire WIRE_SB_T3_SOUTH_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T3_WEST_SB_IN_B17_O;
	wire WIRE_SB_T3_WEST_SB_IN_B17_ready_out;
	wire WIRE_SB_T3_WEST_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T4_EAST_SB_IN_B17_O;
	wire WIRE_SB_T4_EAST_SB_IN_B17_ready_out;
	wire WIRE_SB_T4_EAST_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T4_NORTH_SB_IN_B17_O;
	wire WIRE_SB_T4_NORTH_SB_IN_B17_ready_out;
	wire WIRE_SB_T4_NORTH_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T4_SOUTH_SB_IN_B17_O;
	wire WIRE_SB_T4_SOUTH_SB_IN_B17_ready_out;
	wire WIRE_SB_T4_SOUTH_SB_IN_B17_valid_out;
	wire [16:0] WIRE_SB_T4_WEST_SB_IN_B17_O;
	wire WIRE_SB_T4_WEST_SB_IN_B17_ready_out;
	wire WIRE_SB_T4_WEST_SB_IN_B17_valid_out;
	wire ZextWrapper_23_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_23_32_inst0$self_O_in;
	wire ZextWrapper_30_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_30_32_inst0$self_O_in;
	wire ZextWrapper_31_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_31_32_inst0$self_O_in;
	wire [0:0] and1_inst0_out;
	wire [0:0] and1_inst1_out;
	wire [0:0] and1_inst10_out;
	wire [0:0] and1_inst11_out;
	wire [0:0] and1_inst12_out;
	wire [0:0] and1_inst13_out;
	wire [0:0] and1_inst14_out;
	wire [0:0] and1_inst15_out;
	wire [0:0] and1_inst16_out;
	wire [0:0] and1_inst17_out;
	wire [0:0] and1_inst18_out;
	wire [0:0] and1_inst19_out;
	wire [0:0] and1_inst2_out;
	wire [0:0] and1_inst3_out;
	wire [0:0] and1_inst4_out;
	wire [0:0] and1_inst5_out;
	wire [0:0] and1_inst6_out;
	wire [0:0] and1_inst7_out;
	wire [0:0] and1_inst8_out;
	wire [0:0] and1_inst9_out;
	wire [31:0] config_reg_0_O;
	wire [31:0] config_reg_1_O;
	wire [31:0] config_reg_2_O;
	wire [30:0] config_reg_3_O;
	wire [29:0] config_reg_4_O;
	wire [22:0] config_reg_5_O;
	wire [0:0] const_1_1_out;
	wire coreir_eq_1_inst0_out;
	wire coreir_eq_1_inst1_out;
	wire coreir_eq_1_inst10_out;
	wire coreir_eq_1_inst11_out;
	wire coreir_eq_1_inst12_out;
	wire coreir_eq_1_inst13_out;
	wire coreir_eq_1_inst14_out;
	wire coreir_eq_1_inst15_out;
	wire coreir_eq_1_inst16_out;
	wire coreir_eq_1_inst17_out;
	wire coreir_eq_1_inst18_out;
	wire coreir_eq_1_inst19_out;
	wire coreir_eq_1_inst2_out;
	wire coreir_eq_1_inst3_out;
	wire coreir_eq_1_inst4_out;
	wire coreir_eq_1_inst5_out;
	wire coreir_eq_1_inst6_out;
	wire coreir_eq_1_inst7_out;
	wire coreir_eq_1_inst8_out;
	wire coreir_eq_1_inst9_out;
	wire [31:0] mux_aoi_6_32_inst0_O;
	wire [7:0] mux_aoi_6_32_inst0_out_sel;
	wire [7:0] self_config_config_addr_out;
	FanoutHash_E70AF988E4250F5 CB_MEM_output_width_17_num_0_fan_in(
		.I13(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
		.E8(SB_T2_NORTH_SB_OUT_B17_enable_value_O),
		.E17(SB_T4_SOUTH_SB_OUT_B17_enable_value_O),
		.I15(MUX_SB_T3_WEST_SB_OUT_B17_ready_out),
		.I12(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out),
		.E6(SB_T1_EAST_SB_OUT_B17_enable_value_O),
		.I9(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
		.I16(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
		.E3(SB_T0_WEST_SB_OUT_B17_enable_value_O),
		.S14(MUX_SB_T3_EAST_SB_OUT_B17_out_sel),
		.E10(SB_T2_EAST_SB_OUT_B17_enable_value_O),
		.I5(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
		.S6(MUX_SB_T1_EAST_SB_OUT_B17_out_sel),
		.E0(SB_T0_NORTH_SB_OUT_B17_enable_value_O),
		.E18(SB_T4_EAST_SB_OUT_B17_enable_value_O),
		.I19(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
		.I10(MUX_SB_T2_EAST_SB_OUT_B17_ready_out),
		.S5(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel),
		.I6(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
		.I8(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
		.S3(MUX_SB_T0_WEST_SB_OUT_B17_out_sel),
		.S10(MUX_SB_T2_EAST_SB_OUT_B17_out_sel),
		.E16(SB_T4_NORTH_SB_OUT_B17_enable_value_O),
		.S4(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel),
		.E11(SB_T2_WEST_SB_OUT_B17_enable_value_O),
		.S19(MUX_SB_T4_WEST_SB_OUT_B17_out_sel),
		.E15(SB_T3_WEST_SB_OUT_B17_enable_value_O),
		.E19(SB_T4_WEST_SB_OUT_B17_enable_value_O),
		.I3(MUX_SB_T0_WEST_SB_OUT_B17_ready_out),
		.I4(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out),
		.S1(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel),
		.E13(SB_T3_SOUTH_SB_OUT_B17_enable_value_O),
		.S0(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T0_EAST_SB_OUT_B17_out_sel),
		.I11(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
		.S8(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel),
		.E2(SB_T0_EAST_SB_OUT_B17_enable_value_O),
		.E14(SB_T3_EAST_SB_OUT_B17_enable_value_O),
		.S17(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel),
		.E5(SB_T1_SOUTH_SB_OUT_B17_enable_value_O),
		.E4(SB_T1_NORTH_SB_OUT_B17_enable_value_O),
		.I1(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
		.I2(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
		.I17(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
		.O(CB_MEM_output_width_17_num_0_fan_in_O),
		.E9(SB_T2_SOUTH_SB_OUT_B17_enable_value_O),
		.S13(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel),
		.S11(MUX_SB_T2_WEST_SB_OUT_B17_out_sel),
		.S7(MUX_SB_T1_WEST_SB_OUT_B17_out_sel),
		.E1(SB_T0_SOUTH_SB_OUT_B17_enable_value_O),
		.S15(MUX_SB_T3_WEST_SB_OUT_B17_out_sel),
		.S9(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel),
		.S18(MUX_SB_T4_EAST_SB_OUT_B17_out_sel),
		.S12(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel),
		.I14(MUX_SB_T3_EAST_SB_OUT_B17_ready_out),
		.I7(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
		.S16(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel),
		.E12(SB_T3_NORTH_SB_OUT_B17_enable_value_O),
		.I0(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out),
		.E7(SB_T1_WEST_SB_OUT_B17_enable_value_O),
		.I18(MUX_SB_T4_EAST_SB_OUT_B17_ready_out)
	);
	FanoutHash_82899D6851EDC11 CB_MEM_output_width_17_num_1_fan_in(
		.I13(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
		.E8(SB_T2_NORTH_SB_OUT_B17_enable_value_O),
		.E17(SB_T4_SOUTH_SB_OUT_B17_enable_value_O),
		.I15(MUX_SB_T3_WEST_SB_OUT_B17_ready_out),
		.I12(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out),
		.E6(SB_T1_EAST_SB_OUT_B17_enable_value_O),
		.I9(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
		.I16(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
		.E3(SB_T0_WEST_SB_OUT_B17_enable_value_O),
		.S14(MUX_SB_T3_EAST_SB_OUT_B17_out_sel),
		.E10(SB_T2_EAST_SB_OUT_B17_enable_value_O),
		.I5(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
		.S6(MUX_SB_T1_EAST_SB_OUT_B17_out_sel),
		.E0(SB_T0_NORTH_SB_OUT_B17_enable_value_O),
		.E18(SB_T4_EAST_SB_OUT_B17_enable_value_O),
		.I19(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
		.I10(MUX_SB_T2_EAST_SB_OUT_B17_ready_out),
		.S5(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel),
		.I6(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
		.I8(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
		.S3(MUX_SB_T0_WEST_SB_OUT_B17_out_sel),
		.S10(MUX_SB_T2_EAST_SB_OUT_B17_out_sel),
		.E16(SB_T4_NORTH_SB_OUT_B17_enable_value_O),
		.S4(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel),
		.E11(SB_T2_WEST_SB_OUT_B17_enable_value_O),
		.S19(MUX_SB_T4_WEST_SB_OUT_B17_out_sel),
		.E15(SB_T3_WEST_SB_OUT_B17_enable_value_O),
		.E19(SB_T4_WEST_SB_OUT_B17_enable_value_O),
		.I3(MUX_SB_T0_WEST_SB_OUT_B17_ready_out),
		.I4(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out),
		.S1(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel),
		.E13(SB_T3_SOUTH_SB_OUT_B17_enable_value_O),
		.S0(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T0_EAST_SB_OUT_B17_out_sel),
		.I11(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
		.S8(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel),
		.E2(SB_T0_EAST_SB_OUT_B17_enable_value_O),
		.E14(SB_T3_EAST_SB_OUT_B17_enable_value_O),
		.S17(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel),
		.E5(SB_T1_SOUTH_SB_OUT_B17_enable_value_O),
		.E4(SB_T1_NORTH_SB_OUT_B17_enable_value_O),
		.I1(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
		.I2(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
		.I17(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
		.O(CB_MEM_output_width_17_num_1_fan_in_O),
		.E9(SB_T2_SOUTH_SB_OUT_B17_enable_value_O),
		.S13(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel),
		.S11(MUX_SB_T2_WEST_SB_OUT_B17_out_sel),
		.S7(MUX_SB_T1_WEST_SB_OUT_B17_out_sel),
		.E1(SB_T0_SOUTH_SB_OUT_B17_enable_value_O),
		.S15(MUX_SB_T3_WEST_SB_OUT_B17_out_sel),
		.S9(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel),
		.S18(MUX_SB_T4_EAST_SB_OUT_B17_out_sel),
		.S12(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel),
		.I14(MUX_SB_T3_EAST_SB_OUT_B17_ready_out),
		.I7(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
		.S16(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel),
		.E12(SB_T3_NORTH_SB_OUT_B17_enable_value_O),
		.I0(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out),
		.E7(SB_T1_WEST_SB_OUT_B17_enable_value_O),
		.I18(MUX_SB_T4_EAST_SB_OUT_B17_ready_out)
	);
	FanoutHash_CE1AA874B742213 CB_MEM_output_width_17_num_2_fan_in(
		.I13(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
		.E8(SB_T2_NORTH_SB_OUT_B17_enable_value_O),
		.E17(SB_T4_SOUTH_SB_OUT_B17_enable_value_O),
		.I15(MUX_SB_T3_WEST_SB_OUT_B17_ready_out),
		.I12(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out),
		.E6(SB_T1_EAST_SB_OUT_B17_enable_value_O),
		.I9(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
		.I16(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
		.E3(SB_T0_WEST_SB_OUT_B17_enable_value_O),
		.S14(MUX_SB_T3_EAST_SB_OUT_B17_out_sel),
		.E10(SB_T2_EAST_SB_OUT_B17_enable_value_O),
		.I5(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
		.S6(MUX_SB_T1_EAST_SB_OUT_B17_out_sel),
		.E0(SB_T0_NORTH_SB_OUT_B17_enable_value_O),
		.E18(SB_T4_EAST_SB_OUT_B17_enable_value_O),
		.I19(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
		.I10(MUX_SB_T2_EAST_SB_OUT_B17_ready_out),
		.S5(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel),
		.I6(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
		.I8(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
		.S3(MUX_SB_T0_WEST_SB_OUT_B17_out_sel),
		.S10(MUX_SB_T2_EAST_SB_OUT_B17_out_sel),
		.E16(SB_T4_NORTH_SB_OUT_B17_enable_value_O),
		.S4(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel),
		.E11(SB_T2_WEST_SB_OUT_B17_enable_value_O),
		.S19(MUX_SB_T4_WEST_SB_OUT_B17_out_sel),
		.E15(SB_T3_WEST_SB_OUT_B17_enable_value_O),
		.E19(SB_T4_WEST_SB_OUT_B17_enable_value_O),
		.I3(MUX_SB_T0_WEST_SB_OUT_B17_ready_out),
		.I4(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out),
		.S1(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel),
		.E13(SB_T3_SOUTH_SB_OUT_B17_enable_value_O),
		.S0(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T0_EAST_SB_OUT_B17_out_sel),
		.I11(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
		.S8(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel),
		.E2(SB_T0_EAST_SB_OUT_B17_enable_value_O),
		.E14(SB_T3_EAST_SB_OUT_B17_enable_value_O),
		.S17(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel),
		.E5(SB_T1_SOUTH_SB_OUT_B17_enable_value_O),
		.E4(SB_T1_NORTH_SB_OUT_B17_enable_value_O),
		.I1(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
		.I2(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
		.I17(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
		.O(CB_MEM_output_width_17_num_2_fan_in_O),
		.E9(SB_T2_SOUTH_SB_OUT_B17_enable_value_O),
		.S13(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel),
		.S11(MUX_SB_T2_WEST_SB_OUT_B17_out_sel),
		.S7(MUX_SB_T1_WEST_SB_OUT_B17_out_sel),
		.E1(SB_T0_SOUTH_SB_OUT_B17_enable_value_O),
		.S15(MUX_SB_T3_WEST_SB_OUT_B17_out_sel),
		.S9(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel),
		.S18(MUX_SB_T4_EAST_SB_OUT_B17_out_sel),
		.S12(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel),
		.I14(MUX_SB_T3_EAST_SB_OUT_B17_ready_out),
		.I7(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
		.S16(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel),
		.E12(SB_T3_NORTH_SB_OUT_B17_enable_value_O),
		.I0(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out),
		.E7(SB_T1_WEST_SB_OUT_B17_enable_value_O),
		.I18(MUX_SB_T4_EAST_SB_OUT_B17_ready_out)
	);
	coreir_not #(.width(1)) Invert1_inst0(
		.in(stall),
		.out(Invert1_inst0_out)
	);
	wire [101:0] MUX_SB_T0_EAST_SB_OUT_B17_I;
	assign MUX_SB_T0_EAST_SB_OUT_B17_I[85+:17] = MEM_output_width_17_num_2;
	assign MUX_SB_T0_EAST_SB_OUT_B17_I[68+:17] = MEM_output_width_17_num_1;
	assign MUX_SB_T0_EAST_SB_OUT_B17_I[51+:17] = MEM_output_width_17_num_0;
	assign MUX_SB_T0_EAST_SB_OUT_B17_I[34+:17] = WIRE_SB_T4_NORTH_SB_IN_B17_O;
	assign MUX_SB_T0_EAST_SB_OUT_B17_I[17+:17] = WIRE_SB_T3_SOUTH_SB_IN_B17_O;
	assign MUX_SB_T0_EAST_SB_OUT_B17_I[0+:17] = WIRE_SB_T0_WEST_SB_IN_B17_O;
	wire [5:0] MUX_SB_T0_EAST_SB_OUT_B17_valid_in;
	assign MUX_SB_T0_EAST_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid, MEM_output_width_17_num_1_valid, MEM_output_width_17_num_0_valid, WIRE_SB_T4_NORTH_SB_IN_B17_valid_out, WIRE_SB_T3_SOUTH_SB_IN_B17_valid_out, WIRE_SB_T0_WEST_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_6_17 MUX_SB_T0_EAST_SB_OUT_B17(
		.I(MUX_SB_T0_EAST_SB_OUT_B17_I),
		.O(MUX_SB_T0_EAST_SB_OUT_B17_O),
		.ready_in(SB_T0_EAST_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T0_EAST_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T0_EAST_SB_OUT_B17_valid_out),
		.S(SB_T0_EAST_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T0_EAST_SB_OUT_B17_out_sel)
	);
	wire [101:0] MUX_SB_T0_NORTH_SB_OUT_B17_I;
	assign MUX_SB_T0_NORTH_SB_OUT_B17_I[85+:17] = MEM_output_width_17_num_2;
	assign MUX_SB_T0_NORTH_SB_OUT_B17_I[68+:17] = MEM_output_width_17_num_1;
	assign MUX_SB_T0_NORTH_SB_OUT_B17_I[51+:17] = MEM_output_width_17_num_0;
	assign MUX_SB_T0_NORTH_SB_OUT_B17_I[34+:17] = WIRE_SB_T0_SOUTH_SB_IN_B17_O;
	assign MUX_SB_T0_NORTH_SB_OUT_B17_I[17+:17] = WIRE_SB_T1_EAST_SB_IN_B17_O;
	assign MUX_SB_T0_NORTH_SB_OUT_B17_I[0+:17] = WIRE_SB_T0_WEST_SB_IN_B17_O;
	wire [5:0] MUX_SB_T0_NORTH_SB_OUT_B17_valid_in;
	assign MUX_SB_T0_NORTH_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid, MEM_output_width_17_num_1_valid, MEM_output_width_17_num_0_valid, WIRE_SB_T0_SOUTH_SB_IN_B17_valid_out, WIRE_SB_T1_EAST_SB_IN_B17_valid_out, WIRE_SB_T0_WEST_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_6_17 MUX_SB_T0_NORTH_SB_OUT_B17(
		.I(MUX_SB_T0_NORTH_SB_OUT_B17_I),
		.O(MUX_SB_T0_NORTH_SB_OUT_B17_O),
		.ready_in(SB_T0_NORTH_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T0_NORTH_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T0_NORTH_SB_OUT_B17_valid_out),
		.S(SB_T0_NORTH_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel)
	);
	wire [101:0] MUX_SB_T0_SOUTH_SB_OUT_B17_I;
	assign MUX_SB_T0_SOUTH_SB_OUT_B17_I[85+:17] = MEM_output_width_17_num_2;
	assign MUX_SB_T0_SOUTH_SB_OUT_B17_I[68+:17] = MEM_output_width_17_num_1;
	assign MUX_SB_T0_SOUTH_SB_OUT_B17_I[51+:17] = MEM_output_width_17_num_0;
	assign MUX_SB_T0_SOUTH_SB_OUT_B17_I[34+:17] = WIRE_SB_T1_WEST_SB_IN_B17_O;
	assign MUX_SB_T0_SOUTH_SB_OUT_B17_I[17+:17] = WIRE_SB_T0_NORTH_SB_IN_B17_O;
	assign MUX_SB_T0_SOUTH_SB_OUT_B17_I[0+:17] = WIRE_SB_T3_EAST_SB_IN_B17_O;
	wire [5:0] MUX_SB_T0_SOUTH_SB_OUT_B17_valid_in;
	assign MUX_SB_T0_SOUTH_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid, MEM_output_width_17_num_1_valid, MEM_output_width_17_num_0_valid, WIRE_SB_T1_WEST_SB_IN_B17_valid_out, WIRE_SB_T0_NORTH_SB_IN_B17_valid_out, WIRE_SB_T3_EAST_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_6_17 MUX_SB_T0_SOUTH_SB_OUT_B17(
		.I(MUX_SB_T0_SOUTH_SB_OUT_B17_I),
		.O(MUX_SB_T0_SOUTH_SB_OUT_B17_O),
		.ready_in(SB_T0_SOUTH_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T0_SOUTH_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T0_SOUTH_SB_OUT_B17_valid_out),
		.S(SB_T0_SOUTH_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel)
	);
	wire [101:0] MUX_SB_T0_WEST_SB_OUT_B17_I;
	assign MUX_SB_T0_WEST_SB_OUT_B17_I[85+:17] = MEM_output_width_17_num_2;
	assign MUX_SB_T0_WEST_SB_OUT_B17_I[68+:17] = MEM_output_width_17_num_1;
	assign MUX_SB_T0_WEST_SB_OUT_B17_I[51+:17] = MEM_output_width_17_num_0;
	assign MUX_SB_T0_WEST_SB_OUT_B17_I[34+:17] = WIRE_SB_T0_EAST_SB_IN_B17_O;
	assign MUX_SB_T0_WEST_SB_OUT_B17_I[17+:17] = WIRE_SB_T4_SOUTH_SB_IN_B17_O;
	assign MUX_SB_T0_WEST_SB_OUT_B17_I[0+:17] = WIRE_SB_T0_NORTH_SB_IN_B17_O;
	wire [5:0] MUX_SB_T0_WEST_SB_OUT_B17_valid_in;
	assign MUX_SB_T0_WEST_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid, MEM_output_width_17_num_1_valid, MEM_output_width_17_num_0_valid, WIRE_SB_T0_EAST_SB_IN_B17_valid_out, WIRE_SB_T4_SOUTH_SB_IN_B17_valid_out, WIRE_SB_T0_NORTH_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_6_17 MUX_SB_T0_WEST_SB_OUT_B17(
		.I(MUX_SB_T0_WEST_SB_OUT_B17_I),
		.O(MUX_SB_T0_WEST_SB_OUT_B17_O),
		.ready_in(SB_T0_WEST_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T0_WEST_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T0_WEST_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T0_WEST_SB_OUT_B17_valid_out),
		.S(SB_T0_WEST_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T0_WEST_SB_OUT_B17_out_sel)
	);
	wire [101:0] MUX_SB_T1_EAST_SB_OUT_B17_I;
	assign MUX_SB_T1_EAST_SB_OUT_B17_I[85+:17] = MEM_output_width_17_num_2;
	assign MUX_SB_T1_EAST_SB_OUT_B17_I[68+:17] = MEM_output_width_17_num_1;
	assign MUX_SB_T1_EAST_SB_OUT_B17_I[51+:17] = MEM_output_width_17_num_0;
	assign MUX_SB_T1_EAST_SB_OUT_B17_I[34+:17] = WIRE_SB_T2_SOUTH_SB_IN_B17_O;
	assign MUX_SB_T1_EAST_SB_OUT_B17_I[17+:17] = WIRE_SB_T1_WEST_SB_IN_B17_O;
	assign MUX_SB_T1_EAST_SB_OUT_B17_I[0+:17] = WIRE_SB_T0_NORTH_SB_IN_B17_O;
	wire [5:0] MUX_SB_T1_EAST_SB_OUT_B17_valid_in;
	assign MUX_SB_T1_EAST_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid, MEM_output_width_17_num_1_valid, MEM_output_width_17_num_0_valid, WIRE_SB_T2_SOUTH_SB_IN_B17_valid_out, WIRE_SB_T1_WEST_SB_IN_B17_valid_out, WIRE_SB_T0_NORTH_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_6_17 MUX_SB_T1_EAST_SB_OUT_B17(
		.I(MUX_SB_T1_EAST_SB_OUT_B17_I),
		.O(MUX_SB_T1_EAST_SB_OUT_B17_O),
		.ready_in(SB_T1_EAST_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T1_EAST_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T1_EAST_SB_OUT_B17_valid_out),
		.S(SB_T1_EAST_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T1_EAST_SB_OUT_B17_out_sel)
	);
	wire [101:0] MUX_SB_T1_NORTH_SB_OUT_B17_I;
	assign MUX_SB_T1_NORTH_SB_OUT_B17_I[85+:17] = MEM_output_width_17_num_2;
	assign MUX_SB_T1_NORTH_SB_OUT_B17_I[68+:17] = MEM_output_width_17_num_1;
	assign MUX_SB_T1_NORTH_SB_OUT_B17_I[51+:17] = MEM_output_width_17_num_0;
	assign MUX_SB_T1_NORTH_SB_OUT_B17_I[34+:17] = WIRE_SB_T4_WEST_SB_IN_B17_O;
	assign MUX_SB_T1_NORTH_SB_OUT_B17_I[17+:17] = WIRE_SB_T1_SOUTH_SB_IN_B17_O;
	assign MUX_SB_T1_NORTH_SB_OUT_B17_I[0+:17] = WIRE_SB_T2_EAST_SB_IN_B17_O;
	wire [5:0] MUX_SB_T1_NORTH_SB_OUT_B17_valid_in;
	assign MUX_SB_T1_NORTH_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid, MEM_output_width_17_num_1_valid, MEM_output_width_17_num_0_valid, WIRE_SB_T4_WEST_SB_IN_B17_valid_out, WIRE_SB_T1_SOUTH_SB_IN_B17_valid_out, WIRE_SB_T2_EAST_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_6_17 MUX_SB_T1_NORTH_SB_OUT_B17(
		.I(MUX_SB_T1_NORTH_SB_OUT_B17_I),
		.O(MUX_SB_T1_NORTH_SB_OUT_B17_O),
		.ready_in(SB_T1_NORTH_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T1_NORTH_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T1_NORTH_SB_OUT_B17_valid_out),
		.S(SB_T1_NORTH_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel)
	);
	wire [101:0] MUX_SB_T1_SOUTH_SB_OUT_B17_I;
	assign MUX_SB_T1_SOUTH_SB_OUT_B17_I[85+:17] = MEM_output_width_17_num_2;
	assign MUX_SB_T1_SOUTH_SB_OUT_B17_I[68+:17] = MEM_output_width_17_num_1;
	assign MUX_SB_T1_SOUTH_SB_OUT_B17_I[51+:17] = MEM_output_width_17_num_0;
	assign MUX_SB_T1_SOUTH_SB_OUT_B17_I[34+:17] = WIRE_SB_T2_WEST_SB_IN_B17_O;
	assign MUX_SB_T1_SOUTH_SB_OUT_B17_I[17+:17] = WIRE_SB_T1_NORTH_SB_IN_B17_O;
	assign MUX_SB_T1_SOUTH_SB_OUT_B17_I[0+:17] = WIRE_SB_T2_EAST_SB_IN_B17_O;
	wire [5:0] MUX_SB_T1_SOUTH_SB_OUT_B17_valid_in;
	assign MUX_SB_T1_SOUTH_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid, MEM_output_width_17_num_1_valid, MEM_output_width_17_num_0_valid, WIRE_SB_T2_WEST_SB_IN_B17_valid_out, WIRE_SB_T1_NORTH_SB_IN_B17_valid_out, WIRE_SB_T2_EAST_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_6_17 MUX_SB_T1_SOUTH_SB_OUT_B17(
		.I(MUX_SB_T1_SOUTH_SB_OUT_B17_I),
		.O(MUX_SB_T1_SOUTH_SB_OUT_B17_O),
		.ready_in(SB_T1_SOUTH_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T1_SOUTH_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T1_SOUTH_SB_OUT_B17_valid_out),
		.S(SB_T1_SOUTH_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel)
	);
	wire [101:0] MUX_SB_T1_WEST_SB_OUT_B17_I;
	assign MUX_SB_T1_WEST_SB_OUT_B17_I[85+:17] = MEM_output_width_17_num_2;
	assign MUX_SB_T1_WEST_SB_OUT_B17_I[68+:17] = MEM_output_width_17_num_1;
	assign MUX_SB_T1_WEST_SB_OUT_B17_I[51+:17] = MEM_output_width_17_num_0;
	assign MUX_SB_T1_WEST_SB_OUT_B17_I[34+:17] = WIRE_SB_T1_EAST_SB_IN_B17_O;
	assign MUX_SB_T1_WEST_SB_OUT_B17_I[17+:17] = WIRE_SB_T0_SOUTH_SB_IN_B17_O;
	assign MUX_SB_T1_WEST_SB_OUT_B17_I[0+:17] = WIRE_SB_T4_NORTH_SB_IN_B17_O;
	wire [5:0] MUX_SB_T1_WEST_SB_OUT_B17_valid_in;
	assign MUX_SB_T1_WEST_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid, MEM_output_width_17_num_1_valid, MEM_output_width_17_num_0_valid, WIRE_SB_T1_EAST_SB_IN_B17_valid_out, WIRE_SB_T0_SOUTH_SB_IN_B17_valid_out, WIRE_SB_T4_NORTH_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_6_17 MUX_SB_T1_WEST_SB_OUT_B17(
		.I(MUX_SB_T1_WEST_SB_OUT_B17_I),
		.O(MUX_SB_T1_WEST_SB_OUT_B17_O),
		.ready_in(SB_T1_WEST_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T1_WEST_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T1_WEST_SB_OUT_B17_valid_out),
		.S(SB_T1_WEST_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T1_WEST_SB_OUT_B17_out_sel)
	);
	wire [101:0] MUX_SB_T2_EAST_SB_OUT_B17_I;
	assign MUX_SB_T2_EAST_SB_OUT_B17_I[85+:17] = MEM_output_width_17_num_2;
	assign MUX_SB_T2_EAST_SB_OUT_B17_I[68+:17] = MEM_output_width_17_num_1;
	assign MUX_SB_T2_EAST_SB_OUT_B17_I[51+:17] = MEM_output_width_17_num_0;
	assign MUX_SB_T2_EAST_SB_OUT_B17_I[34+:17] = WIRE_SB_T2_WEST_SB_IN_B17_O;
	assign MUX_SB_T2_EAST_SB_OUT_B17_I[17+:17] = WIRE_SB_T1_SOUTH_SB_IN_B17_O;
	assign MUX_SB_T2_EAST_SB_OUT_B17_I[0+:17] = WIRE_SB_T1_NORTH_SB_IN_B17_O;
	wire [5:0] MUX_SB_T2_EAST_SB_OUT_B17_valid_in;
	assign MUX_SB_T2_EAST_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid, MEM_output_width_17_num_1_valid, MEM_output_width_17_num_0_valid, WIRE_SB_T2_WEST_SB_IN_B17_valid_out, WIRE_SB_T1_SOUTH_SB_IN_B17_valid_out, WIRE_SB_T1_NORTH_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_6_17 MUX_SB_T2_EAST_SB_OUT_B17(
		.I(MUX_SB_T2_EAST_SB_OUT_B17_I),
		.O(MUX_SB_T2_EAST_SB_OUT_B17_O),
		.ready_in(SB_T2_EAST_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T2_EAST_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T2_EAST_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T2_EAST_SB_OUT_B17_valid_out),
		.S(SB_T2_EAST_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T2_EAST_SB_OUT_B17_out_sel)
	);
	wire [101:0] MUX_SB_T2_NORTH_SB_OUT_B17_I;
	assign MUX_SB_T2_NORTH_SB_OUT_B17_I[85+:17] = MEM_output_width_17_num_2;
	assign MUX_SB_T2_NORTH_SB_OUT_B17_I[68+:17] = MEM_output_width_17_num_1;
	assign MUX_SB_T2_NORTH_SB_OUT_B17_I[51+:17] = MEM_output_width_17_num_0;
	assign MUX_SB_T2_NORTH_SB_OUT_B17_I[34+:17] = WIRE_SB_T3_WEST_SB_IN_B17_O;
	assign MUX_SB_T2_NORTH_SB_OUT_B17_I[17+:17] = WIRE_SB_T2_SOUTH_SB_IN_B17_O;
	assign MUX_SB_T2_NORTH_SB_OUT_B17_I[0+:17] = WIRE_SB_T3_EAST_SB_IN_B17_O;
	wire [5:0] MUX_SB_T2_NORTH_SB_OUT_B17_valid_in;
	assign MUX_SB_T2_NORTH_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid, MEM_output_width_17_num_1_valid, MEM_output_width_17_num_0_valid, WIRE_SB_T3_WEST_SB_IN_B17_valid_out, WIRE_SB_T2_SOUTH_SB_IN_B17_valid_out, WIRE_SB_T3_EAST_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_6_17 MUX_SB_T2_NORTH_SB_OUT_B17(
		.I(MUX_SB_T2_NORTH_SB_OUT_B17_I),
		.O(MUX_SB_T2_NORTH_SB_OUT_B17_O),
		.ready_in(SB_T2_NORTH_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T2_NORTH_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T2_NORTH_SB_OUT_B17_valid_out),
		.S(SB_T2_NORTH_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel)
	);
	wire [101:0] MUX_SB_T2_SOUTH_SB_OUT_B17_I;
	assign MUX_SB_T2_SOUTH_SB_OUT_B17_I[85+:17] = MEM_output_width_17_num_2;
	assign MUX_SB_T2_SOUTH_SB_OUT_B17_I[68+:17] = MEM_output_width_17_num_1;
	assign MUX_SB_T2_SOUTH_SB_OUT_B17_I[51+:17] = MEM_output_width_17_num_0;
	assign MUX_SB_T2_SOUTH_SB_OUT_B17_I[34+:17] = WIRE_SB_T3_WEST_SB_IN_B17_O;
	assign MUX_SB_T2_SOUTH_SB_OUT_B17_I[17+:17] = WIRE_SB_T2_NORTH_SB_IN_B17_O;
	assign MUX_SB_T2_SOUTH_SB_OUT_B17_I[0+:17] = WIRE_SB_T1_EAST_SB_IN_B17_O;
	wire [5:0] MUX_SB_T2_SOUTH_SB_OUT_B17_valid_in;
	assign MUX_SB_T2_SOUTH_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid, MEM_output_width_17_num_1_valid, MEM_output_width_17_num_0_valid, WIRE_SB_T3_WEST_SB_IN_B17_valid_out, WIRE_SB_T2_NORTH_SB_IN_B17_valid_out, WIRE_SB_T1_EAST_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_6_17 MUX_SB_T2_SOUTH_SB_OUT_B17(
		.I(MUX_SB_T2_SOUTH_SB_OUT_B17_I),
		.O(MUX_SB_T2_SOUTH_SB_OUT_B17_O),
		.ready_in(SB_T2_SOUTH_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T2_SOUTH_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T2_SOUTH_SB_OUT_B17_valid_out),
		.S(SB_T2_SOUTH_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel)
	);
	wire [101:0] MUX_SB_T2_WEST_SB_OUT_B17_I;
	assign MUX_SB_T2_WEST_SB_OUT_B17_I[85+:17] = MEM_output_width_17_num_2;
	assign MUX_SB_T2_WEST_SB_OUT_B17_I[68+:17] = MEM_output_width_17_num_1;
	assign MUX_SB_T2_WEST_SB_OUT_B17_I[51+:17] = MEM_output_width_17_num_0;
	assign MUX_SB_T2_WEST_SB_OUT_B17_I[34+:17] = WIRE_SB_T2_EAST_SB_IN_B17_O;
	assign MUX_SB_T2_WEST_SB_OUT_B17_I[17+:17] = WIRE_SB_T1_SOUTH_SB_IN_B17_O;
	assign MUX_SB_T2_WEST_SB_OUT_B17_I[0+:17] = WIRE_SB_T3_NORTH_SB_IN_B17_O;
	wire [5:0] MUX_SB_T2_WEST_SB_OUT_B17_valid_in;
	assign MUX_SB_T2_WEST_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid, MEM_output_width_17_num_1_valid, MEM_output_width_17_num_0_valid, WIRE_SB_T2_EAST_SB_IN_B17_valid_out, WIRE_SB_T1_SOUTH_SB_IN_B17_valid_out, WIRE_SB_T3_NORTH_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_6_17 MUX_SB_T2_WEST_SB_OUT_B17(
		.I(MUX_SB_T2_WEST_SB_OUT_B17_I),
		.O(MUX_SB_T2_WEST_SB_OUT_B17_O),
		.ready_in(SB_T2_WEST_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T2_WEST_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T2_WEST_SB_OUT_B17_valid_out),
		.S(SB_T2_WEST_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T2_WEST_SB_OUT_B17_out_sel)
	);
	wire [101:0] MUX_SB_T3_EAST_SB_OUT_B17_I;
	assign MUX_SB_T3_EAST_SB_OUT_B17_I[85+:17] = MEM_output_width_17_num_2;
	assign MUX_SB_T3_EAST_SB_OUT_B17_I[68+:17] = MEM_output_width_17_num_1;
	assign MUX_SB_T3_EAST_SB_OUT_B17_I[51+:17] = MEM_output_width_17_num_0;
	assign MUX_SB_T3_EAST_SB_OUT_B17_I[34+:17] = WIRE_SB_T3_WEST_SB_IN_B17_O;
	assign MUX_SB_T3_EAST_SB_OUT_B17_I[17+:17] = WIRE_SB_T2_NORTH_SB_IN_B17_O;
	assign MUX_SB_T3_EAST_SB_OUT_B17_I[0+:17] = WIRE_SB_T0_SOUTH_SB_IN_B17_O;
	wire [5:0] MUX_SB_T3_EAST_SB_OUT_B17_valid_in;
	assign MUX_SB_T3_EAST_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid, MEM_output_width_17_num_1_valid, MEM_output_width_17_num_0_valid, WIRE_SB_T3_WEST_SB_IN_B17_valid_out, WIRE_SB_T2_NORTH_SB_IN_B17_valid_out, WIRE_SB_T0_SOUTH_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_6_17 MUX_SB_T3_EAST_SB_OUT_B17(
		.I(MUX_SB_T3_EAST_SB_OUT_B17_I),
		.O(MUX_SB_T3_EAST_SB_OUT_B17_O),
		.ready_in(SB_T3_EAST_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T3_EAST_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T3_EAST_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T3_EAST_SB_OUT_B17_valid_out),
		.S(SB_T3_EAST_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T3_EAST_SB_OUT_B17_out_sel)
	);
	wire [101:0] MUX_SB_T3_NORTH_SB_OUT_B17_I;
	assign MUX_SB_T3_NORTH_SB_OUT_B17_I[85+:17] = MEM_output_width_17_num_2;
	assign MUX_SB_T3_NORTH_SB_OUT_B17_I[68+:17] = MEM_output_width_17_num_1;
	assign MUX_SB_T3_NORTH_SB_OUT_B17_I[51+:17] = MEM_output_width_17_num_0;
	assign MUX_SB_T3_NORTH_SB_OUT_B17_I[34+:17] = WIRE_SB_T3_SOUTH_SB_IN_B17_O;
	assign MUX_SB_T3_NORTH_SB_OUT_B17_I[17+:17] = WIRE_SB_T4_EAST_SB_IN_B17_O;
	assign MUX_SB_T3_NORTH_SB_OUT_B17_I[0+:17] = WIRE_SB_T2_WEST_SB_IN_B17_O;
	wire [5:0] MUX_SB_T3_NORTH_SB_OUT_B17_valid_in;
	assign MUX_SB_T3_NORTH_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid, MEM_output_width_17_num_1_valid, MEM_output_width_17_num_0_valid, WIRE_SB_T3_SOUTH_SB_IN_B17_valid_out, WIRE_SB_T4_EAST_SB_IN_B17_valid_out, WIRE_SB_T2_WEST_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_6_17 MUX_SB_T3_NORTH_SB_OUT_B17(
		.I(MUX_SB_T3_NORTH_SB_OUT_B17_I),
		.O(MUX_SB_T3_NORTH_SB_OUT_B17_O),
		.ready_in(SB_T3_NORTH_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T3_NORTH_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T3_NORTH_SB_OUT_B17_valid_out),
		.S(SB_T3_NORTH_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel)
	);
	wire [101:0] MUX_SB_T3_SOUTH_SB_OUT_B17_I;
	assign MUX_SB_T3_SOUTH_SB_OUT_B17_I[85+:17] = MEM_output_width_17_num_2;
	assign MUX_SB_T3_SOUTH_SB_OUT_B17_I[68+:17] = MEM_output_width_17_num_1;
	assign MUX_SB_T3_SOUTH_SB_OUT_B17_I[51+:17] = MEM_output_width_17_num_0;
	assign MUX_SB_T3_SOUTH_SB_OUT_B17_I[34+:17] = WIRE_SB_T4_WEST_SB_IN_B17_O;
	assign MUX_SB_T3_SOUTH_SB_OUT_B17_I[17+:17] = WIRE_SB_T3_NORTH_SB_IN_B17_O;
	assign MUX_SB_T3_SOUTH_SB_OUT_B17_I[0+:17] = WIRE_SB_T0_EAST_SB_IN_B17_O;
	wire [5:0] MUX_SB_T3_SOUTH_SB_OUT_B17_valid_in;
	assign MUX_SB_T3_SOUTH_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid, MEM_output_width_17_num_1_valid, MEM_output_width_17_num_0_valid, WIRE_SB_T4_WEST_SB_IN_B17_valid_out, WIRE_SB_T3_NORTH_SB_IN_B17_valid_out, WIRE_SB_T0_EAST_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_6_17 MUX_SB_T3_SOUTH_SB_OUT_B17(
		.I(MUX_SB_T3_SOUTH_SB_OUT_B17_I),
		.O(MUX_SB_T3_SOUTH_SB_OUT_B17_O),
		.ready_in(SB_T3_SOUTH_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T3_SOUTH_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T3_SOUTH_SB_OUT_B17_valid_out),
		.S(SB_T3_SOUTH_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel)
	);
	wire [101:0] MUX_SB_T3_WEST_SB_OUT_B17_I;
	assign MUX_SB_T3_WEST_SB_OUT_B17_I[85+:17] = MEM_output_width_17_num_2;
	assign MUX_SB_T3_WEST_SB_OUT_B17_I[68+:17] = MEM_output_width_17_num_1;
	assign MUX_SB_T3_WEST_SB_OUT_B17_I[51+:17] = MEM_output_width_17_num_0;
	assign MUX_SB_T3_WEST_SB_OUT_B17_I[34+:17] = WIRE_SB_T3_EAST_SB_IN_B17_O;
	assign MUX_SB_T3_WEST_SB_OUT_B17_I[17+:17] = WIRE_SB_T2_SOUTH_SB_IN_B17_O;
	assign MUX_SB_T3_WEST_SB_OUT_B17_I[0+:17] = WIRE_SB_T2_NORTH_SB_IN_B17_O;
	wire [5:0] MUX_SB_T3_WEST_SB_OUT_B17_valid_in;
	assign MUX_SB_T3_WEST_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid, MEM_output_width_17_num_1_valid, MEM_output_width_17_num_0_valid, WIRE_SB_T3_EAST_SB_IN_B17_valid_out, WIRE_SB_T2_SOUTH_SB_IN_B17_valid_out, WIRE_SB_T2_NORTH_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_6_17 MUX_SB_T3_WEST_SB_OUT_B17(
		.I(MUX_SB_T3_WEST_SB_OUT_B17_I),
		.O(MUX_SB_T3_WEST_SB_OUT_B17_O),
		.ready_in(SB_T3_WEST_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T3_WEST_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T3_WEST_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T3_WEST_SB_OUT_B17_valid_out),
		.S(SB_T3_WEST_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T3_WEST_SB_OUT_B17_out_sel)
	);
	wire [101:0] MUX_SB_T4_EAST_SB_OUT_B17_I;
	assign MUX_SB_T4_EAST_SB_OUT_B17_I[85+:17] = MEM_output_width_17_num_2;
	assign MUX_SB_T4_EAST_SB_OUT_B17_I[68+:17] = MEM_output_width_17_num_1;
	assign MUX_SB_T4_EAST_SB_OUT_B17_I[51+:17] = MEM_output_width_17_num_0;
	assign MUX_SB_T4_EAST_SB_OUT_B17_I[34+:17] = WIRE_SB_T4_WEST_SB_IN_B17_O;
	assign MUX_SB_T4_EAST_SB_OUT_B17_I[17+:17] = WIRE_SB_T4_SOUTH_SB_IN_B17_O;
	assign MUX_SB_T4_EAST_SB_OUT_B17_I[0+:17] = WIRE_SB_T3_NORTH_SB_IN_B17_O;
	wire [5:0] MUX_SB_T4_EAST_SB_OUT_B17_valid_in;
	assign MUX_SB_T4_EAST_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid, MEM_output_width_17_num_1_valid, MEM_output_width_17_num_0_valid, WIRE_SB_T4_WEST_SB_IN_B17_valid_out, WIRE_SB_T4_SOUTH_SB_IN_B17_valid_out, WIRE_SB_T3_NORTH_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_6_17 MUX_SB_T4_EAST_SB_OUT_B17(
		.I(MUX_SB_T4_EAST_SB_OUT_B17_I),
		.O(MUX_SB_T4_EAST_SB_OUT_B17_O),
		.ready_in(SB_T4_EAST_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T4_EAST_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T4_EAST_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T4_EAST_SB_OUT_B17_valid_out),
		.S(SB_T4_EAST_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T4_EAST_SB_OUT_B17_out_sel)
	);
	wire [101:0] MUX_SB_T4_NORTH_SB_OUT_B17_I;
	assign MUX_SB_T4_NORTH_SB_OUT_B17_I[85+:17] = MEM_output_width_17_num_2;
	assign MUX_SB_T4_NORTH_SB_OUT_B17_I[68+:17] = MEM_output_width_17_num_1;
	assign MUX_SB_T4_NORTH_SB_OUT_B17_I[51+:17] = MEM_output_width_17_num_0;
	assign MUX_SB_T4_NORTH_SB_OUT_B17_I[34+:17] = WIRE_SB_T4_SOUTH_SB_IN_B17_O;
	assign MUX_SB_T4_NORTH_SB_OUT_B17_I[17+:17] = WIRE_SB_T0_EAST_SB_IN_B17_O;
	assign MUX_SB_T4_NORTH_SB_OUT_B17_I[0+:17] = WIRE_SB_T1_WEST_SB_IN_B17_O;
	wire [5:0] MUX_SB_T4_NORTH_SB_OUT_B17_valid_in;
	assign MUX_SB_T4_NORTH_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid, MEM_output_width_17_num_1_valid, MEM_output_width_17_num_0_valid, WIRE_SB_T4_SOUTH_SB_IN_B17_valid_out, WIRE_SB_T0_EAST_SB_IN_B17_valid_out, WIRE_SB_T1_WEST_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_6_17 MUX_SB_T4_NORTH_SB_OUT_B17(
		.I(MUX_SB_T4_NORTH_SB_OUT_B17_I),
		.O(MUX_SB_T4_NORTH_SB_OUT_B17_O),
		.ready_in(SB_T4_NORTH_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T4_NORTH_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T4_NORTH_SB_OUT_B17_valid_out),
		.S(SB_T4_NORTH_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel)
	);
	wire [101:0] MUX_SB_T4_SOUTH_SB_OUT_B17_I;
	assign MUX_SB_T4_SOUTH_SB_OUT_B17_I[85+:17] = MEM_output_width_17_num_2;
	assign MUX_SB_T4_SOUTH_SB_OUT_B17_I[68+:17] = MEM_output_width_17_num_1;
	assign MUX_SB_T4_SOUTH_SB_OUT_B17_I[51+:17] = MEM_output_width_17_num_0;
	assign MUX_SB_T4_SOUTH_SB_OUT_B17_I[34+:17] = WIRE_SB_T4_NORTH_SB_IN_B17_O;
	assign MUX_SB_T4_SOUTH_SB_OUT_B17_I[17+:17] = WIRE_SB_T4_EAST_SB_IN_B17_O;
	assign MUX_SB_T4_SOUTH_SB_OUT_B17_I[0+:17] = WIRE_SB_T0_WEST_SB_IN_B17_O;
	wire [5:0] MUX_SB_T4_SOUTH_SB_OUT_B17_valid_in;
	assign MUX_SB_T4_SOUTH_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid, MEM_output_width_17_num_1_valid, MEM_output_width_17_num_0_valid, WIRE_SB_T4_NORTH_SB_IN_B17_valid_out, WIRE_SB_T4_EAST_SB_IN_B17_valid_out, WIRE_SB_T0_WEST_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_6_17 MUX_SB_T4_SOUTH_SB_OUT_B17(
		.I(MUX_SB_T4_SOUTH_SB_OUT_B17_I),
		.O(MUX_SB_T4_SOUTH_SB_OUT_B17_O),
		.ready_in(SB_T4_SOUTH_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T4_SOUTH_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T4_SOUTH_SB_OUT_B17_valid_out),
		.S(SB_T4_SOUTH_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel)
	);
	wire [101:0] MUX_SB_T4_WEST_SB_OUT_B17_I;
	assign MUX_SB_T4_WEST_SB_OUT_B17_I[85+:17] = MEM_output_width_17_num_2;
	assign MUX_SB_T4_WEST_SB_OUT_B17_I[68+:17] = MEM_output_width_17_num_1;
	assign MUX_SB_T4_WEST_SB_OUT_B17_I[51+:17] = MEM_output_width_17_num_0;
	assign MUX_SB_T4_WEST_SB_OUT_B17_I[34+:17] = WIRE_SB_T4_EAST_SB_IN_B17_O;
	assign MUX_SB_T4_WEST_SB_OUT_B17_I[17+:17] = WIRE_SB_T3_SOUTH_SB_IN_B17_O;
	assign MUX_SB_T4_WEST_SB_OUT_B17_I[0+:17] = WIRE_SB_T1_NORTH_SB_IN_B17_O;
	wire [5:0] MUX_SB_T4_WEST_SB_OUT_B17_valid_in;
	assign MUX_SB_T4_WEST_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid, MEM_output_width_17_num_1_valid, MEM_output_width_17_num_0_valid, WIRE_SB_T4_EAST_SB_IN_B17_valid_out, WIRE_SB_T3_SOUTH_SB_IN_B17_valid_out, WIRE_SB_T1_NORTH_SB_IN_B17_valid_out};
	mux_aoi_ready_valid_6_17 MUX_SB_T4_WEST_SB_OUT_B17(
		.I(MUX_SB_T4_WEST_SB_OUT_B17_I),
		.O(MUX_SB_T4_WEST_SB_OUT_B17_O),
		.ready_in(SB_T4_WEST_SB_OUT_B17_FANOUT_O[0]),
		.ready_out(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
		.valid_in(MUX_SB_T4_WEST_SB_OUT_B17_valid_in),
		.valid_out(MUX_SB_T4_WEST_SB_OUT_B17_valid_out),
		.S(SB_T4_WEST_SB_OUT_B17_sel_value_O),
		.out_sel(MUX_SB_T4_WEST_SB_OUT_B17_out_sel)
	);
	SplitFifo_17 REG_T0_EAST_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T0_EAST_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T0_EAST_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T0_EAST_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T0_EAST_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst2_out[0]),
		.end_fifo(REG_T0_EAST_B17_end_value_O[0]),
		.valid0(MUX_SB_T0_EAST_SB_OUT_B17_valid_out),
		.valid1(REG_T0_EAST_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T0_EAST_B17_ready_out),
		.fifo_en(REG_T0_EAST_B17_fifo_value_O[0])
	);
	SliceWrapper_32_0_1 REG_T0_EAST_B17_end_value(
		.I(config_reg_0_O),
		.O(REG_T0_EAST_B17_end_value_O)
	);
	SliceWrapper_32_1_2 REG_T0_EAST_B17_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T0_EAST_B17_fifo_value_O)
	);
	SliceWrapper_32_2_3 REG_T0_EAST_B17_start_value(
		.I(config_reg_0_O),
		.O(REG_T0_EAST_B17_start_value_O)
	);
	SplitFifo_17 REG_T0_NORTH_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T0_NORTH_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T0_NORTH_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T0_NORTH_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T0_NORTH_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst0_out[0]),
		.end_fifo(REG_T0_NORTH_B17_end_value_O[0]),
		.valid0(MUX_SB_T0_NORTH_SB_OUT_B17_valid_out),
		.valid1(REG_T0_NORTH_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T0_NORTH_B17_ready_out),
		.fifo_en(REG_T0_NORTH_B17_fifo_value_O[0])
	);
	SliceWrapper_32_3_4 REG_T0_NORTH_B17_end_value(
		.I(config_reg_0_O),
		.O(REG_T0_NORTH_B17_end_value_O)
	);
	SliceWrapper_32_4_5 REG_T0_NORTH_B17_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T0_NORTH_B17_fifo_value_O)
	);
	SliceWrapper_32_5_6 REG_T0_NORTH_B17_start_value(
		.I(config_reg_0_O),
		.O(REG_T0_NORTH_B17_start_value_O)
	);
	SplitFifo_17 REG_T0_SOUTH_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T0_SOUTH_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T0_SOUTH_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T0_SOUTH_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T0_SOUTH_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst1_out[0]),
		.end_fifo(REG_T0_SOUTH_B17_end_value_O[0]),
		.valid0(MUX_SB_T0_SOUTH_SB_OUT_B17_valid_out),
		.valid1(REG_T0_SOUTH_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T0_SOUTH_B17_ready_out),
		.fifo_en(REG_T0_SOUTH_B17_fifo_value_O[0])
	);
	SliceWrapper_32_6_7 REG_T0_SOUTH_B17_end_value(
		.I(config_reg_0_O),
		.O(REG_T0_SOUTH_B17_end_value_O)
	);
	SliceWrapper_32_7_8 REG_T0_SOUTH_B17_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T0_SOUTH_B17_fifo_value_O)
	);
	SliceWrapper_32_8_9 REG_T0_SOUTH_B17_start_value(
		.I(config_reg_0_O),
		.O(REG_T0_SOUTH_B17_start_value_O)
	);
	SplitFifo_17 REG_T0_WEST_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T0_WEST_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T0_WEST_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T0_WEST_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T0_WEST_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst3_out[0]),
		.end_fifo(REG_T0_WEST_B17_end_value_O[0]),
		.valid0(MUX_SB_T0_WEST_SB_OUT_B17_valid_out),
		.valid1(REG_T0_WEST_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T0_WEST_B17_ready_out),
		.fifo_en(REG_T0_WEST_B17_fifo_value_O[0])
	);
	SliceWrapper_32_9_10 REG_T0_WEST_B17_end_value(
		.I(config_reg_0_O),
		.O(REG_T0_WEST_B17_end_value_O)
	);
	SliceWrapper_32_10_11 REG_T0_WEST_B17_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T0_WEST_B17_fifo_value_O)
	);
	SliceWrapper_32_11_12 REG_T0_WEST_B17_start_value(
		.I(config_reg_0_O),
		.O(REG_T0_WEST_B17_start_value_O)
	);
	SplitFifo_17 REG_T1_EAST_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T1_EAST_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T1_EAST_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T1_EAST_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T1_EAST_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst6_out[0]),
		.end_fifo(REG_T1_EAST_B17_end_value_O[0]),
		.valid0(MUX_SB_T1_EAST_SB_OUT_B17_valid_out),
		.valid1(REG_T1_EAST_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T1_EAST_B17_ready_out),
		.fifo_en(REG_T1_EAST_B17_fifo_value_O[0])
	);
	SliceWrapper_32_12_13 REG_T1_EAST_B17_end_value(
		.I(config_reg_0_O),
		.O(REG_T1_EAST_B17_end_value_O)
	);
	SliceWrapper_32_13_14 REG_T1_EAST_B17_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T1_EAST_B17_fifo_value_O)
	);
	SliceWrapper_32_14_15 REG_T1_EAST_B17_start_value(
		.I(config_reg_0_O),
		.O(REG_T1_EAST_B17_start_value_O)
	);
	SplitFifo_17 REG_T1_NORTH_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T1_NORTH_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T1_NORTH_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T1_NORTH_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T1_NORTH_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst4_out[0]),
		.end_fifo(REG_T1_NORTH_B17_end_value_O[0]),
		.valid0(MUX_SB_T1_NORTH_SB_OUT_B17_valid_out),
		.valid1(REG_T1_NORTH_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T1_NORTH_B17_ready_out),
		.fifo_en(REG_T1_NORTH_B17_fifo_value_O[0])
	);
	SliceWrapper_32_15_16 REG_T1_NORTH_B17_end_value(
		.I(config_reg_0_O),
		.O(REG_T1_NORTH_B17_end_value_O)
	);
	SliceWrapper_32_16_17 REG_T1_NORTH_B17_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T1_NORTH_B17_fifo_value_O)
	);
	SliceWrapper_32_17_18 REG_T1_NORTH_B17_start_value(
		.I(config_reg_0_O),
		.O(REG_T1_NORTH_B17_start_value_O)
	);
	SplitFifo_17 REG_T1_SOUTH_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T1_SOUTH_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T1_SOUTH_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T1_SOUTH_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T1_SOUTH_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst5_out[0]),
		.end_fifo(REG_T1_SOUTH_B17_end_value_O[0]),
		.valid0(MUX_SB_T1_SOUTH_SB_OUT_B17_valid_out),
		.valid1(REG_T1_SOUTH_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T1_SOUTH_B17_ready_out),
		.fifo_en(REG_T1_SOUTH_B17_fifo_value_O[0])
	);
	SliceWrapper_32_18_19 REG_T1_SOUTH_B17_end_value(
		.I(config_reg_0_O),
		.O(REG_T1_SOUTH_B17_end_value_O)
	);
	SliceWrapper_32_19_20 REG_T1_SOUTH_B17_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T1_SOUTH_B17_fifo_value_O)
	);
	SliceWrapper_32_20_21 REG_T1_SOUTH_B17_start_value(
		.I(config_reg_0_O),
		.O(REG_T1_SOUTH_B17_start_value_O)
	);
	SplitFifo_17 REG_T1_WEST_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T1_WEST_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T1_WEST_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T1_WEST_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T1_WEST_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst7_out[0]),
		.end_fifo(REG_T1_WEST_B17_end_value_O[0]),
		.valid0(MUX_SB_T1_WEST_SB_OUT_B17_valid_out),
		.valid1(REG_T1_WEST_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T1_WEST_B17_ready_out),
		.fifo_en(REG_T1_WEST_B17_fifo_value_O[0])
	);
	SliceWrapper_32_21_22 REG_T1_WEST_B17_end_value(
		.I(config_reg_0_O),
		.O(REG_T1_WEST_B17_end_value_O)
	);
	SliceWrapper_32_22_23 REG_T1_WEST_B17_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T1_WEST_B17_fifo_value_O)
	);
	SliceWrapper_32_23_24 REG_T1_WEST_B17_start_value(
		.I(config_reg_0_O),
		.O(REG_T1_WEST_B17_start_value_O)
	);
	SplitFifo_17 REG_T2_EAST_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T2_EAST_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T2_EAST_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T2_EAST_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T2_EAST_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst10_out[0]),
		.end_fifo(REG_T2_EAST_B17_end_value_O[0]),
		.valid0(MUX_SB_T2_EAST_SB_OUT_B17_valid_out),
		.valid1(REG_T2_EAST_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T2_EAST_B17_ready_out),
		.fifo_en(REG_T2_EAST_B17_fifo_value_O[0])
	);
	SliceWrapper_32_24_25 REG_T2_EAST_B17_end_value(
		.I(config_reg_0_O),
		.O(REG_T2_EAST_B17_end_value_O)
	);
	SliceWrapper_32_25_26 REG_T2_EAST_B17_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T2_EAST_B17_fifo_value_O)
	);
	SliceWrapper_32_26_27 REG_T2_EAST_B17_start_value(
		.I(config_reg_0_O),
		.O(REG_T2_EAST_B17_start_value_O)
	);
	SplitFifo_17 REG_T2_NORTH_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T2_NORTH_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T2_NORTH_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T2_NORTH_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T2_NORTH_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst8_out[0]),
		.end_fifo(REG_T2_NORTH_B17_end_value_O[0]),
		.valid0(MUX_SB_T2_NORTH_SB_OUT_B17_valid_out),
		.valid1(REG_T2_NORTH_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T2_NORTH_B17_ready_out),
		.fifo_en(REG_T2_NORTH_B17_fifo_value_O[0])
	);
	SliceWrapper_32_27_28 REG_T2_NORTH_B17_end_value(
		.I(config_reg_0_O),
		.O(REG_T2_NORTH_B17_end_value_O)
	);
	SliceWrapper_32_28_29 REG_T2_NORTH_B17_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T2_NORTH_B17_fifo_value_O)
	);
	SliceWrapper_32_29_30 REG_T2_NORTH_B17_start_value(
		.I(config_reg_0_O),
		.O(REG_T2_NORTH_B17_start_value_O)
	);
	SplitFifo_17 REG_T2_SOUTH_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T2_SOUTH_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T2_SOUTH_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T2_SOUTH_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T2_SOUTH_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst9_out[0]),
		.end_fifo(REG_T2_SOUTH_B17_end_value_O[0]),
		.valid0(MUX_SB_T2_SOUTH_SB_OUT_B17_valid_out),
		.valid1(REG_T2_SOUTH_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T2_SOUTH_B17_ready_out),
		.fifo_en(REG_T2_SOUTH_B17_fifo_value_O[0])
	);
	SliceWrapper_32_30_31 REG_T2_SOUTH_B17_end_value(
		.I(config_reg_0_O),
		.O(REG_T2_SOUTH_B17_end_value_O)
	);
	SliceWrapper_32_31_32 REG_T2_SOUTH_B17_fifo_value(
		.I(config_reg_0_O),
		.O(REG_T2_SOUTH_B17_fifo_value_O)
	);
	SliceWrapper_32_0_1 REG_T2_SOUTH_B17_start_value(
		.I(config_reg_1_O),
		.O(REG_T2_SOUTH_B17_start_value_O)
	);
	SplitFifo_17 REG_T2_WEST_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T2_WEST_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T2_WEST_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T2_WEST_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T2_WEST_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst11_out[0]),
		.end_fifo(REG_T2_WEST_B17_end_value_O[0]),
		.valid0(MUX_SB_T2_WEST_SB_OUT_B17_valid_out),
		.valid1(REG_T2_WEST_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T2_WEST_B17_ready_out),
		.fifo_en(REG_T2_WEST_B17_fifo_value_O[0])
	);
	SliceWrapper_32_1_2 REG_T2_WEST_B17_end_value(
		.I(config_reg_1_O),
		.O(REG_T2_WEST_B17_end_value_O)
	);
	SliceWrapper_32_2_3 REG_T2_WEST_B17_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T2_WEST_B17_fifo_value_O)
	);
	SliceWrapper_32_3_4 REG_T2_WEST_B17_start_value(
		.I(config_reg_1_O),
		.O(REG_T2_WEST_B17_start_value_O)
	);
	SplitFifo_17 REG_T3_EAST_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T3_EAST_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T3_EAST_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T3_EAST_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T3_EAST_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst14_out[0]),
		.end_fifo(REG_T3_EAST_B17_end_value_O[0]),
		.valid0(MUX_SB_T3_EAST_SB_OUT_B17_valid_out),
		.valid1(REG_T3_EAST_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T3_EAST_B17_ready_out),
		.fifo_en(REG_T3_EAST_B17_fifo_value_O[0])
	);
	SliceWrapper_32_4_5 REG_T3_EAST_B17_end_value(
		.I(config_reg_1_O),
		.O(REG_T3_EAST_B17_end_value_O)
	);
	SliceWrapper_32_5_6 REG_T3_EAST_B17_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T3_EAST_B17_fifo_value_O)
	);
	SliceWrapper_32_6_7 REG_T3_EAST_B17_start_value(
		.I(config_reg_1_O),
		.O(REG_T3_EAST_B17_start_value_O)
	);
	SplitFifo_17 REG_T3_NORTH_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T3_NORTH_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T3_NORTH_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T3_NORTH_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T3_NORTH_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst12_out[0]),
		.end_fifo(REG_T3_NORTH_B17_end_value_O[0]),
		.valid0(MUX_SB_T3_NORTH_SB_OUT_B17_valid_out),
		.valid1(REG_T3_NORTH_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T3_NORTH_B17_ready_out),
		.fifo_en(REG_T3_NORTH_B17_fifo_value_O[0])
	);
	SliceWrapper_32_7_8 REG_T3_NORTH_B17_end_value(
		.I(config_reg_1_O),
		.O(REG_T3_NORTH_B17_end_value_O)
	);
	SliceWrapper_32_8_9 REG_T3_NORTH_B17_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T3_NORTH_B17_fifo_value_O)
	);
	SliceWrapper_32_9_10 REG_T3_NORTH_B17_start_value(
		.I(config_reg_1_O),
		.O(REG_T3_NORTH_B17_start_value_O)
	);
	SplitFifo_17 REG_T3_SOUTH_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T3_SOUTH_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T3_SOUTH_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T3_SOUTH_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T3_SOUTH_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst13_out[0]),
		.end_fifo(REG_T3_SOUTH_B17_end_value_O[0]),
		.valid0(MUX_SB_T3_SOUTH_SB_OUT_B17_valid_out),
		.valid1(REG_T3_SOUTH_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T3_SOUTH_B17_ready_out),
		.fifo_en(REG_T3_SOUTH_B17_fifo_value_O[0])
	);
	SliceWrapper_32_10_11 REG_T3_SOUTH_B17_end_value(
		.I(config_reg_1_O),
		.O(REG_T3_SOUTH_B17_end_value_O)
	);
	SliceWrapper_32_11_12 REG_T3_SOUTH_B17_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T3_SOUTH_B17_fifo_value_O)
	);
	SliceWrapper_32_12_13 REG_T3_SOUTH_B17_start_value(
		.I(config_reg_1_O),
		.O(REG_T3_SOUTH_B17_start_value_O)
	);
	SplitFifo_17 REG_T3_WEST_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T3_WEST_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T3_WEST_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T3_WEST_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T3_WEST_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst15_out[0]),
		.end_fifo(REG_T3_WEST_B17_end_value_O[0]),
		.valid0(MUX_SB_T3_WEST_SB_OUT_B17_valid_out),
		.valid1(REG_T3_WEST_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T3_WEST_B17_ready_out),
		.fifo_en(REG_T3_WEST_B17_fifo_value_O[0])
	);
	SliceWrapper_32_13_14 REG_T3_WEST_B17_end_value(
		.I(config_reg_1_O),
		.O(REG_T3_WEST_B17_end_value_O)
	);
	SliceWrapper_32_14_15 REG_T3_WEST_B17_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T3_WEST_B17_fifo_value_O)
	);
	SliceWrapper_32_15_16 REG_T3_WEST_B17_start_value(
		.I(config_reg_1_O),
		.O(REG_T3_WEST_B17_start_value_O)
	);
	SplitFifo_17 REG_T4_EAST_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T4_EAST_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T4_EAST_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T4_EAST_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T4_EAST_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst18_out[0]),
		.end_fifo(REG_T4_EAST_B17_end_value_O[0]),
		.valid0(MUX_SB_T4_EAST_SB_OUT_B17_valid_out),
		.valid1(REG_T4_EAST_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T4_EAST_B17_ready_out),
		.fifo_en(REG_T4_EAST_B17_fifo_value_O[0])
	);
	SliceWrapper_32_16_17 REG_T4_EAST_B17_end_value(
		.I(config_reg_1_O),
		.O(REG_T4_EAST_B17_end_value_O)
	);
	SliceWrapper_32_17_18 REG_T4_EAST_B17_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T4_EAST_B17_fifo_value_O)
	);
	SliceWrapper_32_18_19 REG_T4_EAST_B17_start_value(
		.I(config_reg_1_O),
		.O(REG_T4_EAST_B17_start_value_O)
	);
	SplitFifo_17 REG_T4_NORTH_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T4_NORTH_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T4_NORTH_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T4_NORTH_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T4_NORTH_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst16_out[0]),
		.end_fifo(REG_T4_NORTH_B17_end_value_O[0]),
		.valid0(MUX_SB_T4_NORTH_SB_OUT_B17_valid_out),
		.valid1(REG_T4_NORTH_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T4_NORTH_B17_ready_out),
		.fifo_en(REG_T4_NORTH_B17_fifo_value_O[0])
	);
	SliceWrapper_32_19_20 REG_T4_NORTH_B17_end_value(
		.I(config_reg_1_O),
		.O(REG_T4_NORTH_B17_end_value_O)
	);
	SliceWrapper_32_20_21 REG_T4_NORTH_B17_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T4_NORTH_B17_fifo_value_O)
	);
	SliceWrapper_32_21_22 REG_T4_NORTH_B17_start_value(
		.I(config_reg_1_O),
		.O(REG_T4_NORTH_B17_start_value_O)
	);
	SplitFifo_17 REG_T4_SOUTH_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T4_SOUTH_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T4_SOUTH_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T4_SOUTH_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T4_SOUTH_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst17_out[0]),
		.end_fifo(REG_T4_SOUTH_B17_end_value_O[0]),
		.valid0(MUX_SB_T4_SOUTH_SB_OUT_B17_valid_out),
		.valid1(REG_T4_SOUTH_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T4_SOUTH_B17_ready_out),
		.fifo_en(REG_T4_SOUTH_B17_fifo_value_O[0])
	);
	SliceWrapper_32_22_23 REG_T4_SOUTH_B17_end_value(
		.I(config_reg_1_O),
		.O(REG_T4_SOUTH_B17_end_value_O)
	);
	SliceWrapper_32_23_24 REG_T4_SOUTH_B17_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T4_SOUTH_B17_fifo_value_O)
	);
	SliceWrapper_32_24_25 REG_T4_SOUTH_B17_start_value(
		.I(config_reg_1_O),
		.O(REG_T4_SOUTH_B17_start_value_O)
	);
	SplitFifo_17 REG_T4_WEST_B17$SplitFifo_17_inst0(
		.data_in(MUX_SB_T4_WEST_SB_OUT_B17_O),
		.rst(reset),
		.start_fifo(REG_T4_WEST_B17_start_value_O[0]),
		.clk(clk),
		.ready0(REG_T4_WEST_B17$SplitFifo_17_inst0_ready0),
		.data_out(REG_T4_WEST_B17$SplitFifo_17_inst0_data_out),
		.clk_en(and1_inst19_out[0]),
		.end_fifo(REG_T4_WEST_B17_end_value_O[0]),
		.valid0(MUX_SB_T4_WEST_SB_OUT_B17_valid_out),
		.valid1(REG_T4_WEST_B17$SplitFifo_17_inst0_valid1),
		.ready1(RMUX_T4_WEST_B17_ready_out),
		.fifo_en(REG_T4_WEST_B17_fifo_value_O[0])
	);
	SliceWrapper_32_25_26 REG_T4_WEST_B17_end_value(
		.I(config_reg_1_O),
		.O(REG_T4_WEST_B17_end_value_O)
	);
	SliceWrapper_32_26_27 REG_T4_WEST_B17_fifo_value(
		.I(config_reg_1_O),
		.O(REG_T4_WEST_B17_fifo_value_O)
	);
	SliceWrapper_32_27_28 REG_T4_WEST_B17_start_value(
		.I(config_reg_1_O),
		.O(REG_T4_WEST_B17_start_value_O)
	);
	wire [33:0] RMUX_T0_EAST_B17_I;
	assign RMUX_T0_EAST_B17_I[17+:17] = REG_T0_EAST_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T0_EAST_B17_I[0+:17] = MUX_SB_T0_EAST_SB_OUT_B17_O;
	wire [1:0] RMUX_T0_EAST_B17_valid_in;
	assign RMUX_T0_EAST_B17_valid_in = {REG_T0_EAST_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T0_EAST_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T0_EAST_B17(
		.I(RMUX_T0_EAST_B17_I),
		.O(RMUX_T0_EAST_B17_O),
		.ready_in(SB_T0_EAST_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T0_EAST_B17_ready_out),
		.valid_in(RMUX_T0_EAST_B17_valid_in),
		.valid_out(RMUX_T0_EAST_B17_valid_out),
		.S(RMUX_T0_EAST_B17_sel_value_O),
		.out_sel(RMUX_T0_EAST_B17_out_sel)
	);
	SliceWrapper_32_28_29 RMUX_T0_EAST_B17_sel_value(
		.I(config_reg_1_O),
		.O(RMUX_T0_EAST_B17_sel_value_O)
	);
	wire [33:0] RMUX_T0_NORTH_B17_I;
	assign RMUX_T0_NORTH_B17_I[17+:17] = REG_T0_NORTH_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T0_NORTH_B17_I[0+:17] = MUX_SB_T0_NORTH_SB_OUT_B17_O;
	wire [1:0] RMUX_T0_NORTH_B17_valid_in;
	assign RMUX_T0_NORTH_B17_valid_in = {REG_T0_NORTH_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T0_NORTH_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T0_NORTH_B17(
		.I(RMUX_T0_NORTH_B17_I),
		.O(RMUX_T0_NORTH_B17_O),
		.ready_in(SB_T0_NORTH_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T0_NORTH_B17_ready_out),
		.valid_in(RMUX_T0_NORTH_B17_valid_in),
		.valid_out(RMUX_T0_NORTH_B17_valid_out),
		.S(RMUX_T0_NORTH_B17_sel_value_O),
		.out_sel(RMUX_T0_NORTH_B17_out_sel)
	);
	SliceWrapper_32_29_30 RMUX_T0_NORTH_B17_sel_value(
		.I(config_reg_1_O),
		.O(RMUX_T0_NORTH_B17_sel_value_O)
	);
	wire [33:0] RMUX_T0_SOUTH_B17_I;
	assign RMUX_T0_SOUTH_B17_I[17+:17] = REG_T0_SOUTH_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T0_SOUTH_B17_I[0+:17] = MUX_SB_T0_SOUTH_SB_OUT_B17_O;
	wire [1:0] RMUX_T0_SOUTH_B17_valid_in;
	assign RMUX_T0_SOUTH_B17_valid_in = {REG_T0_SOUTH_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T0_SOUTH_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T0_SOUTH_B17(
		.I(RMUX_T0_SOUTH_B17_I),
		.O(RMUX_T0_SOUTH_B17_O),
		.ready_in(SB_T0_SOUTH_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T0_SOUTH_B17_ready_out),
		.valid_in(RMUX_T0_SOUTH_B17_valid_in),
		.valid_out(RMUX_T0_SOUTH_B17_valid_out),
		.S(RMUX_T0_SOUTH_B17_sel_value_O),
		.out_sel(RMUX_T0_SOUTH_B17_out_sel)
	);
	SliceWrapper_32_30_31 RMUX_T0_SOUTH_B17_sel_value(
		.I(config_reg_1_O),
		.O(RMUX_T0_SOUTH_B17_sel_value_O)
	);
	wire [33:0] RMUX_T0_WEST_B17_I;
	assign RMUX_T0_WEST_B17_I[17+:17] = REG_T0_WEST_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T0_WEST_B17_I[0+:17] = MUX_SB_T0_WEST_SB_OUT_B17_O;
	wire [1:0] RMUX_T0_WEST_B17_valid_in;
	assign RMUX_T0_WEST_B17_valid_in = {REG_T0_WEST_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T0_WEST_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T0_WEST_B17(
		.I(RMUX_T0_WEST_B17_I),
		.O(RMUX_T0_WEST_B17_O),
		.ready_in(SB_T0_WEST_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T0_WEST_B17_ready_out),
		.valid_in(RMUX_T0_WEST_B17_valid_in),
		.valid_out(RMUX_T0_WEST_B17_valid_out),
		.S(RMUX_T0_WEST_B17_sel_value_O),
		.out_sel(RMUX_T0_WEST_B17_out_sel)
	);
	SliceWrapper_32_31_32 RMUX_T0_WEST_B17_sel_value(
		.I(config_reg_1_O),
		.O(RMUX_T0_WEST_B17_sel_value_O)
	);
	wire [33:0] RMUX_T1_EAST_B17_I;
	assign RMUX_T1_EAST_B17_I[17+:17] = REG_T1_EAST_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T1_EAST_B17_I[0+:17] = MUX_SB_T1_EAST_SB_OUT_B17_O;
	wire [1:0] RMUX_T1_EAST_B17_valid_in;
	assign RMUX_T1_EAST_B17_valid_in = {REG_T1_EAST_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T1_EAST_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T1_EAST_B17(
		.I(RMUX_T1_EAST_B17_I),
		.O(RMUX_T1_EAST_B17_O),
		.ready_in(SB_T1_EAST_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T1_EAST_B17_ready_out),
		.valid_in(RMUX_T1_EAST_B17_valid_in),
		.valid_out(RMUX_T1_EAST_B17_valid_out),
		.S(RMUX_T1_EAST_B17_sel_value_O),
		.out_sel(RMUX_T1_EAST_B17_out_sel)
	);
	SliceWrapper_32_0_1 RMUX_T1_EAST_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T1_EAST_B17_sel_value_O)
	);
	wire [33:0] RMUX_T1_NORTH_B17_I;
	assign RMUX_T1_NORTH_B17_I[17+:17] = REG_T1_NORTH_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T1_NORTH_B17_I[0+:17] = MUX_SB_T1_NORTH_SB_OUT_B17_O;
	wire [1:0] RMUX_T1_NORTH_B17_valid_in;
	assign RMUX_T1_NORTH_B17_valid_in = {REG_T1_NORTH_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T1_NORTH_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T1_NORTH_B17(
		.I(RMUX_T1_NORTH_B17_I),
		.O(RMUX_T1_NORTH_B17_O),
		.ready_in(SB_T1_NORTH_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T1_NORTH_B17_ready_out),
		.valid_in(RMUX_T1_NORTH_B17_valid_in),
		.valid_out(RMUX_T1_NORTH_B17_valid_out),
		.S(RMUX_T1_NORTH_B17_sel_value_O),
		.out_sel(RMUX_T1_NORTH_B17_out_sel)
	);
	SliceWrapper_32_1_2 RMUX_T1_NORTH_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T1_NORTH_B17_sel_value_O)
	);
	wire [33:0] RMUX_T1_SOUTH_B17_I;
	assign RMUX_T1_SOUTH_B17_I[17+:17] = REG_T1_SOUTH_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T1_SOUTH_B17_I[0+:17] = MUX_SB_T1_SOUTH_SB_OUT_B17_O;
	wire [1:0] RMUX_T1_SOUTH_B17_valid_in;
	assign RMUX_T1_SOUTH_B17_valid_in = {REG_T1_SOUTH_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T1_SOUTH_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T1_SOUTH_B17(
		.I(RMUX_T1_SOUTH_B17_I),
		.O(RMUX_T1_SOUTH_B17_O),
		.ready_in(SB_T1_SOUTH_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T1_SOUTH_B17_ready_out),
		.valid_in(RMUX_T1_SOUTH_B17_valid_in),
		.valid_out(RMUX_T1_SOUTH_B17_valid_out),
		.S(RMUX_T1_SOUTH_B17_sel_value_O),
		.out_sel(RMUX_T1_SOUTH_B17_out_sel)
	);
	SliceWrapper_32_2_3 RMUX_T1_SOUTH_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T1_SOUTH_B17_sel_value_O)
	);
	wire [33:0] RMUX_T1_WEST_B17_I;
	assign RMUX_T1_WEST_B17_I[17+:17] = REG_T1_WEST_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T1_WEST_B17_I[0+:17] = MUX_SB_T1_WEST_SB_OUT_B17_O;
	wire [1:0] RMUX_T1_WEST_B17_valid_in;
	assign RMUX_T1_WEST_B17_valid_in = {REG_T1_WEST_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T1_WEST_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T1_WEST_B17(
		.I(RMUX_T1_WEST_B17_I),
		.O(RMUX_T1_WEST_B17_O),
		.ready_in(SB_T1_WEST_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T1_WEST_B17_ready_out),
		.valid_in(RMUX_T1_WEST_B17_valid_in),
		.valid_out(RMUX_T1_WEST_B17_valid_out),
		.S(RMUX_T1_WEST_B17_sel_value_O),
		.out_sel(RMUX_T1_WEST_B17_out_sel)
	);
	SliceWrapper_32_3_4 RMUX_T1_WEST_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T1_WEST_B17_sel_value_O)
	);
	wire [33:0] RMUX_T2_EAST_B17_I;
	assign RMUX_T2_EAST_B17_I[17+:17] = REG_T2_EAST_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T2_EAST_B17_I[0+:17] = MUX_SB_T2_EAST_SB_OUT_B17_O;
	wire [1:0] RMUX_T2_EAST_B17_valid_in;
	assign RMUX_T2_EAST_B17_valid_in = {REG_T2_EAST_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T2_EAST_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T2_EAST_B17(
		.I(RMUX_T2_EAST_B17_I),
		.O(RMUX_T2_EAST_B17_O),
		.ready_in(SB_T2_EAST_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T2_EAST_B17_ready_out),
		.valid_in(RMUX_T2_EAST_B17_valid_in),
		.valid_out(RMUX_T2_EAST_B17_valid_out),
		.S(RMUX_T2_EAST_B17_sel_value_O),
		.out_sel(RMUX_T2_EAST_B17_out_sel)
	);
	SliceWrapper_32_4_5 RMUX_T2_EAST_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T2_EAST_B17_sel_value_O)
	);
	wire [33:0] RMUX_T2_NORTH_B17_I;
	assign RMUX_T2_NORTH_B17_I[17+:17] = REG_T2_NORTH_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T2_NORTH_B17_I[0+:17] = MUX_SB_T2_NORTH_SB_OUT_B17_O;
	wire [1:0] RMUX_T2_NORTH_B17_valid_in;
	assign RMUX_T2_NORTH_B17_valid_in = {REG_T2_NORTH_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T2_NORTH_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T2_NORTH_B17(
		.I(RMUX_T2_NORTH_B17_I),
		.O(RMUX_T2_NORTH_B17_O),
		.ready_in(SB_T2_NORTH_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T2_NORTH_B17_ready_out),
		.valid_in(RMUX_T2_NORTH_B17_valid_in),
		.valid_out(RMUX_T2_NORTH_B17_valid_out),
		.S(RMUX_T2_NORTH_B17_sel_value_O),
		.out_sel(RMUX_T2_NORTH_B17_out_sel)
	);
	SliceWrapper_32_5_6 RMUX_T2_NORTH_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T2_NORTH_B17_sel_value_O)
	);
	wire [33:0] RMUX_T2_SOUTH_B17_I;
	assign RMUX_T2_SOUTH_B17_I[17+:17] = REG_T2_SOUTH_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T2_SOUTH_B17_I[0+:17] = MUX_SB_T2_SOUTH_SB_OUT_B17_O;
	wire [1:0] RMUX_T2_SOUTH_B17_valid_in;
	assign RMUX_T2_SOUTH_B17_valid_in = {REG_T2_SOUTH_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T2_SOUTH_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T2_SOUTH_B17(
		.I(RMUX_T2_SOUTH_B17_I),
		.O(RMUX_T2_SOUTH_B17_O),
		.ready_in(SB_T2_SOUTH_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T2_SOUTH_B17_ready_out),
		.valid_in(RMUX_T2_SOUTH_B17_valid_in),
		.valid_out(RMUX_T2_SOUTH_B17_valid_out),
		.S(RMUX_T2_SOUTH_B17_sel_value_O),
		.out_sel(RMUX_T2_SOUTH_B17_out_sel)
	);
	SliceWrapper_32_6_7 RMUX_T2_SOUTH_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T2_SOUTH_B17_sel_value_O)
	);
	wire [33:0] RMUX_T2_WEST_B17_I;
	assign RMUX_T2_WEST_B17_I[17+:17] = REG_T2_WEST_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T2_WEST_B17_I[0+:17] = MUX_SB_T2_WEST_SB_OUT_B17_O;
	wire [1:0] RMUX_T2_WEST_B17_valid_in;
	assign RMUX_T2_WEST_B17_valid_in = {REG_T2_WEST_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T2_WEST_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T2_WEST_B17(
		.I(RMUX_T2_WEST_B17_I),
		.O(RMUX_T2_WEST_B17_O),
		.ready_in(SB_T2_WEST_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T2_WEST_B17_ready_out),
		.valid_in(RMUX_T2_WEST_B17_valid_in),
		.valid_out(RMUX_T2_WEST_B17_valid_out),
		.S(RMUX_T2_WEST_B17_sel_value_O),
		.out_sel(RMUX_T2_WEST_B17_out_sel)
	);
	SliceWrapper_32_7_8 RMUX_T2_WEST_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T2_WEST_B17_sel_value_O)
	);
	wire [33:0] RMUX_T3_EAST_B17_I;
	assign RMUX_T3_EAST_B17_I[17+:17] = REG_T3_EAST_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T3_EAST_B17_I[0+:17] = MUX_SB_T3_EAST_SB_OUT_B17_O;
	wire [1:0] RMUX_T3_EAST_B17_valid_in;
	assign RMUX_T3_EAST_B17_valid_in = {REG_T3_EAST_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T3_EAST_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T3_EAST_B17(
		.I(RMUX_T3_EAST_B17_I),
		.O(RMUX_T3_EAST_B17_O),
		.ready_in(SB_T3_EAST_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T3_EAST_B17_ready_out),
		.valid_in(RMUX_T3_EAST_B17_valid_in),
		.valid_out(RMUX_T3_EAST_B17_valid_out),
		.S(RMUX_T3_EAST_B17_sel_value_O),
		.out_sel(RMUX_T3_EAST_B17_out_sel)
	);
	SliceWrapper_32_8_9 RMUX_T3_EAST_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T3_EAST_B17_sel_value_O)
	);
	wire [33:0] RMUX_T3_NORTH_B17_I;
	assign RMUX_T3_NORTH_B17_I[17+:17] = REG_T3_NORTH_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T3_NORTH_B17_I[0+:17] = MUX_SB_T3_NORTH_SB_OUT_B17_O;
	wire [1:0] RMUX_T3_NORTH_B17_valid_in;
	assign RMUX_T3_NORTH_B17_valid_in = {REG_T3_NORTH_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T3_NORTH_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T3_NORTH_B17(
		.I(RMUX_T3_NORTH_B17_I),
		.O(RMUX_T3_NORTH_B17_O),
		.ready_in(SB_T3_NORTH_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T3_NORTH_B17_ready_out),
		.valid_in(RMUX_T3_NORTH_B17_valid_in),
		.valid_out(RMUX_T3_NORTH_B17_valid_out),
		.S(RMUX_T3_NORTH_B17_sel_value_O),
		.out_sel(RMUX_T3_NORTH_B17_out_sel)
	);
	SliceWrapper_32_9_10 RMUX_T3_NORTH_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T3_NORTH_B17_sel_value_O)
	);
	wire [33:0] RMUX_T3_SOUTH_B17_I;
	assign RMUX_T3_SOUTH_B17_I[17+:17] = REG_T3_SOUTH_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T3_SOUTH_B17_I[0+:17] = MUX_SB_T3_SOUTH_SB_OUT_B17_O;
	wire [1:0] RMUX_T3_SOUTH_B17_valid_in;
	assign RMUX_T3_SOUTH_B17_valid_in = {REG_T3_SOUTH_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T3_SOUTH_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T3_SOUTH_B17(
		.I(RMUX_T3_SOUTH_B17_I),
		.O(RMUX_T3_SOUTH_B17_O),
		.ready_in(SB_T3_SOUTH_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T3_SOUTH_B17_ready_out),
		.valid_in(RMUX_T3_SOUTH_B17_valid_in),
		.valid_out(RMUX_T3_SOUTH_B17_valid_out),
		.S(RMUX_T3_SOUTH_B17_sel_value_O),
		.out_sel(RMUX_T3_SOUTH_B17_out_sel)
	);
	SliceWrapper_32_10_11 RMUX_T3_SOUTH_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T3_SOUTH_B17_sel_value_O)
	);
	wire [33:0] RMUX_T3_WEST_B17_I;
	assign RMUX_T3_WEST_B17_I[17+:17] = REG_T3_WEST_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T3_WEST_B17_I[0+:17] = MUX_SB_T3_WEST_SB_OUT_B17_O;
	wire [1:0] RMUX_T3_WEST_B17_valid_in;
	assign RMUX_T3_WEST_B17_valid_in = {REG_T3_WEST_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T3_WEST_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T3_WEST_B17(
		.I(RMUX_T3_WEST_B17_I),
		.O(RMUX_T3_WEST_B17_O),
		.ready_in(SB_T3_WEST_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T3_WEST_B17_ready_out),
		.valid_in(RMUX_T3_WEST_B17_valid_in),
		.valid_out(RMUX_T3_WEST_B17_valid_out),
		.S(RMUX_T3_WEST_B17_sel_value_O),
		.out_sel(RMUX_T3_WEST_B17_out_sel)
	);
	SliceWrapper_32_11_12 RMUX_T3_WEST_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T3_WEST_B17_sel_value_O)
	);
	wire [33:0] RMUX_T4_EAST_B17_I;
	assign RMUX_T4_EAST_B17_I[17+:17] = REG_T4_EAST_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T4_EAST_B17_I[0+:17] = MUX_SB_T4_EAST_SB_OUT_B17_O;
	wire [1:0] RMUX_T4_EAST_B17_valid_in;
	assign RMUX_T4_EAST_B17_valid_in = {REG_T4_EAST_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T4_EAST_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T4_EAST_B17(
		.I(RMUX_T4_EAST_B17_I),
		.O(RMUX_T4_EAST_B17_O),
		.ready_in(SB_T4_EAST_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T4_EAST_B17_ready_out),
		.valid_in(RMUX_T4_EAST_B17_valid_in),
		.valid_out(RMUX_T4_EAST_B17_valid_out),
		.S(RMUX_T4_EAST_B17_sel_value_O),
		.out_sel(RMUX_T4_EAST_B17_out_sel)
	);
	SliceWrapper_32_12_13 RMUX_T4_EAST_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T4_EAST_B17_sel_value_O)
	);
	wire [33:0] RMUX_T4_NORTH_B17_I;
	assign RMUX_T4_NORTH_B17_I[17+:17] = REG_T4_NORTH_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T4_NORTH_B17_I[0+:17] = MUX_SB_T4_NORTH_SB_OUT_B17_O;
	wire [1:0] RMUX_T4_NORTH_B17_valid_in;
	assign RMUX_T4_NORTH_B17_valid_in = {REG_T4_NORTH_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T4_NORTH_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T4_NORTH_B17(
		.I(RMUX_T4_NORTH_B17_I),
		.O(RMUX_T4_NORTH_B17_O),
		.ready_in(SB_T4_NORTH_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T4_NORTH_B17_ready_out),
		.valid_in(RMUX_T4_NORTH_B17_valid_in),
		.valid_out(RMUX_T4_NORTH_B17_valid_out),
		.S(RMUX_T4_NORTH_B17_sel_value_O),
		.out_sel(RMUX_T4_NORTH_B17_out_sel)
	);
	SliceWrapper_32_13_14 RMUX_T4_NORTH_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T4_NORTH_B17_sel_value_O)
	);
	wire [33:0] RMUX_T4_SOUTH_B17_I;
	assign RMUX_T4_SOUTH_B17_I[17+:17] = REG_T4_SOUTH_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T4_SOUTH_B17_I[0+:17] = MUX_SB_T4_SOUTH_SB_OUT_B17_O;
	wire [1:0] RMUX_T4_SOUTH_B17_valid_in;
	assign RMUX_T4_SOUTH_B17_valid_in = {REG_T4_SOUTH_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T4_SOUTH_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T4_SOUTH_B17(
		.I(RMUX_T4_SOUTH_B17_I),
		.O(RMUX_T4_SOUTH_B17_O),
		.ready_in(SB_T4_SOUTH_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T4_SOUTH_B17_ready_out),
		.valid_in(RMUX_T4_SOUTH_B17_valid_in),
		.valid_out(RMUX_T4_SOUTH_B17_valid_out),
		.S(RMUX_T4_SOUTH_B17_sel_value_O),
		.out_sel(RMUX_T4_SOUTH_B17_out_sel)
	);
	SliceWrapper_32_14_15 RMUX_T4_SOUTH_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T4_SOUTH_B17_sel_value_O)
	);
	wire [33:0] RMUX_T4_WEST_B17_I;
	assign RMUX_T4_WEST_B17_I[17+:17] = REG_T4_WEST_B17$SplitFifo_17_inst0_data_out;
	assign RMUX_T4_WEST_B17_I[0+:17] = MUX_SB_T4_WEST_SB_OUT_B17_O;
	wire [1:0] RMUX_T4_WEST_B17_valid_in;
	assign RMUX_T4_WEST_B17_valid_in = {REG_T4_WEST_B17$SplitFifo_17_inst0_valid1[0], MUX_SB_T4_WEST_SB_OUT_B17_valid_out};
	mux_aoi_ready_valid_2_17 RMUX_T4_WEST_B17(
		.I(RMUX_T4_WEST_B17_I),
		.O(RMUX_T4_WEST_B17_O),
		.ready_in(SB_T4_WEST_SB_OUT_B17_ready_in),
		.ready_out(RMUX_T4_WEST_B17_ready_out),
		.valid_in(RMUX_T4_WEST_B17_valid_in),
		.valid_out(RMUX_T4_WEST_B17_valid_out),
		.S(RMUX_T4_WEST_B17_sel_value_O),
		.out_sel(RMUX_T4_WEST_B17_out_sel)
	);
	SliceWrapper_32_15_16 RMUX_T4_WEST_B17_sel_value(
		.I(config_reg_2_O),
		.O(RMUX_T4_WEST_B17_sel_value_O)
	);
	SliceWrapper_32_16_17 SB_T0_EAST_SB_IN_B17_enable_value(
		.I(config_reg_2_O),
		.O(SB_T0_EAST_SB_IN_B17_enable_value_O)
	);
	FanoutHash_302974B49BE3F0C4 SB_T0_EAST_SB_IN_B17_fan_in(
		.E6(MEM_input_width_17_num_3_enable),
		.E3(MEM_input_width_17_num_0_enable),
		.I5(MEM_input_width_17_num_2_ready),
		.S6(MEM_input_width_17_num_3_out_sel),
		.E0(SB_T0_WEST_SB_OUT_B17_enable_value_O),
		.S5(MEM_input_width_17_num_2_out_sel),
		.I6(MEM_input_width_17_num_3_ready),
		.S3(MEM_input_width_17_num_0_out_sel),
		.S4(MEM_input_width_17_num_1_out_sel),
		.I3(MEM_input_width_17_num_0_ready),
		.I4(MEM_input_width_17_num_1_ready),
		.S1(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T0_WEST_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel),
		.E2(SB_T4_NORTH_SB_OUT_B17_enable_value_O),
		.E5(MEM_input_width_17_num_2_enable),
		.E4(MEM_input_width_17_num_1_enable),
		.I2(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
		.O(SB_T0_EAST_SB_IN_B17_fan_in_O),
		.E1(SB_T3_SOUTH_SB_OUT_B17_enable_value_O),
		.I0(MUX_SB_T0_WEST_SB_OUT_B17_ready_out)
	);
	wire [1:0] SB_T0_EAST_SB_OUT_B17_FANOUT_I;
	assign SB_T0_EAST_SB_OUT_B17_FANOUT_I = {REG_T0_EAST_B17$SplitFifo_17_inst0_ready0[0], RMUX_T0_EAST_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T0_EAST_SB_OUT_B17_FANOUT(
		.O(SB_T0_EAST_SB_OUT_B17_FANOUT_O),
		.I(SB_T0_EAST_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T0_EAST_B17_out_sel)
	);
	SliceWrapper_32_17_18 SB_T0_EAST_SB_OUT_B17_enable_value(
		.I(config_reg_2_O),
		.O(SB_T0_EAST_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_32_18_21 SB_T0_EAST_SB_OUT_B17_sel_value(
		.I(config_reg_2_O),
		.O(SB_T0_EAST_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_32_21_22 SB_T0_NORTH_SB_IN_B17_enable_value(
		.I(config_reg_2_O),
		.O(SB_T0_NORTH_SB_IN_B17_enable_value_O)
	);
	FanoutHash_47712AAC902ADA2 SB_T0_NORTH_SB_IN_B17_fan_in(
		.E6(MEM_input_width_17_num_3_enable),
		.E3(MEM_input_width_17_num_0_enable),
		.I5(MEM_input_width_17_num_2_ready),
		.S6(MEM_input_width_17_num_3_out_sel),
		.E0(SB_T0_WEST_SB_OUT_B17_enable_value_O),
		.S5(MEM_input_width_17_num_2_out_sel),
		.I6(MEM_input_width_17_num_3_ready),
		.S3(MEM_input_width_17_num_0_out_sel),
		.S4(MEM_input_width_17_num_1_out_sel),
		.I3(MEM_input_width_17_num_0_ready),
		.I4(MEM_input_width_17_num_1_ready),
		.S1(MUX_SB_T1_EAST_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T0_WEST_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel),
		.E2(SB_T0_SOUTH_SB_OUT_B17_enable_value_O),
		.E5(MEM_input_width_17_num_2_enable),
		.E4(MEM_input_width_17_num_1_enable),
		.I2(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
		.O(SB_T0_NORTH_SB_IN_B17_fan_in_O),
		.E1(SB_T1_EAST_SB_OUT_B17_enable_value_O),
		.I0(MUX_SB_T0_WEST_SB_OUT_B17_ready_out)
	);
	wire [1:0] SB_T0_NORTH_SB_OUT_B17_FANOUT_I;
	assign SB_T0_NORTH_SB_OUT_B17_FANOUT_I = {REG_T0_NORTH_B17$SplitFifo_17_inst0_ready0[0], RMUX_T0_NORTH_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T0_NORTH_SB_OUT_B17_FANOUT(
		.O(SB_T0_NORTH_SB_OUT_B17_FANOUT_O),
		.I(SB_T0_NORTH_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T0_NORTH_B17_out_sel)
	);
	SliceWrapper_32_22_23 SB_T0_NORTH_SB_OUT_B17_enable_value(
		.I(config_reg_2_O),
		.O(SB_T0_NORTH_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_32_23_26 SB_T0_NORTH_SB_OUT_B17_sel_value(
		.I(config_reg_2_O),
		.O(SB_T0_NORTH_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_32_26_27 SB_T0_SOUTH_SB_IN_B17_enable_value(
		.I(config_reg_2_O),
		.O(SB_T0_SOUTH_SB_IN_B17_enable_value_O)
	);
	FanoutHash_2785CE916183C5C SB_T0_SOUTH_SB_IN_B17_fan_in(
		.E6(MEM_input_width_17_num_3_enable),
		.E3(MEM_input_width_17_num_0_enable),
		.I5(MEM_input_width_17_num_2_ready),
		.S6(MEM_input_width_17_num_3_out_sel),
		.E0(SB_T3_EAST_SB_OUT_B17_enable_value_O),
		.S5(MEM_input_width_17_num_2_out_sel),
		.I6(MEM_input_width_17_num_3_ready),
		.S3(MEM_input_width_17_num_0_out_sel),
		.S4(MEM_input_width_17_num_1_out_sel),
		.I3(MEM_input_width_17_num_0_ready),
		.I4(MEM_input_width_17_num_1_ready),
		.S1(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T3_EAST_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T1_WEST_SB_OUT_B17_out_sel),
		.E2(SB_T1_WEST_SB_OUT_B17_enable_value_O),
		.E5(MEM_input_width_17_num_2_enable),
		.E4(MEM_input_width_17_num_1_enable),
		.I2(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out),
		.O(SB_T0_SOUTH_SB_IN_B17_fan_in_O),
		.E1(SB_T0_NORTH_SB_OUT_B17_enable_value_O),
		.I0(MUX_SB_T3_EAST_SB_OUT_B17_ready_out)
	);
	wire [1:0] SB_T0_SOUTH_SB_OUT_B17_FANOUT_I;
	assign SB_T0_SOUTH_SB_OUT_B17_FANOUT_I = {REG_T0_SOUTH_B17$SplitFifo_17_inst0_ready0[0], RMUX_T0_SOUTH_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T0_SOUTH_SB_OUT_B17_FANOUT(
		.O(SB_T0_SOUTH_SB_OUT_B17_FANOUT_O),
		.I(SB_T0_SOUTH_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T0_SOUTH_B17_out_sel)
	);
	SliceWrapper_32_27_28 SB_T0_SOUTH_SB_OUT_B17_enable_value(
		.I(config_reg_2_O),
		.O(SB_T0_SOUTH_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_32_28_31 SB_T0_SOUTH_SB_OUT_B17_sel_value(
		.I(config_reg_2_O),
		.O(SB_T0_SOUTH_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_32_31_32 SB_T0_WEST_SB_IN_B17_enable_value(
		.I(config_reg_2_O),
		.O(SB_T0_WEST_SB_IN_B17_enable_value_O)
	);
	FanoutHash_65A468071775C7BB SB_T0_WEST_SB_IN_B17_fan_in(
		.E6(MEM_input_width_17_num_3_enable),
		.E3(MEM_input_width_17_num_0_enable),
		.I5(MEM_input_width_17_num_2_ready),
		.S6(MEM_input_width_17_num_3_out_sel),
		.E0(SB_T0_NORTH_SB_OUT_B17_enable_value_O),
		.S5(MEM_input_width_17_num_2_out_sel),
		.I6(MEM_input_width_17_num_3_ready),
		.S3(MEM_input_width_17_num_0_out_sel),
		.S4(MEM_input_width_17_num_1_out_sel),
		.I3(MEM_input_width_17_num_0_ready),
		.I4(MEM_input_width_17_num_1_ready),
		.S1(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T0_EAST_SB_OUT_B17_out_sel),
		.E2(SB_T0_EAST_SB_OUT_B17_enable_value_O),
		.E5(MEM_input_width_17_num_2_enable),
		.E4(MEM_input_width_17_num_1_enable),
		.I2(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
		.O(SB_T0_WEST_SB_IN_B17_fan_in_O),
		.E1(SB_T4_SOUTH_SB_OUT_B17_enable_value_O),
		.I0(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out)
	);
	wire [1:0] SB_T0_WEST_SB_OUT_B17_FANOUT_I;
	assign SB_T0_WEST_SB_OUT_B17_FANOUT_I = {REG_T0_WEST_B17$SplitFifo_17_inst0_ready0[0], RMUX_T0_WEST_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T0_WEST_SB_OUT_B17_FANOUT(
		.O(SB_T0_WEST_SB_OUT_B17_FANOUT_O),
		.I(SB_T0_WEST_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T0_WEST_B17_out_sel)
	);
	SliceWrapper_31_0_1 SB_T0_WEST_SB_OUT_B17_enable_value(
		.I(config_reg_3_O),
		.O(SB_T0_WEST_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_31_1_4 SB_T0_WEST_SB_OUT_B17_sel_value(
		.I(config_reg_3_O),
		.O(SB_T0_WEST_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_31_4_5 SB_T1_EAST_SB_IN_B17_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_EAST_SB_IN_B17_enable_value_O)
	);
	FanoutHash_4F83851A40824F89 SB_T1_EAST_SB_IN_B17_fan_in(
		.E6(MEM_input_width_17_num_3_enable),
		.E3(MEM_input_width_17_num_0_enable),
		.I5(MEM_input_width_17_num_2_ready),
		.S6(MEM_input_width_17_num_3_out_sel),
		.E0(SB_T0_NORTH_SB_OUT_B17_enable_value_O),
		.S5(MEM_input_width_17_num_2_out_sel),
		.I6(MEM_input_width_17_num_3_ready),
		.S3(MEM_input_width_17_num_0_out_sel),
		.S4(MEM_input_width_17_num_1_out_sel),
		.I3(MEM_input_width_17_num_0_ready),
		.I4(MEM_input_width_17_num_1_ready),
		.S1(MUX_SB_T1_WEST_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel),
		.E2(SB_T2_SOUTH_SB_OUT_B17_enable_value_O),
		.E5(MEM_input_width_17_num_2_enable),
		.E4(MEM_input_width_17_num_1_enable),
		.I2(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
		.O(SB_T1_EAST_SB_IN_B17_fan_in_O),
		.E1(SB_T1_WEST_SB_OUT_B17_enable_value_O),
		.I0(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out)
	);
	wire [1:0] SB_T1_EAST_SB_OUT_B17_FANOUT_I;
	assign SB_T1_EAST_SB_OUT_B17_FANOUT_I = {REG_T1_EAST_B17$SplitFifo_17_inst0_ready0[0], RMUX_T1_EAST_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T1_EAST_SB_OUT_B17_FANOUT(
		.O(SB_T1_EAST_SB_OUT_B17_FANOUT_O),
		.I(SB_T1_EAST_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T1_EAST_B17_out_sel)
	);
	SliceWrapper_31_5_6 SB_T1_EAST_SB_OUT_B17_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_EAST_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_31_6_9 SB_T1_EAST_SB_OUT_B17_sel_value(
		.I(config_reg_3_O),
		.O(SB_T1_EAST_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_31_9_10 SB_T1_NORTH_SB_IN_B17_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_NORTH_SB_IN_B17_enable_value_O)
	);
	FanoutHash_4FADDC8F90390680 SB_T1_NORTH_SB_IN_B17_fan_in(
		.E6(MEM_input_width_17_num_3_enable),
		.E3(MEM_input_width_17_num_0_enable),
		.I5(MEM_input_width_17_num_2_ready),
		.S6(MEM_input_width_17_num_3_out_sel),
		.E0(SB_T2_EAST_SB_OUT_B17_enable_value_O),
		.S5(MEM_input_width_17_num_2_out_sel),
		.I6(MEM_input_width_17_num_3_ready),
		.S3(MEM_input_width_17_num_0_out_sel),
		.S4(MEM_input_width_17_num_1_out_sel),
		.I3(MEM_input_width_17_num_0_ready),
		.I4(MEM_input_width_17_num_1_ready),
		.S1(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T2_EAST_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T4_WEST_SB_OUT_B17_out_sel),
		.E2(SB_T4_WEST_SB_OUT_B17_enable_value_O),
		.E5(MEM_input_width_17_num_2_enable),
		.E4(MEM_input_width_17_num_1_enable),
		.I2(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
		.O(SB_T1_NORTH_SB_IN_B17_fan_in_O),
		.E1(SB_T1_SOUTH_SB_OUT_B17_enable_value_O),
		.I0(MUX_SB_T2_EAST_SB_OUT_B17_ready_out)
	);
	wire [1:0] SB_T1_NORTH_SB_OUT_B17_FANOUT_I;
	assign SB_T1_NORTH_SB_OUT_B17_FANOUT_I = {REG_T1_NORTH_B17$SplitFifo_17_inst0_ready0[0], RMUX_T1_NORTH_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T1_NORTH_SB_OUT_B17_FANOUT(
		.O(SB_T1_NORTH_SB_OUT_B17_FANOUT_O),
		.I(SB_T1_NORTH_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T1_NORTH_B17_out_sel)
	);
	SliceWrapper_31_10_11 SB_T1_NORTH_SB_OUT_B17_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_NORTH_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_31_11_14 SB_T1_NORTH_SB_OUT_B17_sel_value(
		.I(config_reg_3_O),
		.O(SB_T1_NORTH_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_31_14_15 SB_T1_SOUTH_SB_IN_B17_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_SOUTH_SB_IN_B17_enable_value_O)
	);
	FanoutHash_466EB88CFD0CAD7B SB_T1_SOUTH_SB_IN_B17_fan_in(
		.E6(MEM_input_width_17_num_3_enable),
		.E3(MEM_input_width_17_num_0_enable),
		.I5(MEM_input_width_17_num_2_ready),
		.S6(MEM_input_width_17_num_3_out_sel),
		.E0(SB_T2_EAST_SB_OUT_B17_enable_value_O),
		.S5(MEM_input_width_17_num_2_out_sel),
		.I6(MEM_input_width_17_num_3_ready),
		.S3(MEM_input_width_17_num_0_out_sel),
		.S4(MEM_input_width_17_num_1_out_sel),
		.I3(MEM_input_width_17_num_0_ready),
		.I4(MEM_input_width_17_num_1_ready),
		.S1(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T2_EAST_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T2_WEST_SB_OUT_B17_out_sel),
		.E2(SB_T2_WEST_SB_OUT_B17_enable_value_O),
		.E5(MEM_input_width_17_num_2_enable),
		.E4(MEM_input_width_17_num_1_enable),
		.I2(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out),
		.O(SB_T1_SOUTH_SB_IN_B17_fan_in_O),
		.E1(SB_T1_NORTH_SB_OUT_B17_enable_value_O),
		.I0(MUX_SB_T2_EAST_SB_OUT_B17_ready_out)
	);
	wire [1:0] SB_T1_SOUTH_SB_OUT_B17_FANOUT_I;
	assign SB_T1_SOUTH_SB_OUT_B17_FANOUT_I = {REG_T1_SOUTH_B17$SplitFifo_17_inst0_ready0[0], RMUX_T1_SOUTH_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T1_SOUTH_SB_OUT_B17_FANOUT(
		.O(SB_T1_SOUTH_SB_OUT_B17_FANOUT_O),
		.I(SB_T1_SOUTH_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T1_SOUTH_B17_out_sel)
	);
	SliceWrapper_31_15_16 SB_T1_SOUTH_SB_OUT_B17_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_SOUTH_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_31_16_19 SB_T1_SOUTH_SB_OUT_B17_sel_value(
		.I(config_reg_3_O),
		.O(SB_T1_SOUTH_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_31_19_20 SB_T1_WEST_SB_IN_B17_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_WEST_SB_IN_B17_enable_value_O)
	);
	FanoutHash_7ED1C80229B84786 SB_T1_WEST_SB_IN_B17_fan_in(
		.E6(MEM_input_width_17_num_3_enable),
		.E3(MEM_input_width_17_num_0_enable),
		.I5(MEM_input_width_17_num_2_ready),
		.S6(MEM_input_width_17_num_3_out_sel),
		.E0(SB_T4_NORTH_SB_OUT_B17_enable_value_O),
		.S5(MEM_input_width_17_num_2_out_sel),
		.I6(MEM_input_width_17_num_3_ready),
		.S3(MEM_input_width_17_num_0_out_sel),
		.S4(MEM_input_width_17_num_1_out_sel),
		.I3(MEM_input_width_17_num_0_ready),
		.I4(MEM_input_width_17_num_1_ready),
		.S1(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T1_EAST_SB_OUT_B17_out_sel),
		.E2(SB_T1_EAST_SB_OUT_B17_enable_value_O),
		.E5(MEM_input_width_17_num_2_enable),
		.E4(MEM_input_width_17_num_1_enable),
		.I2(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
		.O(SB_T1_WEST_SB_IN_B17_fan_in_O),
		.E1(SB_T0_SOUTH_SB_OUT_B17_enable_value_O),
		.I0(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out)
	);
	wire [1:0] SB_T1_WEST_SB_OUT_B17_FANOUT_I;
	assign SB_T1_WEST_SB_OUT_B17_FANOUT_I = {REG_T1_WEST_B17$SplitFifo_17_inst0_ready0[0], RMUX_T1_WEST_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T1_WEST_SB_OUT_B17_FANOUT(
		.O(SB_T1_WEST_SB_OUT_B17_FANOUT_O),
		.I(SB_T1_WEST_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T1_WEST_B17_out_sel)
	);
	SliceWrapper_31_20_21 SB_T1_WEST_SB_OUT_B17_enable_value(
		.I(config_reg_3_O),
		.O(SB_T1_WEST_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_31_21_24 SB_T1_WEST_SB_OUT_B17_sel_value(
		.I(config_reg_3_O),
		.O(SB_T1_WEST_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_31_24_25 SB_T2_EAST_SB_IN_B17_enable_value(
		.I(config_reg_3_O),
		.O(SB_T2_EAST_SB_IN_B17_enable_value_O)
	);
	FanoutHash_7F4660D1463D9234 SB_T2_EAST_SB_IN_B17_fan_in(
		.E6(MEM_input_width_17_num_3_enable),
		.E3(MEM_input_width_17_num_0_enable),
		.I5(MEM_input_width_17_num_2_ready),
		.S6(MEM_input_width_17_num_3_out_sel),
		.E0(SB_T1_NORTH_SB_OUT_B17_enable_value_O),
		.S5(MEM_input_width_17_num_2_out_sel),
		.I6(MEM_input_width_17_num_3_ready),
		.S3(MEM_input_width_17_num_0_out_sel),
		.S4(MEM_input_width_17_num_1_out_sel),
		.I3(MEM_input_width_17_num_0_ready),
		.I4(MEM_input_width_17_num_1_ready),
		.S1(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T2_WEST_SB_OUT_B17_out_sel),
		.E2(SB_T2_WEST_SB_OUT_B17_enable_value_O),
		.E5(MEM_input_width_17_num_2_enable),
		.E4(MEM_input_width_17_num_1_enable),
		.I2(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
		.O(SB_T2_EAST_SB_IN_B17_fan_in_O),
		.E1(SB_T1_SOUTH_SB_OUT_B17_enable_value_O),
		.I0(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out)
	);
	wire [1:0] SB_T2_EAST_SB_OUT_B17_FANOUT_I;
	assign SB_T2_EAST_SB_OUT_B17_FANOUT_I = {REG_T2_EAST_B17$SplitFifo_17_inst0_ready0[0], RMUX_T2_EAST_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T2_EAST_SB_OUT_B17_FANOUT(
		.O(SB_T2_EAST_SB_OUT_B17_FANOUT_O),
		.I(SB_T2_EAST_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T2_EAST_B17_out_sel)
	);
	SliceWrapper_31_25_26 SB_T2_EAST_SB_OUT_B17_enable_value(
		.I(config_reg_3_O),
		.O(SB_T2_EAST_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_31_26_29 SB_T2_EAST_SB_OUT_B17_sel_value(
		.I(config_reg_3_O),
		.O(SB_T2_EAST_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_31_29_30 SB_T2_NORTH_SB_IN_B17_enable_value(
		.I(config_reg_3_O),
		.O(SB_T2_NORTH_SB_IN_B17_enable_value_O)
	);
	FanoutHash_3B67229CB02928BA SB_T2_NORTH_SB_IN_B17_fan_in(
		.E6(MEM_input_width_17_num_3_enable),
		.E3(MEM_input_width_17_num_0_enable),
		.I5(MEM_input_width_17_num_2_ready),
		.S6(MEM_input_width_17_num_3_out_sel),
		.E0(SB_T3_EAST_SB_OUT_B17_enable_value_O),
		.S5(MEM_input_width_17_num_2_out_sel),
		.I6(MEM_input_width_17_num_3_ready),
		.S3(MEM_input_width_17_num_0_out_sel),
		.S4(MEM_input_width_17_num_1_out_sel),
		.I3(MEM_input_width_17_num_0_ready),
		.I4(MEM_input_width_17_num_1_ready),
		.S1(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T3_EAST_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T3_WEST_SB_OUT_B17_out_sel),
		.E2(SB_T3_WEST_SB_OUT_B17_enable_value_O),
		.E5(MEM_input_width_17_num_2_enable),
		.E4(MEM_input_width_17_num_1_enable),
		.I2(MUX_SB_T3_WEST_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
		.O(SB_T2_NORTH_SB_IN_B17_fan_in_O),
		.E1(SB_T2_SOUTH_SB_OUT_B17_enable_value_O),
		.I0(MUX_SB_T3_EAST_SB_OUT_B17_ready_out)
	);
	wire [1:0] SB_T2_NORTH_SB_OUT_B17_FANOUT_I;
	assign SB_T2_NORTH_SB_OUT_B17_FANOUT_I = {REG_T2_NORTH_B17$SplitFifo_17_inst0_ready0[0], RMUX_T2_NORTH_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T2_NORTH_SB_OUT_B17_FANOUT(
		.O(SB_T2_NORTH_SB_OUT_B17_FANOUT_O),
		.I(SB_T2_NORTH_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T2_NORTH_B17_out_sel)
	);
	SliceWrapper_31_30_31 SB_T2_NORTH_SB_OUT_B17_enable_value(
		.I(config_reg_3_O),
		.O(SB_T2_NORTH_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_30_0_3 SB_T2_NORTH_SB_OUT_B17_sel_value(
		.I(config_reg_4_O),
		.O(SB_T2_NORTH_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_30_3_4 SB_T2_SOUTH_SB_IN_B17_enable_value(
		.I(config_reg_4_O),
		.O(SB_T2_SOUTH_SB_IN_B17_enable_value_O)
	);
	FanoutHash_28125A548B305607 SB_T2_SOUTH_SB_IN_B17_fan_in(
		.E6(MEM_input_width_17_num_3_enable),
		.E3(MEM_input_width_17_num_0_enable),
		.I5(MEM_input_width_17_num_2_ready),
		.S6(MEM_input_width_17_num_3_out_sel),
		.E0(SB_T1_EAST_SB_OUT_B17_enable_value_O),
		.S5(MEM_input_width_17_num_2_out_sel),
		.I6(MEM_input_width_17_num_3_ready),
		.S3(MEM_input_width_17_num_0_out_sel),
		.S4(MEM_input_width_17_num_1_out_sel),
		.I3(MEM_input_width_17_num_0_ready),
		.I4(MEM_input_width_17_num_1_ready),
		.S1(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T1_EAST_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T3_WEST_SB_OUT_B17_out_sel),
		.E2(SB_T3_WEST_SB_OUT_B17_enable_value_O),
		.E5(MEM_input_width_17_num_2_enable),
		.E4(MEM_input_width_17_num_1_enable),
		.I2(MUX_SB_T3_WEST_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
		.O(SB_T2_SOUTH_SB_IN_B17_fan_in_O),
		.E1(SB_T2_NORTH_SB_OUT_B17_enable_value_O),
		.I0(MUX_SB_T1_EAST_SB_OUT_B17_ready_out)
	);
	wire [1:0] SB_T2_SOUTH_SB_OUT_B17_FANOUT_I;
	assign SB_T2_SOUTH_SB_OUT_B17_FANOUT_I = {REG_T2_SOUTH_B17$SplitFifo_17_inst0_ready0[0], RMUX_T2_SOUTH_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T2_SOUTH_SB_OUT_B17_FANOUT(
		.O(SB_T2_SOUTH_SB_OUT_B17_FANOUT_O),
		.I(SB_T2_SOUTH_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T2_SOUTH_B17_out_sel)
	);
	SliceWrapper_30_4_5 SB_T2_SOUTH_SB_OUT_B17_enable_value(
		.I(config_reg_4_O),
		.O(SB_T2_SOUTH_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_30_5_8 SB_T2_SOUTH_SB_OUT_B17_sel_value(
		.I(config_reg_4_O),
		.O(SB_T2_SOUTH_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_30_8_9 SB_T2_WEST_SB_IN_B17_enable_value(
		.I(config_reg_4_O),
		.O(SB_T2_WEST_SB_IN_B17_enable_value_O)
	);
	FanoutHash_752C11B748DD905C SB_T2_WEST_SB_IN_B17_fan_in(
		.E6(MEM_input_width_17_num_3_enable),
		.E3(MEM_input_width_17_num_0_enable),
		.I5(MEM_input_width_17_num_2_ready),
		.S6(MEM_input_width_17_num_3_out_sel),
		.E0(SB_T3_NORTH_SB_OUT_B17_enable_value_O),
		.S5(MEM_input_width_17_num_2_out_sel),
		.I6(MEM_input_width_17_num_3_ready),
		.S3(MEM_input_width_17_num_0_out_sel),
		.S4(MEM_input_width_17_num_1_out_sel),
		.I3(MEM_input_width_17_num_0_ready),
		.I4(MEM_input_width_17_num_1_ready),
		.S1(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T2_EAST_SB_OUT_B17_out_sel),
		.E2(SB_T2_EAST_SB_OUT_B17_enable_value_O),
		.E5(MEM_input_width_17_num_2_enable),
		.E4(MEM_input_width_17_num_1_enable),
		.I2(MUX_SB_T2_EAST_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
		.O(SB_T2_WEST_SB_IN_B17_fan_in_O),
		.E1(SB_T1_SOUTH_SB_OUT_B17_enable_value_O),
		.I0(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out)
	);
	wire [1:0] SB_T2_WEST_SB_OUT_B17_FANOUT_I;
	assign SB_T2_WEST_SB_OUT_B17_FANOUT_I = {REG_T2_WEST_B17$SplitFifo_17_inst0_ready0[0], RMUX_T2_WEST_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T2_WEST_SB_OUT_B17_FANOUT(
		.O(SB_T2_WEST_SB_OUT_B17_FANOUT_O),
		.I(SB_T2_WEST_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T2_WEST_B17_out_sel)
	);
	SliceWrapper_30_9_10 SB_T2_WEST_SB_OUT_B17_enable_value(
		.I(config_reg_4_O),
		.O(SB_T2_WEST_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_30_10_13 SB_T2_WEST_SB_OUT_B17_sel_value(
		.I(config_reg_4_O),
		.O(SB_T2_WEST_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_30_13_14 SB_T3_EAST_SB_IN_B17_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_EAST_SB_IN_B17_enable_value_O)
	);
	FanoutHash_43D5C80ABD816837 SB_T3_EAST_SB_IN_B17_fan_in(
		.E6(MEM_input_width_17_num_3_enable),
		.E3(MEM_input_width_17_num_0_enable),
		.I5(MEM_input_width_17_num_2_ready),
		.S6(MEM_input_width_17_num_3_out_sel),
		.E0(SB_T0_SOUTH_SB_OUT_B17_enable_value_O),
		.S5(MEM_input_width_17_num_2_out_sel),
		.I6(MEM_input_width_17_num_3_ready),
		.S3(MEM_input_width_17_num_0_out_sel),
		.S4(MEM_input_width_17_num_1_out_sel),
		.I3(MEM_input_width_17_num_0_ready),
		.I4(MEM_input_width_17_num_1_ready),
		.S1(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T3_WEST_SB_OUT_B17_out_sel),
		.E2(SB_T3_WEST_SB_OUT_B17_enable_value_O),
		.E5(MEM_input_width_17_num_2_enable),
		.E4(MEM_input_width_17_num_1_enable),
		.I2(MUX_SB_T3_WEST_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
		.O(SB_T3_EAST_SB_IN_B17_fan_in_O),
		.E1(SB_T2_NORTH_SB_OUT_B17_enable_value_O),
		.I0(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out)
	);
	wire [1:0] SB_T3_EAST_SB_OUT_B17_FANOUT_I;
	assign SB_T3_EAST_SB_OUT_B17_FANOUT_I = {REG_T3_EAST_B17$SplitFifo_17_inst0_ready0[0], RMUX_T3_EAST_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T3_EAST_SB_OUT_B17_FANOUT(
		.O(SB_T3_EAST_SB_OUT_B17_FANOUT_O),
		.I(SB_T3_EAST_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T3_EAST_B17_out_sel)
	);
	SliceWrapper_30_14_15 SB_T3_EAST_SB_OUT_B17_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_EAST_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_30_15_18 SB_T3_EAST_SB_OUT_B17_sel_value(
		.I(config_reg_4_O),
		.O(SB_T3_EAST_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_30_18_19 SB_T3_NORTH_SB_IN_B17_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_NORTH_SB_IN_B17_enable_value_O)
	);
	FanoutHash_69376833A2418E2 SB_T3_NORTH_SB_IN_B17_fan_in(
		.E6(MEM_input_width_17_num_3_enable),
		.E3(MEM_input_width_17_num_0_enable),
		.I5(MEM_input_width_17_num_2_ready),
		.S6(MEM_input_width_17_num_3_out_sel),
		.E0(SB_T2_WEST_SB_OUT_B17_enable_value_O),
		.S5(MEM_input_width_17_num_2_out_sel),
		.I6(MEM_input_width_17_num_3_ready),
		.S3(MEM_input_width_17_num_0_out_sel),
		.S4(MEM_input_width_17_num_1_out_sel),
		.I3(MEM_input_width_17_num_0_ready),
		.I4(MEM_input_width_17_num_1_ready),
		.S1(MUX_SB_T4_EAST_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T2_WEST_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel),
		.E2(SB_T3_SOUTH_SB_OUT_B17_enable_value_O),
		.E5(MEM_input_width_17_num_2_enable),
		.E4(MEM_input_width_17_num_1_enable),
		.I2(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T4_EAST_SB_OUT_B17_ready_out),
		.O(SB_T3_NORTH_SB_IN_B17_fan_in_O),
		.E1(SB_T4_EAST_SB_OUT_B17_enable_value_O),
		.I0(MUX_SB_T2_WEST_SB_OUT_B17_ready_out)
	);
	wire [1:0] SB_T3_NORTH_SB_OUT_B17_FANOUT_I;
	assign SB_T3_NORTH_SB_OUT_B17_FANOUT_I = {REG_T3_NORTH_B17$SplitFifo_17_inst0_ready0[0], RMUX_T3_NORTH_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T3_NORTH_SB_OUT_B17_FANOUT(
		.O(SB_T3_NORTH_SB_OUT_B17_FANOUT_O),
		.I(SB_T3_NORTH_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T3_NORTH_B17_out_sel)
	);
	SliceWrapper_30_19_20 SB_T3_NORTH_SB_OUT_B17_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_NORTH_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_30_20_23 SB_T3_NORTH_SB_OUT_B17_sel_value(
		.I(config_reg_4_O),
		.O(SB_T3_NORTH_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_30_23_24 SB_T3_SOUTH_SB_IN_B17_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_SOUTH_SB_IN_B17_enable_value_O)
	);
	FanoutHash_66A75CC8494A4D6B SB_T3_SOUTH_SB_IN_B17_fan_in(
		.E6(MEM_input_width_17_num_3_enable),
		.E3(MEM_input_width_17_num_0_enable),
		.I5(MEM_input_width_17_num_2_ready),
		.S6(MEM_input_width_17_num_3_out_sel),
		.E0(SB_T0_EAST_SB_OUT_B17_enable_value_O),
		.S5(MEM_input_width_17_num_2_out_sel),
		.I6(MEM_input_width_17_num_3_ready),
		.S3(MEM_input_width_17_num_0_out_sel),
		.S4(MEM_input_width_17_num_1_out_sel),
		.I3(MEM_input_width_17_num_0_ready),
		.I4(MEM_input_width_17_num_1_ready),
		.S1(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T0_EAST_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T4_WEST_SB_OUT_B17_out_sel),
		.E2(SB_T4_WEST_SB_OUT_B17_enable_value_O),
		.E5(MEM_input_width_17_num_2_enable),
		.E4(MEM_input_width_17_num_1_enable),
		.I2(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out),
		.O(SB_T3_SOUTH_SB_IN_B17_fan_in_O),
		.E1(SB_T3_NORTH_SB_OUT_B17_enable_value_O),
		.I0(MUX_SB_T0_EAST_SB_OUT_B17_ready_out)
	);
	wire [1:0] SB_T3_SOUTH_SB_OUT_B17_FANOUT_I;
	assign SB_T3_SOUTH_SB_OUT_B17_FANOUT_I = {REG_T3_SOUTH_B17$SplitFifo_17_inst0_ready0[0], RMUX_T3_SOUTH_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T3_SOUTH_SB_OUT_B17_FANOUT(
		.O(SB_T3_SOUTH_SB_OUT_B17_FANOUT_O),
		.I(SB_T3_SOUTH_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T3_SOUTH_B17_out_sel)
	);
	SliceWrapper_30_24_25 SB_T3_SOUTH_SB_OUT_B17_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_SOUTH_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_30_25_28 SB_T3_SOUTH_SB_OUT_B17_sel_value(
		.I(config_reg_4_O),
		.O(SB_T3_SOUTH_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_30_28_29 SB_T3_WEST_SB_IN_B17_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_WEST_SB_IN_B17_enable_value_O)
	);
	FanoutHash_31AE65CCDD94603 SB_T3_WEST_SB_IN_B17_fan_in(
		.E6(MEM_input_width_17_num_3_enable),
		.E3(MEM_input_width_17_num_0_enable),
		.I5(MEM_input_width_17_num_2_ready),
		.S6(MEM_input_width_17_num_3_out_sel),
		.E0(SB_T2_NORTH_SB_OUT_B17_enable_value_O),
		.S5(MEM_input_width_17_num_2_out_sel),
		.I6(MEM_input_width_17_num_3_ready),
		.S3(MEM_input_width_17_num_0_out_sel),
		.S4(MEM_input_width_17_num_1_out_sel),
		.I3(MEM_input_width_17_num_0_ready),
		.I4(MEM_input_width_17_num_1_ready),
		.S1(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T3_EAST_SB_OUT_B17_out_sel),
		.E2(SB_T3_EAST_SB_OUT_B17_enable_value_O),
		.E5(MEM_input_width_17_num_2_enable),
		.E4(MEM_input_width_17_num_1_enable),
		.I2(MUX_SB_T3_EAST_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
		.O(SB_T3_WEST_SB_IN_B17_fan_in_O),
		.E1(SB_T2_SOUTH_SB_OUT_B17_enable_value_O),
		.I0(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out)
	);
	wire [1:0] SB_T3_WEST_SB_OUT_B17_FANOUT_I;
	assign SB_T3_WEST_SB_OUT_B17_FANOUT_I = {REG_T3_WEST_B17$SplitFifo_17_inst0_ready0[0], RMUX_T3_WEST_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T3_WEST_SB_OUT_B17_FANOUT(
		.O(SB_T3_WEST_SB_OUT_B17_FANOUT_O),
		.I(SB_T3_WEST_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T3_WEST_B17_out_sel)
	);
	SliceWrapper_30_29_30 SB_T3_WEST_SB_OUT_B17_enable_value(
		.I(config_reg_4_O),
		.O(SB_T3_WEST_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_23_0_3 SB_T3_WEST_SB_OUT_B17_sel_value(
		.I(config_reg_5_O),
		.O(SB_T3_WEST_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_23_3_4 SB_T4_EAST_SB_IN_B17_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_EAST_SB_IN_B17_enable_value_O)
	);
	FanoutHash_5D7AEC1255CDC1CC SB_T4_EAST_SB_IN_B17_fan_in(
		.E6(MEM_input_width_17_num_3_enable),
		.E3(MEM_input_width_17_num_0_enable),
		.I5(MEM_input_width_17_num_2_ready),
		.S6(MEM_input_width_17_num_3_out_sel),
		.E0(SB_T3_NORTH_SB_OUT_B17_enable_value_O),
		.S5(MEM_input_width_17_num_2_out_sel),
		.I6(MEM_input_width_17_num_3_ready),
		.S3(MEM_input_width_17_num_0_out_sel),
		.S4(MEM_input_width_17_num_1_out_sel),
		.I3(MEM_input_width_17_num_0_ready),
		.I4(MEM_input_width_17_num_1_ready),
		.S1(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T4_WEST_SB_OUT_B17_out_sel),
		.E2(SB_T4_WEST_SB_OUT_B17_enable_value_O),
		.E5(MEM_input_width_17_num_2_enable),
		.E4(MEM_input_width_17_num_1_enable),
		.I2(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
		.O(SB_T4_EAST_SB_IN_B17_fan_in_O),
		.E1(SB_T4_SOUTH_SB_OUT_B17_enable_value_O),
		.I0(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out)
	);
	wire [1:0] SB_T4_EAST_SB_OUT_B17_FANOUT_I;
	assign SB_T4_EAST_SB_OUT_B17_FANOUT_I = {REG_T4_EAST_B17$SplitFifo_17_inst0_ready0[0], RMUX_T4_EAST_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T4_EAST_SB_OUT_B17_FANOUT(
		.O(SB_T4_EAST_SB_OUT_B17_FANOUT_O),
		.I(SB_T4_EAST_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T4_EAST_B17_out_sel)
	);
	SliceWrapper_23_4_5 SB_T4_EAST_SB_OUT_B17_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_EAST_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_23_5_8 SB_T4_EAST_SB_OUT_B17_sel_value(
		.I(config_reg_5_O),
		.O(SB_T4_EAST_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_23_8_9 SB_T4_NORTH_SB_IN_B17_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_NORTH_SB_IN_B17_enable_value_O)
	);
	FanoutHash_184DFC10DAF19BE9 SB_T4_NORTH_SB_IN_B17_fan_in(
		.E6(MEM_input_width_17_num_3_enable),
		.E3(MEM_input_width_17_num_0_enable),
		.I5(MEM_input_width_17_num_2_ready),
		.S6(MEM_input_width_17_num_3_out_sel),
		.E0(SB_T1_WEST_SB_OUT_B17_enable_value_O),
		.S5(MEM_input_width_17_num_2_out_sel),
		.I6(MEM_input_width_17_num_3_ready),
		.S3(MEM_input_width_17_num_0_out_sel),
		.S4(MEM_input_width_17_num_1_out_sel),
		.I3(MEM_input_width_17_num_0_ready),
		.I4(MEM_input_width_17_num_1_ready),
		.S1(MUX_SB_T0_EAST_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T1_WEST_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel),
		.E2(SB_T4_SOUTH_SB_OUT_B17_enable_value_O),
		.E5(MEM_input_width_17_num_2_enable),
		.E4(MEM_input_width_17_num_1_enable),
		.I2(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
		.O(SB_T4_NORTH_SB_IN_B17_fan_in_O),
		.E1(SB_T0_EAST_SB_OUT_B17_enable_value_O),
		.I0(MUX_SB_T1_WEST_SB_OUT_B17_ready_out)
	);
	wire [1:0] SB_T4_NORTH_SB_OUT_B17_FANOUT_I;
	assign SB_T4_NORTH_SB_OUT_B17_FANOUT_I = {REG_T4_NORTH_B17$SplitFifo_17_inst0_ready0[0], RMUX_T4_NORTH_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T4_NORTH_SB_OUT_B17_FANOUT(
		.O(SB_T4_NORTH_SB_OUT_B17_FANOUT_O),
		.I(SB_T4_NORTH_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T4_NORTH_B17_out_sel)
	);
	SliceWrapper_23_9_10 SB_T4_NORTH_SB_OUT_B17_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_NORTH_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_23_10_13 SB_T4_NORTH_SB_OUT_B17_sel_value(
		.I(config_reg_5_O),
		.O(SB_T4_NORTH_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_23_13_14 SB_T4_SOUTH_SB_IN_B17_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_SOUTH_SB_IN_B17_enable_value_O)
	);
	FanoutHash_26B6474864379B6A SB_T4_SOUTH_SB_IN_B17_fan_in(
		.E6(MEM_input_width_17_num_3_enable),
		.E3(MEM_input_width_17_num_0_enable),
		.I5(MEM_input_width_17_num_2_ready),
		.S6(MEM_input_width_17_num_3_out_sel),
		.E0(SB_T0_WEST_SB_OUT_B17_enable_value_O),
		.S5(MEM_input_width_17_num_2_out_sel),
		.I6(MEM_input_width_17_num_3_ready),
		.S3(MEM_input_width_17_num_0_out_sel),
		.S4(MEM_input_width_17_num_1_out_sel),
		.I3(MEM_input_width_17_num_0_ready),
		.I4(MEM_input_width_17_num_1_ready),
		.S1(MUX_SB_T4_EAST_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T0_WEST_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel),
		.E2(SB_T4_NORTH_SB_OUT_B17_enable_value_O),
		.E5(MEM_input_width_17_num_2_enable),
		.E4(MEM_input_width_17_num_1_enable),
		.I2(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T4_EAST_SB_OUT_B17_ready_out),
		.O(SB_T4_SOUTH_SB_IN_B17_fan_in_O),
		.E1(SB_T4_EAST_SB_OUT_B17_enable_value_O),
		.I0(MUX_SB_T0_WEST_SB_OUT_B17_ready_out)
	);
	wire [1:0] SB_T4_SOUTH_SB_OUT_B17_FANOUT_I;
	assign SB_T4_SOUTH_SB_OUT_B17_FANOUT_I = {REG_T4_SOUTH_B17$SplitFifo_17_inst0_ready0[0], RMUX_T4_SOUTH_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T4_SOUTH_SB_OUT_B17_FANOUT(
		.O(SB_T4_SOUTH_SB_OUT_B17_FANOUT_O),
		.I(SB_T4_SOUTH_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T4_SOUTH_B17_out_sel)
	);
	SliceWrapper_23_14_15 SB_T4_SOUTH_SB_OUT_B17_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_SOUTH_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_23_15_18 SB_T4_SOUTH_SB_OUT_B17_sel_value(
		.I(config_reg_5_O),
		.O(SB_T4_SOUTH_SB_OUT_B17_sel_value_O)
	);
	SliceWrapper_23_18_19 SB_T4_WEST_SB_IN_B17_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_WEST_SB_IN_B17_enable_value_O)
	);
	FanoutHash_1816466D6957000 SB_T4_WEST_SB_IN_B17_fan_in(
		.E6(MEM_input_width_17_num_3_enable),
		.E3(MEM_input_width_17_num_0_enable),
		.I5(MEM_input_width_17_num_2_ready),
		.S6(MEM_input_width_17_num_3_out_sel),
		.E0(SB_T1_NORTH_SB_OUT_B17_enable_value_O),
		.S5(MEM_input_width_17_num_2_out_sel),
		.I6(MEM_input_width_17_num_3_ready),
		.S3(MEM_input_width_17_num_0_out_sel),
		.S4(MEM_input_width_17_num_1_out_sel),
		.I3(MEM_input_width_17_num_0_ready),
		.I4(MEM_input_width_17_num_1_ready),
		.S1(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel),
		.S0(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel),
		.S2(MUX_SB_T4_EAST_SB_OUT_B17_out_sel),
		.E2(SB_T4_EAST_SB_OUT_B17_enable_value_O),
		.E5(MEM_input_width_17_num_2_enable),
		.E4(MEM_input_width_17_num_1_enable),
		.I2(MUX_SB_T4_EAST_SB_OUT_B17_ready_out),
		.I1(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
		.O(SB_T4_WEST_SB_IN_B17_fan_in_O),
		.E1(SB_T3_SOUTH_SB_OUT_B17_enable_value_O),
		.I0(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out)
	);
	wire [1:0] SB_T4_WEST_SB_OUT_B17_FANOUT_I;
	assign SB_T4_WEST_SB_OUT_B17_FANOUT_I = {REG_T4_WEST_B17$SplitFifo_17_inst0_ready0[0], RMUX_T4_WEST_B17_ready_out};
	ExclusiveNodeFanout_H2 SB_T4_WEST_SB_OUT_B17_FANOUT(
		.O(SB_T4_WEST_SB_OUT_B17_FANOUT_O),
		.I(SB_T4_WEST_SB_OUT_B17_FANOUT_I),
		.S(RMUX_T4_WEST_B17_out_sel)
	);
	SliceWrapper_23_19_20 SB_T4_WEST_SB_OUT_B17_enable_value(
		.I(config_reg_5_O),
		.O(SB_T4_WEST_SB_OUT_B17_enable_value_O)
	);
	SliceWrapper_23_20_23 SB_T4_WEST_SB_OUT_B17_sel_value(
		.I(config_reg_5_O),
		.O(SB_T4_WEST_SB_OUT_B17_sel_value_O)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T0_EAST_SB_IN_B17(
		.I(SB_T0_EAST_SB_IN_B17),
		.O(WIRE_SB_T0_EAST_SB_IN_B17_O),
		.ready_in(SB_T0_EAST_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T0_EAST_SB_IN_B17_ready_out),
		.valid_in(SB_T0_EAST_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T0_EAST_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T0_NORTH_SB_IN_B17(
		.I(SB_T0_NORTH_SB_IN_B17),
		.O(WIRE_SB_T0_NORTH_SB_IN_B17_O),
		.ready_in(SB_T0_NORTH_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T0_NORTH_SB_IN_B17_ready_out),
		.valid_in(SB_T0_NORTH_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T0_NORTH_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T0_SOUTH_SB_IN_B17(
		.I(SB_T0_SOUTH_SB_IN_B17),
		.O(WIRE_SB_T0_SOUTH_SB_IN_B17_O),
		.ready_in(SB_T0_SOUTH_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T0_SOUTH_SB_IN_B17_ready_out),
		.valid_in(SB_T0_SOUTH_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T0_SOUTH_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T0_WEST_SB_IN_B17(
		.I(SB_T0_WEST_SB_IN_B17),
		.O(WIRE_SB_T0_WEST_SB_IN_B17_O),
		.ready_in(SB_T0_WEST_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T0_WEST_SB_IN_B17_ready_out),
		.valid_in(SB_T0_WEST_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T0_WEST_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T1_EAST_SB_IN_B17(
		.I(SB_T1_EAST_SB_IN_B17),
		.O(WIRE_SB_T1_EAST_SB_IN_B17_O),
		.ready_in(SB_T1_EAST_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T1_EAST_SB_IN_B17_ready_out),
		.valid_in(SB_T1_EAST_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T1_EAST_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T1_NORTH_SB_IN_B17(
		.I(SB_T1_NORTH_SB_IN_B17),
		.O(WIRE_SB_T1_NORTH_SB_IN_B17_O),
		.ready_in(SB_T1_NORTH_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T1_NORTH_SB_IN_B17_ready_out),
		.valid_in(SB_T1_NORTH_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T1_NORTH_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T1_SOUTH_SB_IN_B17(
		.I(SB_T1_SOUTH_SB_IN_B17),
		.O(WIRE_SB_T1_SOUTH_SB_IN_B17_O),
		.ready_in(SB_T1_SOUTH_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T1_SOUTH_SB_IN_B17_ready_out),
		.valid_in(SB_T1_SOUTH_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T1_SOUTH_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T1_WEST_SB_IN_B17(
		.I(SB_T1_WEST_SB_IN_B17),
		.O(WIRE_SB_T1_WEST_SB_IN_B17_O),
		.ready_in(SB_T1_WEST_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T1_WEST_SB_IN_B17_ready_out),
		.valid_in(SB_T1_WEST_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T1_WEST_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T2_EAST_SB_IN_B17(
		.I(SB_T2_EAST_SB_IN_B17),
		.O(WIRE_SB_T2_EAST_SB_IN_B17_O),
		.ready_in(SB_T2_EAST_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T2_EAST_SB_IN_B17_ready_out),
		.valid_in(SB_T2_EAST_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T2_EAST_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T2_NORTH_SB_IN_B17(
		.I(SB_T2_NORTH_SB_IN_B17),
		.O(WIRE_SB_T2_NORTH_SB_IN_B17_O),
		.ready_in(SB_T2_NORTH_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T2_NORTH_SB_IN_B17_ready_out),
		.valid_in(SB_T2_NORTH_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T2_NORTH_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T2_SOUTH_SB_IN_B17(
		.I(SB_T2_SOUTH_SB_IN_B17),
		.O(WIRE_SB_T2_SOUTH_SB_IN_B17_O),
		.ready_in(SB_T2_SOUTH_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T2_SOUTH_SB_IN_B17_ready_out),
		.valid_in(SB_T2_SOUTH_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T2_SOUTH_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T2_WEST_SB_IN_B17(
		.I(SB_T2_WEST_SB_IN_B17),
		.O(WIRE_SB_T2_WEST_SB_IN_B17_O),
		.ready_in(SB_T2_WEST_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T2_WEST_SB_IN_B17_ready_out),
		.valid_in(SB_T2_WEST_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T2_WEST_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T3_EAST_SB_IN_B17(
		.I(SB_T3_EAST_SB_IN_B17),
		.O(WIRE_SB_T3_EAST_SB_IN_B17_O),
		.ready_in(SB_T3_EAST_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T3_EAST_SB_IN_B17_ready_out),
		.valid_in(SB_T3_EAST_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T3_EAST_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T3_NORTH_SB_IN_B17(
		.I(SB_T3_NORTH_SB_IN_B17),
		.O(WIRE_SB_T3_NORTH_SB_IN_B17_O),
		.ready_in(SB_T3_NORTH_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T3_NORTH_SB_IN_B17_ready_out),
		.valid_in(SB_T3_NORTH_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T3_NORTH_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T3_SOUTH_SB_IN_B17(
		.I(SB_T3_SOUTH_SB_IN_B17),
		.O(WIRE_SB_T3_SOUTH_SB_IN_B17_O),
		.ready_in(SB_T3_SOUTH_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T3_SOUTH_SB_IN_B17_ready_out),
		.valid_in(SB_T3_SOUTH_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T3_SOUTH_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T3_WEST_SB_IN_B17(
		.I(SB_T3_WEST_SB_IN_B17),
		.O(WIRE_SB_T3_WEST_SB_IN_B17_O),
		.ready_in(SB_T3_WEST_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T3_WEST_SB_IN_B17_ready_out),
		.valid_in(SB_T3_WEST_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T3_WEST_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T4_EAST_SB_IN_B17(
		.I(SB_T4_EAST_SB_IN_B17),
		.O(WIRE_SB_T4_EAST_SB_IN_B17_O),
		.ready_in(SB_T4_EAST_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T4_EAST_SB_IN_B17_ready_out),
		.valid_in(SB_T4_EAST_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T4_EAST_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T4_NORTH_SB_IN_B17(
		.I(SB_T4_NORTH_SB_IN_B17),
		.O(WIRE_SB_T4_NORTH_SB_IN_B17_O),
		.ready_in(SB_T4_NORTH_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T4_NORTH_SB_IN_B17_ready_out),
		.valid_in(SB_T4_NORTH_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T4_NORTH_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T4_SOUTH_SB_IN_B17(
		.I(SB_T4_SOUTH_SB_IN_B17),
		.O(WIRE_SB_T4_SOUTH_SB_IN_B17_O),
		.ready_in(SB_T4_SOUTH_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T4_SOUTH_SB_IN_B17_ready_out),
		.valid_in(SB_T4_SOUTH_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T4_SOUTH_SB_IN_B17_valid_out)
	);
	MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T4_WEST_SB_IN_B17(
		.I(SB_T4_WEST_SB_IN_B17),
		.O(WIRE_SB_T4_WEST_SB_IN_B17_O),
		.ready_in(SB_T4_WEST_SB_IN_B17_fan_in_O[0]),
		.ready_out(WIRE_SB_T4_WEST_SB_IN_B17_ready_out),
		.valid_in(SB_T4_WEST_SB_IN_B17_valid_in),
		.valid_out(WIRE_SB_T4_WEST_SB_IN_B17_valid_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_23_32_inst0$bit_const_0_None(.out(ZextWrapper_23_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_23_32_inst0$self_O_out;
	assign ZextWrapper_23_32_inst0$self_O_out = {ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, ZextWrapper_23_32_inst0$bit_const_0_None_out, config_reg_5_O};
	mantle_wire__typeBitIn32 ZextWrapper_23_32_inst0$self_O(
		.in(ZextWrapper_23_32_inst0$self_O_in),
		.out(ZextWrapper_23_32_inst0$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_30_32_inst0$bit_const_0_None(.out(ZextWrapper_30_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_30_32_inst0$self_O_out;
	assign ZextWrapper_30_32_inst0$self_O_out = {ZextWrapper_30_32_inst0$bit_const_0_None_out, ZextWrapper_30_32_inst0$bit_const_0_None_out, config_reg_4_O};
	mantle_wire__typeBitIn32 ZextWrapper_30_32_inst0$self_O(
		.in(ZextWrapper_30_32_inst0$self_O_in),
		.out(ZextWrapper_30_32_inst0$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_31_32_inst0$bit_const_0_None(.out(ZextWrapper_31_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_31_32_inst0$self_O_out;
	assign ZextWrapper_31_32_inst0$self_O_out = {ZextWrapper_31_32_inst0$bit_const_0_None_out, config_reg_3_O};
	mantle_wire__typeBitIn32 ZextWrapper_31_32_inst0$self_O(
		.in(ZextWrapper_31_32_inst0$self_O_in),
		.out(ZextWrapper_31_32_inst0$self_O_out)
	);
	coreir_and #(.width(1)) and1_inst0(
		.in0(coreir_eq_1_inst0_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst0_out)
	);
	coreir_and #(.width(1)) and1_inst1(
		.in0(coreir_eq_1_inst1_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst1_out)
	);
	coreir_and #(.width(1)) and1_inst10(
		.in0(coreir_eq_1_inst10_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst10_out)
	);
	coreir_and #(.width(1)) and1_inst11(
		.in0(coreir_eq_1_inst11_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst11_out)
	);
	coreir_and #(.width(1)) and1_inst12(
		.in0(coreir_eq_1_inst12_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst12_out)
	);
	coreir_and #(.width(1)) and1_inst13(
		.in0(coreir_eq_1_inst13_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst13_out)
	);
	coreir_and #(.width(1)) and1_inst14(
		.in0(coreir_eq_1_inst14_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst14_out)
	);
	coreir_and #(.width(1)) and1_inst15(
		.in0(coreir_eq_1_inst15_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst15_out)
	);
	coreir_and #(.width(1)) and1_inst16(
		.in0(coreir_eq_1_inst16_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst16_out)
	);
	coreir_and #(.width(1)) and1_inst17(
		.in0(coreir_eq_1_inst17_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst17_out)
	);
	coreir_and #(.width(1)) and1_inst18(
		.in0(coreir_eq_1_inst18_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst18_out)
	);
	coreir_and #(.width(1)) and1_inst19(
		.in0(coreir_eq_1_inst19_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst19_out)
	);
	coreir_and #(.width(1)) and1_inst2(
		.in0(coreir_eq_1_inst2_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst2_out)
	);
	coreir_and #(.width(1)) and1_inst3(
		.in0(coreir_eq_1_inst3_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst3_out)
	);
	coreir_and #(.width(1)) and1_inst4(
		.in0(coreir_eq_1_inst4_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst4_out)
	);
	coreir_and #(.width(1)) and1_inst5(
		.in0(coreir_eq_1_inst5_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst5_out)
	);
	coreir_and #(.width(1)) and1_inst6(
		.in0(coreir_eq_1_inst6_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst6_out)
	);
	coreir_and #(.width(1)) and1_inst7(
		.in0(coreir_eq_1_inst7_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst7_out)
	);
	coreir_and #(.width(1)) and1_inst8(
		.in0(coreir_eq_1_inst8_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst8_out)
	);
	coreir_and #(.width(1)) and1_inst9(
		.in0(coreir_eq_1_inst9_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst9_out)
	);
	wire [7:0] config_reg_0_config_addr;
	assign config_reg_0_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4], self_config_config_addr_out[3], self_config_config_addr_out[2:0]};
	ConfigRegister_32_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_reg_0_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_1_config_addr;
	assign config_reg_1_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4], self_config_config_addr_out[3], self_config_config_addr_out[2:0]};
	ConfigRegister_32_8_32_1 config_reg_1(
		.clk(clk),
		.reset(reset),
		.O(config_reg_1_O),
		.config_addr(config_reg_1_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_2_config_addr;
	assign config_reg_2_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4], self_config_config_addr_out[3], self_config_config_addr_out[2:0]};
	ConfigRegister_32_8_32_2 config_reg_2(
		.clk(clk),
		.reset(reset),
		.O(config_reg_2_O),
		.config_addr(config_reg_2_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_3_config_addr;
	assign config_reg_3_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4], self_config_config_addr_out[3], self_config_config_addr_out[2:0]};
	ConfigRegister_31_8_32_3 config_reg_3(
		.clk(clk),
		.reset(reset),
		.O(config_reg_3_O),
		.config_addr(config_reg_3_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_4_config_addr;
	assign config_reg_4_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4], self_config_config_addr_out[3], self_config_config_addr_out[2:0]};
	ConfigRegister_30_8_32_4 config_reg_4(
		.clk(clk),
		.reset(reset),
		.O(config_reg_4_O),
		.config_addr(config_reg_4_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_5_config_addr;
	assign config_reg_5_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4], self_config_config_addr_out[3], self_config_config_addr_out[2:0]};
	ConfigRegister_23_8_32_5 config_reg_5(
		.clk(clk),
		.reset(reset),
		.O(config_reg_5_O),
		.config_addr(config_reg_5_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	coreir_const #(
		.value(1'h1),
		.width(1)
	) const_1_1(.out(const_1_1_out));
	coreir_eq #(.width(1)) coreir_eq_1_inst0(
		.in0(const_1_1_out),
		.in1(RMUX_T0_NORTH_B17_sel_value_O),
		.out(coreir_eq_1_inst0_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst1(
		.in0(const_1_1_out),
		.in1(RMUX_T0_SOUTH_B17_sel_value_O),
		.out(coreir_eq_1_inst1_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst10(
		.in0(const_1_1_out),
		.in1(RMUX_T2_EAST_B17_sel_value_O),
		.out(coreir_eq_1_inst10_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst11(
		.in0(const_1_1_out),
		.in1(RMUX_T2_WEST_B17_sel_value_O),
		.out(coreir_eq_1_inst11_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst12(
		.in0(const_1_1_out),
		.in1(RMUX_T3_NORTH_B17_sel_value_O),
		.out(coreir_eq_1_inst12_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst13(
		.in0(const_1_1_out),
		.in1(RMUX_T3_SOUTH_B17_sel_value_O),
		.out(coreir_eq_1_inst13_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst14(
		.in0(const_1_1_out),
		.in1(RMUX_T3_EAST_B17_sel_value_O),
		.out(coreir_eq_1_inst14_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst15(
		.in0(const_1_1_out),
		.in1(RMUX_T3_WEST_B17_sel_value_O),
		.out(coreir_eq_1_inst15_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst16(
		.in0(const_1_1_out),
		.in1(RMUX_T4_NORTH_B17_sel_value_O),
		.out(coreir_eq_1_inst16_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst17(
		.in0(const_1_1_out),
		.in1(RMUX_T4_SOUTH_B17_sel_value_O),
		.out(coreir_eq_1_inst17_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst18(
		.in0(const_1_1_out),
		.in1(RMUX_T4_EAST_B17_sel_value_O),
		.out(coreir_eq_1_inst18_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst19(
		.in0(const_1_1_out),
		.in1(RMUX_T4_WEST_B17_sel_value_O),
		.out(coreir_eq_1_inst19_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst2(
		.in0(const_1_1_out),
		.in1(RMUX_T0_EAST_B17_sel_value_O),
		.out(coreir_eq_1_inst2_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst3(
		.in0(const_1_1_out),
		.in1(RMUX_T0_WEST_B17_sel_value_O),
		.out(coreir_eq_1_inst3_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst4(
		.in0(const_1_1_out),
		.in1(RMUX_T1_NORTH_B17_sel_value_O),
		.out(coreir_eq_1_inst4_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst5(
		.in0(const_1_1_out),
		.in1(RMUX_T1_SOUTH_B17_sel_value_O),
		.out(coreir_eq_1_inst5_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst6(
		.in0(const_1_1_out),
		.in1(RMUX_T1_EAST_B17_sel_value_O),
		.out(coreir_eq_1_inst6_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst7(
		.in0(const_1_1_out),
		.in1(RMUX_T1_WEST_B17_sel_value_O),
		.out(coreir_eq_1_inst7_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst8(
		.in0(const_1_1_out),
		.in1(RMUX_T2_NORTH_B17_sel_value_O),
		.out(coreir_eq_1_inst8_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst9(
		.in0(const_1_1_out),
		.in1(RMUX_T2_SOUTH_B17_sel_value_O),
		.out(coreir_eq_1_inst9_out)
	);
	wire [191:0] mux_aoi_6_32_inst0_I;
	assign mux_aoi_6_32_inst0_I[160+:32] = ZextWrapper_23_32_inst0$self_O_in;
	assign mux_aoi_6_32_inst0_I[128+:32] = ZextWrapper_30_32_inst0$self_O_in;
	assign mux_aoi_6_32_inst0_I[96+:32] = ZextWrapper_31_32_inst0$self_O_in;
	assign mux_aoi_6_32_inst0_I[64+:32] = config_reg_2_O;
	assign mux_aoi_6_32_inst0_I[32+:32] = config_reg_1_O;
	assign mux_aoi_6_32_inst0_I[0+:32] = config_reg_0_O;
	mux_aoi_6_32 mux_aoi_6_32_inst0(
		.I(mux_aoi_6_32_inst0_I),
		.O(mux_aoi_6_32_inst0_O),
		.S(self_config_config_addr_out[2:0]),
		.out_sel(mux_aoi_6_32_inst0_out_sel)
	);
	mantle_wire__typeBit8 self_config_config_addr(
		.in(config_config_addr),
		.out(self_config_config_addr_out)
	);
	assign MEM_output_width_17_num_0_ready_out = CB_MEM_output_width_17_num_0_fan_in_O[0];
	assign MEM_output_width_17_num_1_ready_out = CB_MEM_output_width_17_num_1_fan_in_O[0];
	assign MEM_output_width_17_num_2_ready_out = CB_MEM_output_width_17_num_2_fan_in_O[0];
	assign SB_T0_EAST_SB_IN_B17_enable = SB_T0_EAST_SB_IN_B17_enable_value_O[0];
	assign SB_T0_EAST_SB_IN_B17_ready_out = WIRE_SB_T0_EAST_SB_IN_B17_ready_out;
	assign SB_T0_EAST_SB_OUT_B17 = RMUX_T0_EAST_B17_O;
	assign SB_T0_EAST_SB_OUT_B17_enable = SB_T0_EAST_SB_OUT_B17_enable_value_O[0];
	assign SB_T0_EAST_SB_OUT_B17_valid_out = RMUX_T0_EAST_B17_valid_out;
	assign SB_T0_NORTH_SB_IN_B17_enable = SB_T0_NORTH_SB_IN_B17_enable_value_O[0];
	assign SB_T0_NORTH_SB_IN_B17_ready_out = WIRE_SB_T0_NORTH_SB_IN_B17_ready_out;
	assign SB_T0_NORTH_SB_OUT_B17 = RMUX_T0_NORTH_B17_O;
	assign SB_T0_NORTH_SB_OUT_B17_enable = SB_T0_NORTH_SB_OUT_B17_enable_value_O[0];
	assign SB_T0_NORTH_SB_OUT_B17_valid_out = RMUX_T0_NORTH_B17_valid_out;
	assign SB_T0_SOUTH_SB_IN_B17_enable = SB_T0_SOUTH_SB_IN_B17_enable_value_O[0];
	assign SB_T0_SOUTH_SB_IN_B17_ready_out = WIRE_SB_T0_SOUTH_SB_IN_B17_ready_out;
	assign SB_T0_SOUTH_SB_OUT_B17 = RMUX_T0_SOUTH_B17_O;
	assign SB_T0_SOUTH_SB_OUT_B17_enable = SB_T0_SOUTH_SB_OUT_B17_enable_value_O[0];
	assign SB_T0_SOUTH_SB_OUT_B17_valid_out = RMUX_T0_SOUTH_B17_valid_out;
	assign SB_T0_WEST_SB_IN_B17_enable = SB_T0_WEST_SB_IN_B17_enable_value_O[0];
	assign SB_T0_WEST_SB_IN_B17_ready_out = WIRE_SB_T0_WEST_SB_IN_B17_ready_out;
	assign SB_T0_WEST_SB_OUT_B17 = RMUX_T0_WEST_B17_O;
	assign SB_T0_WEST_SB_OUT_B17_enable = SB_T0_WEST_SB_OUT_B17_enable_value_O[0];
	assign SB_T0_WEST_SB_OUT_B17_valid_out = RMUX_T0_WEST_B17_valid_out;
	assign SB_T1_EAST_SB_IN_B17_enable = SB_T1_EAST_SB_IN_B17_enable_value_O[0];
	assign SB_T1_EAST_SB_IN_B17_ready_out = WIRE_SB_T1_EAST_SB_IN_B17_ready_out;
	assign SB_T1_EAST_SB_OUT_B17 = RMUX_T1_EAST_B17_O;
	assign SB_T1_EAST_SB_OUT_B17_enable = SB_T1_EAST_SB_OUT_B17_enable_value_O[0];
	assign SB_T1_EAST_SB_OUT_B17_valid_out = RMUX_T1_EAST_B17_valid_out;
	assign SB_T1_NORTH_SB_IN_B17_enable = SB_T1_NORTH_SB_IN_B17_enable_value_O[0];
	assign SB_T1_NORTH_SB_IN_B17_ready_out = WIRE_SB_T1_NORTH_SB_IN_B17_ready_out;
	assign SB_T1_NORTH_SB_OUT_B17 = RMUX_T1_NORTH_B17_O;
	assign SB_T1_NORTH_SB_OUT_B17_enable = SB_T1_NORTH_SB_OUT_B17_enable_value_O[0];
	assign SB_T1_NORTH_SB_OUT_B17_valid_out = RMUX_T1_NORTH_B17_valid_out;
	assign SB_T1_SOUTH_SB_IN_B17_enable = SB_T1_SOUTH_SB_IN_B17_enable_value_O[0];
	assign SB_T1_SOUTH_SB_IN_B17_ready_out = WIRE_SB_T1_SOUTH_SB_IN_B17_ready_out;
	assign SB_T1_SOUTH_SB_OUT_B17 = RMUX_T1_SOUTH_B17_O;
	assign SB_T1_SOUTH_SB_OUT_B17_enable = SB_T1_SOUTH_SB_OUT_B17_enable_value_O[0];
	assign SB_T1_SOUTH_SB_OUT_B17_valid_out = RMUX_T1_SOUTH_B17_valid_out;
	assign SB_T1_WEST_SB_IN_B17_enable = SB_T1_WEST_SB_IN_B17_enable_value_O[0];
	assign SB_T1_WEST_SB_IN_B17_ready_out = WIRE_SB_T1_WEST_SB_IN_B17_ready_out;
	assign SB_T1_WEST_SB_OUT_B17 = RMUX_T1_WEST_B17_O;
	assign SB_T1_WEST_SB_OUT_B17_enable = SB_T1_WEST_SB_OUT_B17_enable_value_O[0];
	assign SB_T1_WEST_SB_OUT_B17_valid_out = RMUX_T1_WEST_B17_valid_out;
	assign SB_T2_EAST_SB_IN_B17_enable = SB_T2_EAST_SB_IN_B17_enable_value_O[0];
	assign SB_T2_EAST_SB_IN_B17_ready_out = WIRE_SB_T2_EAST_SB_IN_B17_ready_out;
	assign SB_T2_EAST_SB_OUT_B17 = RMUX_T2_EAST_B17_O;
	assign SB_T2_EAST_SB_OUT_B17_enable = SB_T2_EAST_SB_OUT_B17_enable_value_O[0];
	assign SB_T2_EAST_SB_OUT_B17_valid_out = RMUX_T2_EAST_B17_valid_out;
	assign SB_T2_NORTH_SB_IN_B17_enable = SB_T2_NORTH_SB_IN_B17_enable_value_O[0];
	assign SB_T2_NORTH_SB_IN_B17_ready_out = WIRE_SB_T2_NORTH_SB_IN_B17_ready_out;
	assign SB_T2_NORTH_SB_OUT_B17 = RMUX_T2_NORTH_B17_O;
	assign SB_T2_NORTH_SB_OUT_B17_enable = SB_T2_NORTH_SB_OUT_B17_enable_value_O[0];
	assign SB_T2_NORTH_SB_OUT_B17_valid_out = RMUX_T2_NORTH_B17_valid_out;
	assign SB_T2_SOUTH_SB_IN_B17_enable = SB_T2_SOUTH_SB_IN_B17_enable_value_O[0];
	assign SB_T2_SOUTH_SB_IN_B17_ready_out = WIRE_SB_T2_SOUTH_SB_IN_B17_ready_out;
	assign SB_T2_SOUTH_SB_OUT_B17 = RMUX_T2_SOUTH_B17_O;
	assign SB_T2_SOUTH_SB_OUT_B17_enable = SB_T2_SOUTH_SB_OUT_B17_enable_value_O[0];
	assign SB_T2_SOUTH_SB_OUT_B17_valid_out = RMUX_T2_SOUTH_B17_valid_out;
	assign SB_T2_WEST_SB_IN_B17_enable = SB_T2_WEST_SB_IN_B17_enable_value_O[0];
	assign SB_T2_WEST_SB_IN_B17_ready_out = WIRE_SB_T2_WEST_SB_IN_B17_ready_out;
	assign SB_T2_WEST_SB_OUT_B17 = RMUX_T2_WEST_B17_O;
	assign SB_T2_WEST_SB_OUT_B17_enable = SB_T2_WEST_SB_OUT_B17_enable_value_O[0];
	assign SB_T2_WEST_SB_OUT_B17_valid_out = RMUX_T2_WEST_B17_valid_out;
	assign SB_T3_EAST_SB_IN_B17_enable = SB_T3_EAST_SB_IN_B17_enable_value_O[0];
	assign SB_T3_EAST_SB_IN_B17_ready_out = WIRE_SB_T3_EAST_SB_IN_B17_ready_out;
	assign SB_T3_EAST_SB_OUT_B17 = RMUX_T3_EAST_B17_O;
	assign SB_T3_EAST_SB_OUT_B17_enable = SB_T3_EAST_SB_OUT_B17_enable_value_O[0];
	assign SB_T3_EAST_SB_OUT_B17_valid_out = RMUX_T3_EAST_B17_valid_out;
	assign SB_T3_NORTH_SB_IN_B17_enable = SB_T3_NORTH_SB_IN_B17_enable_value_O[0];
	assign SB_T3_NORTH_SB_IN_B17_ready_out = WIRE_SB_T3_NORTH_SB_IN_B17_ready_out;
	assign SB_T3_NORTH_SB_OUT_B17 = RMUX_T3_NORTH_B17_O;
	assign SB_T3_NORTH_SB_OUT_B17_enable = SB_T3_NORTH_SB_OUT_B17_enable_value_O[0];
	assign SB_T3_NORTH_SB_OUT_B17_valid_out = RMUX_T3_NORTH_B17_valid_out;
	assign SB_T3_SOUTH_SB_IN_B17_enable = SB_T3_SOUTH_SB_IN_B17_enable_value_O[0];
	assign SB_T3_SOUTH_SB_IN_B17_ready_out = WIRE_SB_T3_SOUTH_SB_IN_B17_ready_out;
	assign SB_T3_SOUTH_SB_OUT_B17 = RMUX_T3_SOUTH_B17_O;
	assign SB_T3_SOUTH_SB_OUT_B17_enable = SB_T3_SOUTH_SB_OUT_B17_enable_value_O[0];
	assign SB_T3_SOUTH_SB_OUT_B17_valid_out = RMUX_T3_SOUTH_B17_valid_out;
	assign SB_T3_WEST_SB_IN_B17_enable = SB_T3_WEST_SB_IN_B17_enable_value_O[0];
	assign SB_T3_WEST_SB_IN_B17_ready_out = WIRE_SB_T3_WEST_SB_IN_B17_ready_out;
	assign SB_T3_WEST_SB_OUT_B17 = RMUX_T3_WEST_B17_O;
	assign SB_T3_WEST_SB_OUT_B17_enable = SB_T3_WEST_SB_OUT_B17_enable_value_O[0];
	assign SB_T3_WEST_SB_OUT_B17_valid_out = RMUX_T3_WEST_B17_valid_out;
	assign SB_T4_EAST_SB_IN_B17_enable = SB_T4_EAST_SB_IN_B17_enable_value_O[0];
	assign SB_T4_EAST_SB_IN_B17_ready_out = WIRE_SB_T4_EAST_SB_IN_B17_ready_out;
	assign SB_T4_EAST_SB_OUT_B17 = RMUX_T4_EAST_B17_O;
	assign SB_T4_EAST_SB_OUT_B17_enable = SB_T4_EAST_SB_OUT_B17_enable_value_O[0];
	assign SB_T4_EAST_SB_OUT_B17_valid_out = RMUX_T4_EAST_B17_valid_out;
	assign SB_T4_NORTH_SB_IN_B17_enable = SB_T4_NORTH_SB_IN_B17_enable_value_O[0];
	assign SB_T4_NORTH_SB_IN_B17_ready_out = WIRE_SB_T4_NORTH_SB_IN_B17_ready_out;
	assign SB_T4_NORTH_SB_OUT_B17 = RMUX_T4_NORTH_B17_O;
	assign SB_T4_NORTH_SB_OUT_B17_enable = SB_T4_NORTH_SB_OUT_B17_enable_value_O[0];
	assign SB_T4_NORTH_SB_OUT_B17_valid_out = RMUX_T4_NORTH_B17_valid_out;
	assign SB_T4_SOUTH_SB_IN_B17_enable = SB_T4_SOUTH_SB_IN_B17_enable_value_O[0];
	assign SB_T4_SOUTH_SB_IN_B17_ready_out = WIRE_SB_T4_SOUTH_SB_IN_B17_ready_out;
	assign SB_T4_SOUTH_SB_OUT_B17 = RMUX_T4_SOUTH_B17_O;
	assign SB_T4_SOUTH_SB_OUT_B17_enable = SB_T4_SOUTH_SB_OUT_B17_enable_value_O[0];
	assign SB_T4_SOUTH_SB_OUT_B17_valid_out = RMUX_T4_SOUTH_B17_valid_out;
	assign SB_T4_WEST_SB_IN_B17_enable = SB_T4_WEST_SB_IN_B17_enable_value_O[0];
	assign SB_T4_WEST_SB_IN_B17_ready_out = WIRE_SB_T4_WEST_SB_IN_B17_ready_out;
	assign SB_T4_WEST_SB_OUT_B17 = RMUX_T4_WEST_B17_O;
	assign SB_T4_WEST_SB_OUT_B17_enable = SB_T4_WEST_SB_OUT_B17_enable_value_O[0];
	assign SB_T4_WEST_SB_OUT_B17_valid_out = RMUX_T4_WEST_B17_valid_out;
	assign read_config_data = mux_aoi_6_32_inst0_O;
endmodule
module ConfigRegister_20_8_32_3 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [19:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [19:0] Register_inst0_O;
	wire [7:0] const_3_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq1 Register_inst0(
		.I(config_data[19:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h03),
		.width(8)
	) const_3_8(.out(const_3_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_3_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module PE (
	PE_input_width_17_num_0,
	PE_input_width_17_num_0_ready,
	PE_input_width_17_num_0_valid,
	PE_input_width_17_num_1,
	PE_input_width_17_num_1_ready,
	PE_input_width_17_num_1_valid,
	PE_input_width_17_num_2,
	PE_input_width_17_num_2_ready,
	PE_input_width_17_num_2_valid,
	PE_input_width_17_num_3,
	PE_input_width_17_num_3_ready,
	PE_input_width_17_num_3_valid,
	PE_input_width_1_num_0,
	PE_input_width_1_num_0_ready,
	PE_input_width_1_num_0_valid,
	PE_input_width_1_num_1,
	PE_input_width_1_num_1_ready,
	PE_input_width_1_num_1_valid,
	PE_input_width_1_num_2,
	PE_input_width_1_num_2_ready,
	PE_input_width_1_num_2_valid,
	PE_output_width_17_num_0,
	PE_output_width_17_num_0_ready,
	PE_output_width_17_num_0_valid,
	PE_output_width_17_num_1,
	PE_output_width_17_num_1_ready,
	PE_output_width_17_num_1_valid,
	PE_output_width_17_num_2,
	PE_output_width_17_num_2_ready,
	PE_output_width_17_num_2_valid,
	PE_output_width_1_num_0,
	PE_output_width_1_num_0_ready,
	PE_output_width_1_num_0_valid,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	flush,
	flush_core,
	read_config_data,
	reset,
	stall
);
	input [16:0] PE_input_width_17_num_0;
	output wire [0:0] PE_input_width_17_num_0_ready;
	input [0:0] PE_input_width_17_num_0_valid;
	input [16:0] PE_input_width_17_num_1;
	output wire [0:0] PE_input_width_17_num_1_ready;
	input [0:0] PE_input_width_17_num_1_valid;
	input [16:0] PE_input_width_17_num_2;
	output wire [0:0] PE_input_width_17_num_2_ready;
	input [0:0] PE_input_width_17_num_2_valid;
	input [16:0] PE_input_width_17_num_3;
	output wire [0:0] PE_input_width_17_num_3_ready;
	input [0:0] PE_input_width_17_num_3_valid;
	input [0:0] PE_input_width_1_num_0;
	output wire PE_input_width_1_num_0_ready;
	input PE_input_width_1_num_0_valid;
	input [0:0] PE_input_width_1_num_1;
	output wire PE_input_width_1_num_1_ready;
	input PE_input_width_1_num_1_valid;
	input [0:0] PE_input_width_1_num_2;
	output wire PE_input_width_1_num_2_ready;
	input PE_input_width_1_num_2_valid;
	output wire [16:0] PE_output_width_17_num_0;
	input [0:0] PE_output_width_17_num_0_ready;
	output wire [0:0] PE_output_width_17_num_0_valid;
	output wire [16:0] PE_output_width_17_num_1;
	input [0:0] PE_output_width_17_num_1_ready;
	output wire [0:0] PE_output_width_17_num_1_valid;
	output wire [16:0] PE_output_width_17_num_2;
	input [0:0] PE_output_width_17_num_2_ready;
	output wire [0:0] PE_output_width_17_num_2_valid;
	output wire [0:0] PE_output_width_1_num_0;
	input PE_output_width_1_num_0_ready;
	output wire PE_output_width_1_num_0_valid;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	input [0:0] flush;
	input [0:0] flush_core;
	output wire [31:0] read_config_data;
	input reset;
	input [0:0] stall;
	wire [31:0] CONFIG_SPACE_0_value_O;
	wire [31:0] CONFIG_SPACE_1_value_O;
	wire [21:0] CONFIG_SPACE_2_value_O;
	wire [0:0] Invert1_inst0_out;
	wire [0:0] Invert1_inst1_out;
	wire [16:0] PE_inner_W_inst0_PE_output_width_17_num_1;
	wire [0:0] PE_inner_W_inst0_PE_output_width_17_num_0_valid;
	wire [15:0] PE_inner_W_inst0_PE_onyx_inst_onyxpeintf_O3;
	wire [15:0] PE_inner_W_inst0_PE_onyx_inst_onyxpeintf_O4;
	wire [0:0] PE_inner_W_inst0_PE_input_width_17_num_3_ready;
	wire [0:0] PE_inner_W_inst0_PE_input_width_17_num_1_ready;
	wire [15:0] PE_inner_W_inst0_PE_onyx_inst_onyxpeintf_O2;
	wire [16:0] PE_inner_W_inst0_PE_output_width_17_num_2;
	wire [0:0] PE_inner_W_inst0_PE_input_width_17_num_0_ready;
	wire [0:0] PE_inner_W_inst0_PE_input_width_17_num_2_ready;
	wire [0:0] PE_inner_W_inst0_PE_output_width_1_num_0;
	wire [0:0] PE_inner_W_inst0_PE_output_width_17_num_1_valid;
	wire [16:0] PE_inner_W_inst0_PE_output_width_17_num_0;
	wire [0:0] PE_inner_W_inst0_PE_output_width_17_num_2_valid;
	wire [0:0] PE_input_width_17_num_0_dense_value_O;
	wire [0:0] PE_input_width_17_num_0_valid_reg_sel_value_O;
	wire [0:0] PE_input_width_17_num_0_valid_reg_value_value_O;
	wire [0:0] PE_input_width_17_num_0_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] PE_input_width_17_num_1_dense_value_O;
	wire [0:0] PE_input_width_17_num_1_valid_reg_sel_value_O;
	wire [0:0] PE_input_width_17_num_1_valid_reg_value_value_O;
	wire [0:0] PE_input_width_17_num_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] PE_input_width_17_num_2_valid_reg_sel_value_O;
	wire [0:0] PE_input_width_17_num_2_valid_reg_value_value_O;
	wire [0:0] PE_input_width_17_num_2_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] PE_input_width_17_num_3_valid_reg_sel_value_O;
	wire [0:0] PE_input_width_17_num_3_valid_reg_value_value_O;
	wire [0:0] PE_input_width_17_num_3_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] PE_input_width_1_num_0_reg_sel_value_O;
	wire [0:0] PE_input_width_1_num_0_reg_value_value_O;
	wire [0:0] PE_input_width_1_num_0_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] PE_input_width_1_num_1_reg_sel_value_O;
	wire [0:0] PE_input_width_1_num_1_reg_value_value_O;
	wire [0:0] PE_input_width_1_num_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] PE_input_width_1_num_2_reg_sel_value_O;
	wire [0:0] PE_input_width_1_num_2_reg_value_value_O;
	wire [0:0] PE_input_width_1_num_2_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [15:0] PE_onyx_inst_onyxpeintf_O2_value_O;
	wire [15:0] PE_onyx_inst_onyxpeintf_O3_value_O;
	wire [15:0] PE_onyx_inst_onyxpeintf_O4_value_O;
	wire [0:0] PE_output_width_17_num_0_dense_value_O;
	wire [0:0] PE_output_width_17_num_0_ready_reg_sel_value_O;
	wire [0:0] PE_output_width_17_num_0_ready_reg_value_value_O;
	wire [0:0] PE_output_width_17_num_0_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] PE_output_width_17_num_1_ready_reg_sel_value_O;
	wire [0:0] PE_output_width_17_num_1_ready_reg_value_value_O;
	wire [0:0] PE_output_width_17_num_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] PE_output_width_17_num_2_ready_reg_sel_value_O;
	wire [0:0] PE_output_width_17_num_2_ready_reg_value_value_O;
	wire [0:0] PE_output_width_17_num_2_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire ZextWrapper_16_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_16_32_inst0$self_O_in;
	wire ZextWrapper_16_32_inst1$bit_const_0_None_out;
	wire [31:0] ZextWrapper_16_32_inst1$self_O_in;
	wire ZextWrapper_16_32_inst2$bit_const_0_None_out;
	wire [31:0] ZextWrapper_16_32_inst2$self_O_in;
	wire ZextWrapper_20_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_20_32_inst0$self_O_in;
	wire bit_const_1_None_out;
	wire [31:0] config_reg_0_O;
	wire [31:0] config_reg_1_O;
	wire [31:0] config_reg_2_O;
	wire [19:0] config_reg_3_O;
	wire coreir_wrapInAsyncReset_inst0_out;
	wire coreir_wrapOutAsyncReset_inst0_out;
	wire [0:0] flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] flush_mux_sel_value_O;
	wire [0:0] flush_reg_sel_value_O;
	wire [0:0] flush_reg_value_value_O;
	wire [0:0] flush_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [2:0] mode_value_O;
	wire [31:0] mux_aoi_7_32_inst0_O;
	wire [7:0] mux_aoi_7_32_inst0_out_sel;
	wire [7:0] self_config_config_addr_out;
	wire [0:0] tile_en_value_O;
	SliceWrapper_32_0_32 CONFIG_SPACE_0_value(
		.I(config_reg_0_O),
		.O(CONFIG_SPACE_0_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_1_value(
		.I(config_reg_1_O),
		.O(CONFIG_SPACE_1_value_O)
	);
	SliceWrapper_32_0_22 CONFIG_SPACE_2_value(
		.I(config_reg_2_O),
		.O(CONFIG_SPACE_2_value_O)
	);
	coreir_not #(.width(1)) Invert1_inst0(
		.in(coreir_wrapInAsyncReset_inst0_out),
		.out(Invert1_inst0_out)
	);
	coreir_not #(.width(1)) Invert1_inst1(
		.in(stall),
		.out(Invert1_inst1_out)
	);
	PE_inner_W PE_inner_W_inst0(
		.PE_output_width_17_num_1(PE_inner_W_inst0_PE_output_width_17_num_1),
		.PE_output_width_17_num_0_valid(PE_inner_W_inst0_PE_output_width_17_num_0_valid),
		.PE_input_width_17_num_1_valid(PE_input_width_17_num_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.PE_input_width_17_num_1(PE_input_width_17_num_1),
		.PE_onyx_inst_onyxpeintf_O3(PE_inner_W_inst0_PE_onyx_inst_onyxpeintf_O3),
		.PE_input_width_17_num_0(PE_input_width_17_num_0),
		.PE_onyx_inst_onyxpeintf_O4(PE_inner_W_inst0_PE_onyx_inst_onyxpeintf_O4),
		.PE_input_width_17_num_0_valid(PE_input_width_17_num_0_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.clk_en(Invert1_inst1_out),
		.PE_input_width_17_num_3_ready(PE_inner_W_inst0_PE_input_width_17_num_3_ready),
		.PE_output_width_17_num_0_ready(PE_output_width_17_num_0_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.PE_input_width_17_num_1_ready(PE_inner_W_inst0_PE_input_width_17_num_1_ready),
		.PE_onyx_inst_onyxpeintf_O2(PE_inner_W_inst0_PE_onyx_inst_onyxpeintf_O2),
		.PE_input_width_17_num_1_dense(PE_input_width_17_num_1_dense_value_O),
		.PE_input_width_17_num_3_valid(PE_input_width_17_num_3_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.PE_input_width_1_num_0(PE_input_width_1_num_0_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.PE_input_width_1_num_1(PE_input_width_1_num_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.PE_output_width_17_num_0_dense(PE_output_width_17_num_0_dense_value_O),
		.PE_input_width_17_num_2(PE_input_width_17_num_2),
		.PE_output_width_17_num_2(PE_inner_W_inst0_PE_output_width_17_num_2),
		.PE_input_width_1_num_2(PE_input_width_1_num_2_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.tile_en(tile_en_value_O),
		.PE_input_width_17_num_3(PE_input_width_17_num_3),
		.PE_input_width_17_num_0_ready(PE_inner_W_inst0_PE_input_width_17_num_0_ready),
		.PE_input_width_17_num_2_valid(PE_input_width_17_num_2_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.CONFIG_SPACE_0(CONFIG_SPACE_0_value_O),
		.PE_input_width_17_num_2_ready(PE_inner_W_inst0_PE_input_width_17_num_2_ready),
		.mode(mode_value_O),
		.clk(clk),
		.flush(flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.PE_output_width_17_num_2_ready(PE_output_width_17_num_2_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.PE_output_width_1_num_0(PE_inner_W_inst0_PE_output_width_1_num_0),
		.CONFIG_SPACE_2(CONFIG_SPACE_2_value_O),
		.PE_output_width_17_num_1_valid(PE_inner_W_inst0_PE_output_width_17_num_1_valid),
		.PE_output_width_17_num_0(PE_inner_W_inst0_PE_output_width_17_num_0),
		.PE_input_width_17_num_0_dense(PE_input_width_17_num_0_dense_value_O),
		.rst_n(coreir_wrapOutAsyncReset_inst0_out),
		.CONFIG_SPACE_1(CONFIG_SPACE_1_value_O),
		.PE_output_width_17_num_1_ready(PE_output_width_17_num_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.PE_output_width_17_num_2_valid(PE_inner_W_inst0_PE_output_width_17_num_2_valid)
	);
	SliceWrapper_32_22_23 PE_input_width_17_num_0_dense_value(
		.I(config_reg_2_O),
		.O(PE_input_width_17_num_0_dense_value_O)
	);
	SliceWrapper_32_23_24 PE_input_width_17_num_0_valid_reg_sel_value(
		.I(config_reg_2_O),
		.O(PE_input_width_17_num_0_valid_reg_sel_value_O)
	);
	SliceWrapper_32_24_25 PE_input_width_17_num_0_valid_reg_value_value(
		.I(config_reg_2_O),
		.O(PE_input_width_17_num_0_valid_reg_value_value_O)
	);
	coreir_mux #(.width(1)) PE_input_width_17_num_0_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(PE_input_width_17_num_0_valid),
		.in1(PE_input_width_17_num_0_valid_reg_value_value_O),
		.sel(PE_input_width_17_num_0_valid_reg_sel_value_O[0]),
		.out(PE_input_width_17_num_0_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_32_25_26 PE_input_width_17_num_1_dense_value(
		.I(config_reg_2_O),
		.O(PE_input_width_17_num_1_dense_value_O)
	);
	SliceWrapper_32_26_27 PE_input_width_17_num_1_valid_reg_sel_value(
		.I(config_reg_2_O),
		.O(PE_input_width_17_num_1_valid_reg_sel_value_O)
	);
	SliceWrapper_32_27_28 PE_input_width_17_num_1_valid_reg_value_value(
		.I(config_reg_2_O),
		.O(PE_input_width_17_num_1_valid_reg_value_value_O)
	);
	coreir_mux #(.width(1)) PE_input_width_17_num_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(PE_input_width_17_num_1_valid),
		.in1(PE_input_width_17_num_1_valid_reg_value_value_O),
		.sel(PE_input_width_17_num_1_valid_reg_sel_value_O[0]),
		.out(PE_input_width_17_num_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_32_28_29 PE_input_width_17_num_2_valid_reg_sel_value(
		.I(config_reg_2_O),
		.O(PE_input_width_17_num_2_valid_reg_sel_value_O)
	);
	SliceWrapper_32_29_30 PE_input_width_17_num_2_valid_reg_value_value(
		.I(config_reg_2_O),
		.O(PE_input_width_17_num_2_valid_reg_value_value_O)
	);
	coreir_mux #(.width(1)) PE_input_width_17_num_2_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(PE_input_width_17_num_2_valid),
		.in1(PE_input_width_17_num_2_valid_reg_value_value_O),
		.sel(PE_input_width_17_num_2_valid_reg_sel_value_O[0]),
		.out(PE_input_width_17_num_2_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_32_30_31 PE_input_width_17_num_3_valid_reg_sel_value(
		.I(config_reg_2_O),
		.O(PE_input_width_17_num_3_valid_reg_sel_value_O)
	);
	SliceWrapper_32_31_32 PE_input_width_17_num_3_valid_reg_value_value(
		.I(config_reg_2_O),
		.O(PE_input_width_17_num_3_valid_reg_value_value_O)
	);
	coreir_mux #(.width(1)) PE_input_width_17_num_3_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(PE_input_width_17_num_3_valid),
		.in1(PE_input_width_17_num_3_valid_reg_value_value_O),
		.sel(PE_input_width_17_num_3_valid_reg_sel_value_O[0]),
		.out(PE_input_width_17_num_3_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_20_0_1 PE_input_width_1_num_0_reg_sel_value(
		.I(config_reg_3_O),
		.O(PE_input_width_1_num_0_reg_sel_value_O)
	);
	SliceWrapper_20_1_2 PE_input_width_1_num_0_reg_value_value(
		.I(config_reg_3_O),
		.O(PE_input_width_1_num_0_reg_value_value_O)
	);
	coreir_mux #(.width(1)) PE_input_width_1_num_0_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(PE_input_width_1_num_0),
		.in1(PE_input_width_1_num_0_reg_value_value_O),
		.sel(PE_input_width_1_num_0_reg_sel_value_O[0]),
		.out(PE_input_width_1_num_0_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_20_2_3 PE_input_width_1_num_1_reg_sel_value(
		.I(config_reg_3_O),
		.O(PE_input_width_1_num_1_reg_sel_value_O)
	);
	SliceWrapper_20_3_4 PE_input_width_1_num_1_reg_value_value(
		.I(config_reg_3_O),
		.O(PE_input_width_1_num_1_reg_value_value_O)
	);
	coreir_mux #(.width(1)) PE_input_width_1_num_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(PE_input_width_1_num_1),
		.in1(PE_input_width_1_num_1_reg_value_value_O),
		.sel(PE_input_width_1_num_1_reg_sel_value_O[0]),
		.out(PE_input_width_1_num_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_20_4_5 PE_input_width_1_num_2_reg_sel_value(
		.I(config_reg_3_O),
		.O(PE_input_width_1_num_2_reg_sel_value_O)
	);
	SliceWrapper_20_5_6 PE_input_width_1_num_2_reg_value_value(
		.I(config_reg_3_O),
		.O(PE_input_width_1_num_2_reg_value_value_O)
	);
	coreir_mux #(.width(1)) PE_input_width_1_num_2_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(PE_input_width_1_num_2),
		.in1(PE_input_width_1_num_2_reg_value_value_O),
		.sel(PE_input_width_1_num_2_reg_sel_value_O[0]),
		.out(PE_input_width_1_num_2_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_16_0_16 PE_onyx_inst_onyxpeintf_O2_value(
		.I(PE_inner_W_inst0_PE_onyx_inst_onyxpeintf_O2),
		.O(PE_onyx_inst_onyxpeintf_O2_value_O)
	);
	SliceWrapper_16_0_16 PE_onyx_inst_onyxpeintf_O3_value(
		.I(PE_inner_W_inst0_PE_onyx_inst_onyxpeintf_O3),
		.O(PE_onyx_inst_onyxpeintf_O3_value_O)
	);
	SliceWrapper_16_0_16 PE_onyx_inst_onyxpeintf_O4_value(
		.I(PE_inner_W_inst0_PE_onyx_inst_onyxpeintf_O4),
		.O(PE_onyx_inst_onyxpeintf_O4_value_O)
	);
	SliceWrapper_20_6_7 PE_output_width_17_num_0_dense_value(
		.I(config_reg_3_O),
		.O(PE_output_width_17_num_0_dense_value_O)
	);
	SliceWrapper_20_7_8 PE_output_width_17_num_0_ready_reg_sel_value(
		.I(config_reg_3_O),
		.O(PE_output_width_17_num_0_ready_reg_sel_value_O)
	);
	SliceWrapper_20_8_9 PE_output_width_17_num_0_ready_reg_value_value(
		.I(config_reg_3_O),
		.O(PE_output_width_17_num_0_ready_reg_value_value_O)
	);
	coreir_mux #(.width(1)) PE_output_width_17_num_0_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(PE_output_width_17_num_0_ready),
		.in1(PE_output_width_17_num_0_ready_reg_value_value_O),
		.sel(PE_output_width_17_num_0_ready_reg_sel_value_O[0]),
		.out(PE_output_width_17_num_0_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_20_9_10 PE_output_width_17_num_1_ready_reg_sel_value(
		.I(config_reg_3_O),
		.O(PE_output_width_17_num_1_ready_reg_sel_value_O)
	);
	SliceWrapper_20_10_11 PE_output_width_17_num_1_ready_reg_value_value(
		.I(config_reg_3_O),
		.O(PE_output_width_17_num_1_ready_reg_value_value_O)
	);
	coreir_mux #(.width(1)) PE_output_width_17_num_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(PE_output_width_17_num_1_ready),
		.in1(PE_output_width_17_num_1_ready_reg_value_value_O),
		.sel(PE_output_width_17_num_1_ready_reg_sel_value_O[0]),
		.out(PE_output_width_17_num_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_20_11_12 PE_output_width_17_num_2_ready_reg_sel_value(
		.I(config_reg_3_O),
		.O(PE_output_width_17_num_2_ready_reg_sel_value_O)
	);
	SliceWrapper_20_12_13 PE_output_width_17_num_2_ready_reg_value_value(
		.I(config_reg_3_O),
		.O(PE_output_width_17_num_2_ready_reg_value_value_O)
	);
	coreir_mux #(.width(1)) PE_output_width_17_num_2_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(PE_output_width_17_num_2_ready),
		.in1(PE_output_width_17_num_2_ready_reg_value_value_O),
		.sel(PE_output_width_17_num_2_ready_reg_sel_value_O[0]),
		.out(PE_output_width_17_num_2_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_16_32_inst0$bit_const_0_None(.out(ZextWrapper_16_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_16_32_inst0$self_O_out;
	assign ZextWrapper_16_32_inst0$self_O_out = {ZextWrapper_16_32_inst0$bit_const_0_None_out, ZextWrapper_16_32_inst0$bit_const_0_None_out, ZextWrapper_16_32_inst0$bit_const_0_None_out, ZextWrapper_16_32_inst0$bit_const_0_None_out, ZextWrapper_16_32_inst0$bit_const_0_None_out, ZextWrapper_16_32_inst0$bit_const_0_None_out, ZextWrapper_16_32_inst0$bit_const_0_None_out, ZextWrapper_16_32_inst0$bit_const_0_None_out, ZextWrapper_16_32_inst0$bit_const_0_None_out, ZextWrapper_16_32_inst0$bit_const_0_None_out, ZextWrapper_16_32_inst0$bit_const_0_None_out, ZextWrapper_16_32_inst0$bit_const_0_None_out, ZextWrapper_16_32_inst0$bit_const_0_None_out, ZextWrapper_16_32_inst0$bit_const_0_None_out, ZextWrapper_16_32_inst0$bit_const_0_None_out, ZextWrapper_16_32_inst0$bit_const_0_None_out, PE_onyx_inst_onyxpeintf_O3_value_O};
	mantle_wire__typeBitIn32 ZextWrapper_16_32_inst0$self_O(
		.in(ZextWrapper_16_32_inst0$self_O_in),
		.out(ZextWrapper_16_32_inst0$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_16_32_inst1$bit_const_0_None(.out(ZextWrapper_16_32_inst1$bit_const_0_None_out));
	wire [31:0] ZextWrapper_16_32_inst1$self_O_out;
	assign ZextWrapper_16_32_inst1$self_O_out = {ZextWrapper_16_32_inst1$bit_const_0_None_out, ZextWrapper_16_32_inst1$bit_const_0_None_out, ZextWrapper_16_32_inst1$bit_const_0_None_out, ZextWrapper_16_32_inst1$bit_const_0_None_out, ZextWrapper_16_32_inst1$bit_const_0_None_out, ZextWrapper_16_32_inst1$bit_const_0_None_out, ZextWrapper_16_32_inst1$bit_const_0_None_out, ZextWrapper_16_32_inst1$bit_const_0_None_out, ZextWrapper_16_32_inst1$bit_const_0_None_out, ZextWrapper_16_32_inst1$bit_const_0_None_out, ZextWrapper_16_32_inst1$bit_const_0_None_out, ZextWrapper_16_32_inst1$bit_const_0_None_out, ZextWrapper_16_32_inst1$bit_const_0_None_out, ZextWrapper_16_32_inst1$bit_const_0_None_out, ZextWrapper_16_32_inst1$bit_const_0_None_out, ZextWrapper_16_32_inst1$bit_const_0_None_out, PE_onyx_inst_onyxpeintf_O4_value_O};
	mantle_wire__typeBitIn32 ZextWrapper_16_32_inst1$self_O(
		.in(ZextWrapper_16_32_inst1$self_O_in),
		.out(ZextWrapper_16_32_inst1$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_16_32_inst2$bit_const_0_None(.out(ZextWrapper_16_32_inst2$bit_const_0_None_out));
	wire [31:0] ZextWrapper_16_32_inst2$self_O_out;
	assign ZextWrapper_16_32_inst2$self_O_out = {ZextWrapper_16_32_inst2$bit_const_0_None_out, ZextWrapper_16_32_inst2$bit_const_0_None_out, ZextWrapper_16_32_inst2$bit_const_0_None_out, ZextWrapper_16_32_inst2$bit_const_0_None_out, ZextWrapper_16_32_inst2$bit_const_0_None_out, ZextWrapper_16_32_inst2$bit_const_0_None_out, ZextWrapper_16_32_inst2$bit_const_0_None_out, ZextWrapper_16_32_inst2$bit_const_0_None_out, ZextWrapper_16_32_inst2$bit_const_0_None_out, ZextWrapper_16_32_inst2$bit_const_0_None_out, ZextWrapper_16_32_inst2$bit_const_0_None_out, ZextWrapper_16_32_inst2$bit_const_0_None_out, ZextWrapper_16_32_inst2$bit_const_0_None_out, ZextWrapper_16_32_inst2$bit_const_0_None_out, ZextWrapper_16_32_inst2$bit_const_0_None_out, ZextWrapper_16_32_inst2$bit_const_0_None_out, PE_onyx_inst_onyxpeintf_O2_value_O};
	mantle_wire__typeBitIn32 ZextWrapper_16_32_inst2$self_O(
		.in(ZextWrapper_16_32_inst2$self_O_in),
		.out(ZextWrapper_16_32_inst2$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_20_32_inst0$bit_const_0_None(.out(ZextWrapper_20_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_20_32_inst0$self_O_out;
	assign ZextWrapper_20_32_inst0$self_O_out = {ZextWrapper_20_32_inst0$bit_const_0_None_out, ZextWrapper_20_32_inst0$bit_const_0_None_out, ZextWrapper_20_32_inst0$bit_const_0_None_out, ZextWrapper_20_32_inst0$bit_const_0_None_out, ZextWrapper_20_32_inst0$bit_const_0_None_out, ZextWrapper_20_32_inst0$bit_const_0_None_out, ZextWrapper_20_32_inst0$bit_const_0_None_out, ZextWrapper_20_32_inst0$bit_const_0_None_out, ZextWrapper_20_32_inst0$bit_const_0_None_out, ZextWrapper_20_32_inst0$bit_const_0_None_out, ZextWrapper_20_32_inst0$bit_const_0_None_out, ZextWrapper_20_32_inst0$bit_const_0_None_out, config_reg_3_O};
	mantle_wire__typeBitIn32 ZextWrapper_20_32_inst0$self_O(
		.in(ZextWrapper_20_32_inst0$self_O_in),
		.out(ZextWrapper_20_32_inst0$self_O_out)
	);
	corebit_const #(.value(1'b1)) bit_const_1_None(.out(bit_const_1_None_out));
	wire [7:0] config_reg_0_config_addr;
	assign config_reg_0_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4], self_config_config_addr_out[3], self_config_config_addr_out[2:0]};
	ConfigRegister_32_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_reg_0_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_1_config_addr;
	assign config_reg_1_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4], self_config_config_addr_out[3], self_config_config_addr_out[2:0]};
	ConfigRegister_32_8_32_1 config_reg_1(
		.clk(clk),
		.reset(reset),
		.O(config_reg_1_O),
		.config_addr(config_reg_1_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_2_config_addr;
	assign config_reg_2_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4], self_config_config_addr_out[3], self_config_config_addr_out[2:0]};
	ConfigRegister_32_8_32_2 config_reg_2(
		.clk(clk),
		.reset(reset),
		.O(config_reg_2_O),
		.config_addr(config_reg_2_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_3_config_addr;
	assign config_reg_3_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4], self_config_config_addr_out[3], self_config_config_addr_out[2:0]};
	ConfigRegister_20_8_32_3 config_reg_3(
		.clk(clk),
		.reset(reset),
		.O(config_reg_3_O),
		.config_addr(config_reg_3_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	coreir_wrap coreir_wrapInAsyncReset_inst0(
		.in(reset),
		.out(coreir_wrapInAsyncReset_inst0_out)
	);
	coreir_wrap coreir_wrapOutAsyncReset_inst0(
		.in(Invert1_inst0_out[0]),
		.out(coreir_wrapOutAsyncReset_inst0_out)
	);
	coreir_mux #(.width(1)) flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(flush_core),
		.in1(flush),
		.sel(flush_mux_sel_value_O[0]),
		.out(flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_20_13_14 flush_mux_sel_value(
		.I(config_reg_3_O),
		.O(flush_mux_sel_value_O)
	);
	SliceWrapper_20_14_15 flush_reg_sel_value(
		.I(config_reg_3_O),
		.O(flush_reg_sel_value_O)
	);
	SliceWrapper_20_15_16 flush_reg_value_value(
		.I(config_reg_3_O),
		.O(flush_reg_value_value_O)
	);
	coreir_mux #(.width(1)) flush_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(flush),
		.in1(flush_reg_value_value_O),
		.sel(flush_reg_sel_value_O[0]),
		.out(flush_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_20_16_19 mode_value(
		.I(config_reg_3_O),
		.O(mode_value_O)
	);
	wire [223:0] mux_aoi_7_32_inst0_I;
	assign mux_aoi_7_32_inst0_I[192+:32] = ZextWrapper_16_32_inst2$self_O_in;
	assign mux_aoi_7_32_inst0_I[160+:32] = ZextWrapper_16_32_inst1$self_O_in;
	assign mux_aoi_7_32_inst0_I[128+:32] = ZextWrapper_16_32_inst0$self_O_in;
	assign mux_aoi_7_32_inst0_I[96+:32] = ZextWrapper_20_32_inst0$self_O_in;
	assign mux_aoi_7_32_inst0_I[64+:32] = config_reg_2_O;
	assign mux_aoi_7_32_inst0_I[32+:32] = config_reg_1_O;
	assign mux_aoi_7_32_inst0_I[0+:32] = config_reg_0_O;
	mux_aoi_7_32 mux_aoi_7_32_inst0(
		.I(mux_aoi_7_32_inst0_I),
		.O(mux_aoi_7_32_inst0_O),
		.S(self_config_config_addr_out[2:0]),
		.out_sel(mux_aoi_7_32_inst0_out_sel)
	);
	mantle_wire__typeBit8 self_config_config_addr(
		.in(config_config_addr),
		.out(self_config_config_addr_out)
	);
	SliceWrapper_20_19_20 tile_en_value(
		.I(config_reg_3_O),
		.O(tile_en_value_O)
	);
	assign PE_input_width_17_num_0_ready = PE_inner_W_inst0_PE_input_width_17_num_0_ready;
	assign PE_input_width_17_num_1_ready = PE_inner_W_inst0_PE_input_width_17_num_1_ready;
	assign PE_input_width_17_num_2_ready = PE_inner_W_inst0_PE_input_width_17_num_2_ready;
	assign PE_input_width_17_num_3_ready = PE_inner_W_inst0_PE_input_width_17_num_3_ready;
	assign PE_input_width_1_num_0_ready = bit_const_1_None_out;
	assign PE_input_width_1_num_1_ready = bit_const_1_None_out;
	assign PE_input_width_1_num_2_ready = bit_const_1_None_out;
	assign PE_output_width_17_num_0 = PE_inner_W_inst0_PE_output_width_17_num_0;
	assign PE_output_width_17_num_0_valid = PE_inner_W_inst0_PE_output_width_17_num_0_valid;
	assign PE_output_width_17_num_1 = PE_inner_W_inst0_PE_output_width_17_num_1;
	assign PE_output_width_17_num_1_valid = PE_inner_W_inst0_PE_output_width_17_num_1_valid;
	assign PE_output_width_17_num_2 = PE_inner_W_inst0_PE_output_width_17_num_2;
	assign PE_output_width_17_num_2_valid = PE_inner_W_inst0_PE_output_width_17_num_2_valid;
	assign PE_output_width_1_num_0 = PE_inner_W_inst0_PE_output_width_1_num_0;
	assign PE_output_width_1_num_0_valid = bit_const_1_None_out;
	assign read_config_data = mux_aoi_7_32_inst0_O;
endmodule
module ConfigRegister_1_8_32_17 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [0:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [0:0] Register_inst0_O;
	wire [7:0] const_17_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq4 Register_inst0(
		.I(config_data[0:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h11),
		.width(8)
	) const_17_8(.out(const_17_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_17_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module PondCore (
	PondTop_input_width_17_num_0,
	PondTop_input_width_17_num_0_ready,
	PondTop_input_width_17_num_0_valid,
	PondTop_input_width_17_num_1,
	PondTop_input_width_17_num_1_ready,
	PondTop_input_width_17_num_1_valid,
	PondTop_output_width_17_num_0,
	PondTop_output_width_17_num_0_ready,
	PondTop_output_width_17_num_0_valid,
	PondTop_output_width_17_num_1,
	PondTop_output_width_17_num_1_ready,
	PondTop_output_width_17_num_1_valid,
	PondTop_output_width_1_num_0,
	PondTop_output_width_1_num_0_ready,
	PondTop_output_width_1_num_0_valid,
	PondTop_output_width_1_num_1,
	PondTop_output_width_1_num_1_ready,
	PondTop_output_width_1_num_1_valid,
	clk,
	config_1_config_addr,
	config_1_config_data,
	config_1_read,
	config_1_write,
	config_config_addr,
	config_config_data,
	config_en_0,
	config_read,
	config_write,
	flush,
	flush_core,
	read_config_data,
	read_config_data_1,
	reset,
	stall
);
	input [16:0] PondTop_input_width_17_num_0;
	output wire PondTop_input_width_17_num_0_ready;
	input PondTop_input_width_17_num_0_valid;
	input [16:0] PondTop_input_width_17_num_1;
	output wire PondTop_input_width_17_num_1_ready;
	input PondTop_input_width_17_num_1_valid;
	output wire [16:0] PondTop_output_width_17_num_0;
	input PondTop_output_width_17_num_0_ready;
	output wire PondTop_output_width_17_num_0_valid;
	output wire [16:0] PondTop_output_width_17_num_1;
	input PondTop_output_width_17_num_1_ready;
	output wire PondTop_output_width_17_num_1_valid;
	output wire [0:0] PondTop_output_width_1_num_0;
	input PondTop_output_width_1_num_0_ready;
	output wire PondTop_output_width_1_num_0_valid;
	output wire [0:0] PondTop_output_width_1_num_1;
	input PondTop_output_width_1_num_1_ready;
	output wire PondTop_output_width_1_num_1_valid;
	input clk;
	input [7:0] config_1_config_addr;
	input [31:0] config_1_config_data;
	input [0:0] config_1_read;
	input [0:0] config_1_write;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input config_en_0;
	input [0:0] config_read;
	input [0:0] config_write;
	input [0:0] flush;
	input [0:0] flush_core;
	output wire [31:0] read_config_data;
	output wire [31:0] read_config_data_1;
	input reset;
	input [0:0] stall;
	wire [0:0] AND_CONFIG_EN_SRAM_0_out;
	wire [31:0] CONFIG_SPACE_0_value_O;
	wire [31:0] CONFIG_SPACE_10_value_O;
	wire [31:0] CONFIG_SPACE_11_value_O;
	wire [31:0] CONFIG_SPACE_12_value_O;
	wire [31:0] CONFIG_SPACE_13_value_O;
	wire [31:0] CONFIG_SPACE_14_value_O;
	wire [31:0] CONFIG_SPACE_15_value_O;
	wire [29:0] CONFIG_SPACE_16_value_O;
	wire [31:0] CONFIG_SPACE_1_value_O;
	wire [31:0] CONFIG_SPACE_2_value_O;
	wire [31:0] CONFIG_SPACE_3_value_O;
	wire [31:0] CONFIG_SPACE_4_value_O;
	wire [31:0] CONFIG_SPACE_5_value_O;
	wire [31:0] CONFIG_SPACE_6_value_O;
	wire [31:0] CONFIG_SPACE_7_value_O;
	wire [31:0] CONFIG_SPACE_8_value_O;
	wire [31:0] CONFIG_SPACE_9_value_O;
	wire [0:0] Invert1_inst0_out;
	wire [0:0] Invert1_inst1_out;
	wire [0:0] OR_CONFIG_EN_SRAM_0_out;
	wire OR_CONFIG_RD_SRAM$orr_inst0_out;
	wire OR_CONFIG_WR_SRAM$orr_inst0_out;
	wire [7:0] OR_config_addr_FEATURE_out;
	wire [31:0] OR_config_data_FEATURE_out;
	wire [0:0] PondTop_W_inst0_PondTop_output_width_1_num_1;
	wire [0:0] PondTop_W_inst0_PondTop_output_width_1_num_0;
	wire [16:0] PondTop_W_inst0_PondTop_output_width_17_num_1;
	wire [31:0] PondTop_W_inst0_config_data_out;
	wire [16:0] PondTop_W_inst0_PondTop_output_width_17_num_0;
	wire ZextWrapper_1_32_inst0$bit_const_0_None_out;
	wire ZextWrapper_30_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_30_32_inst0$self_O_in;
	wire bit_const_1_None_out;
	wire [31:0] config_reg_0_O;
	wire [31:0] config_reg_1_O;
	wire [31:0] config_reg_10_O;
	wire [31:0] config_reg_11_O;
	wire [31:0] config_reg_12_O;
	wire [31:0] config_reg_13_O;
	wire [31:0] config_reg_14_O;
	wire [31:0] config_reg_15_O;
	wire [31:0] config_reg_16_O;
	wire [0:0] config_reg_17_O;
	wire [31:0] config_reg_2_O;
	wire [31:0] config_reg_3_O;
	wire [31:0] config_reg_4_O;
	wire [31:0] config_reg_5_O;
	wire [31:0] config_reg_6_O;
	wire [31:0] config_reg_7_O;
	wire [29:0] config_reg_8_O;
	wire [31:0] config_reg_9_O;
	wire coreir_wrapInAsyncReset_inst0_out;
	wire coreir_wrapOutAsyncReset_inst0_out;
	wire [31:0] mux_aoi_18_32_inst0_O;
	wire [31:0] mux_aoi_18_32_inst0_out_sel;
	wire [0:0] or1_inst0_out;
	wire [7:0] self_config_config_addr_out;
	wire [0:0] tile_en_value_O;
	coreir_and #(.width(1)) AND_CONFIG_EN_SRAM_0(
		.in0(OR_CONFIG_EN_SRAM_0_out),
		.in1(config_en_0),
		.out(AND_CONFIG_EN_SRAM_0_out)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_0_value(
		.I(config_reg_0_O),
		.O(CONFIG_SPACE_0_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_10_value(
		.I(config_reg_2_O),
		.O(CONFIG_SPACE_10_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_11_value(
		.I(config_reg_3_O),
		.O(CONFIG_SPACE_11_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_12_value(
		.I(config_reg_4_O),
		.O(CONFIG_SPACE_12_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_13_value(
		.I(config_reg_5_O),
		.O(CONFIG_SPACE_13_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_14_value(
		.I(config_reg_6_O),
		.O(CONFIG_SPACE_14_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_15_value(
		.I(config_reg_7_O),
		.O(CONFIG_SPACE_15_value_O)
	);
	SliceWrapper_30_0_30 CONFIG_SPACE_16_value(
		.I(config_reg_8_O),
		.O(CONFIG_SPACE_16_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_1_value(
		.I(config_reg_1_O),
		.O(CONFIG_SPACE_1_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_2_value(
		.I(config_reg_9_O),
		.O(CONFIG_SPACE_2_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_3_value(
		.I(config_reg_10_O),
		.O(CONFIG_SPACE_3_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_4_value(
		.I(config_reg_11_O),
		.O(CONFIG_SPACE_4_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_5_value(
		.I(config_reg_12_O),
		.O(CONFIG_SPACE_5_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_6_value(
		.I(config_reg_13_O),
		.O(CONFIG_SPACE_6_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_7_value(
		.I(config_reg_14_O),
		.O(CONFIG_SPACE_7_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_8_value(
		.I(config_reg_15_O),
		.O(CONFIG_SPACE_8_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_9_value(
		.I(config_reg_16_O),
		.O(CONFIG_SPACE_9_value_O)
	);
	coreir_not #(.width(1)) Invert1_inst0(
		.in(coreir_wrapInAsyncReset_inst0_out),
		.out(Invert1_inst0_out)
	);
	coreir_not #(.width(1)) Invert1_inst1(
		.in(stall),
		.out(Invert1_inst1_out)
	);
	coreir_or #(.width(1)) OR_CONFIG_EN_SRAM_0(
		.in0(config_1_write),
		.in1(config_1_read),
		.out(OR_CONFIG_EN_SRAM_0_out)
	);
	coreir_orr #(.width(1)) OR_CONFIG_RD_SRAM$orr_inst0(
		.in(config_1_write),
		.out(OR_CONFIG_RD_SRAM$orr_inst0_out)
	);
	coreir_orr #(.width(1)) OR_CONFIG_WR_SRAM$orr_inst0(
		.in(config_1_read),
		.out(OR_CONFIG_WR_SRAM$orr_inst0_out)
	);
	wire [7:0] OR_config_addr_FEATURE_in0;
	assign OR_config_addr_FEATURE_in0 = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4:0]};
	coreir_or #(.width(8)) OR_config_addr_FEATURE(
		.in0(OR_config_addr_FEATURE_in0),
		.in1(config_1_config_addr),
		.out(OR_config_addr_FEATURE_out)
	);
	coreir_or #(.width(32)) OR_config_data_FEATURE(
		.in0(config_config_data),
		.in1(config_1_config_data),
		.out(OR_config_data_FEATURE_out)
	);
	PondTop_W PondTop_W_inst0(
		.CONFIG_SPACE_7(CONFIG_SPACE_7_value_O),
		.PondTop_input_width_17_num_0(PondTop_input_width_17_num_0),
		.CONFIG_SPACE_5(CONFIG_SPACE_5_value_O),
		.clk_en(Invert1_inst1_out),
		.CONFIG_SPACE_14(CONFIG_SPACE_14_value_O),
		.CONFIG_SPACE_11(CONFIG_SPACE_11_value_O),
		.config_write(OR_CONFIG_RD_SRAM$orr_inst0_out),
		.PondTop_output_width_1_num_1(PondTop_W_inst0_PondTop_output_width_1_num_1),
		.tile_en(tile_en_value_O),
		.config_en(AND_CONFIG_EN_SRAM_0_out),
		.PondTop_input_width_17_num_1(PondTop_input_width_17_num_1),
		.config_data_in(OR_config_data_FEATURE_out),
		.CONFIG_SPACE_0(CONFIG_SPACE_0_value_O),
		.PondTop_output_width_1_num_0(PondTop_W_inst0_PondTop_output_width_1_num_0),
		.CONFIG_SPACE_10(CONFIG_SPACE_10_value_O),
		.CONFIG_SPACE_9(CONFIG_SPACE_9_value_O),
		.clk(clk),
		.flush(or1_inst0_out),
		.CONFIG_SPACE_8(CONFIG_SPACE_8_value_O),
		.CONFIG_SPACE_16(CONFIG_SPACE_16_value_O),
		.CONFIG_SPACE_6(CONFIG_SPACE_6_value_O),
		.PondTop_output_width_17_num_1(PondTop_W_inst0_PondTop_output_width_17_num_1),
		.CONFIG_SPACE_2(CONFIG_SPACE_2_value_O),
		.CONFIG_SPACE_4(CONFIG_SPACE_4_value_O),
		.config_data_out(PondTop_W_inst0_config_data_out),
		.CONFIG_SPACE_13(CONFIG_SPACE_13_value_O),
		.CONFIG_SPACE_3(CONFIG_SPACE_3_value_O),
		.PondTop_output_width_17_num_0(PondTop_W_inst0_PondTop_output_width_17_num_0),
		.CONFIG_SPACE_15(CONFIG_SPACE_15_value_O),
		.CONFIG_SPACE_12(CONFIG_SPACE_12_value_O),
		.config_addr_in(OR_config_addr_FEATURE_out),
		.rst_n(coreir_wrapOutAsyncReset_inst0_out),
		.CONFIG_SPACE_1(CONFIG_SPACE_1_value_O),
		.config_read(OR_CONFIG_WR_SRAM$orr_inst0_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_1_32_inst0$bit_const_0_None(.out(ZextWrapper_1_32_inst0$bit_const_0_None_out));
	corebit_const #(.value(1'b0)) ZextWrapper_30_32_inst0$bit_const_0_None(.out(ZextWrapper_30_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_30_32_inst0$self_O_out;
	assign ZextWrapper_30_32_inst0$self_O_out = {ZextWrapper_30_32_inst0$bit_const_0_None_out, ZextWrapper_30_32_inst0$bit_const_0_None_out, config_reg_8_O};
	mantle_wire__typeBitIn32 ZextWrapper_30_32_inst0$self_O(
		.in(ZextWrapper_30_32_inst0$self_O_in),
		.out(ZextWrapper_30_32_inst0$self_O_out)
	);
	corebit_const #(.value(1'b1)) bit_const_1_None(.out(bit_const_1_None_out));
	wire [7:0] config_reg_0_config_addr;
	assign config_reg_0_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4:0]};
	ConfigRegister_32_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_reg_0_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_1_config_addr;
	assign config_reg_1_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4:0]};
	ConfigRegister_32_8_32_1 config_reg_1(
		.clk(clk),
		.reset(reset),
		.O(config_reg_1_O),
		.config_addr(config_reg_1_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_10_config_addr;
	assign config_reg_10_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4:0]};
	ConfigRegister_32_8_32_10 config_reg_10(
		.clk(clk),
		.reset(reset),
		.O(config_reg_10_O),
		.config_addr(config_reg_10_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_11_config_addr;
	assign config_reg_11_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4:0]};
	ConfigRegister_32_8_32_11 config_reg_11(
		.clk(clk),
		.reset(reset),
		.O(config_reg_11_O),
		.config_addr(config_reg_11_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_12_config_addr;
	assign config_reg_12_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4:0]};
	ConfigRegister_32_8_32_12 config_reg_12(
		.clk(clk),
		.reset(reset),
		.O(config_reg_12_O),
		.config_addr(config_reg_12_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_13_config_addr;
	assign config_reg_13_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4:0]};
	ConfigRegister_32_8_32_13 config_reg_13(
		.clk(clk),
		.reset(reset),
		.O(config_reg_13_O),
		.config_addr(config_reg_13_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_14_config_addr;
	assign config_reg_14_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4:0]};
	ConfigRegister_32_8_32_14 config_reg_14(
		.clk(clk),
		.reset(reset),
		.O(config_reg_14_O),
		.config_addr(config_reg_14_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_15_config_addr;
	assign config_reg_15_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4:0]};
	ConfigRegister_32_8_32_15 config_reg_15(
		.clk(clk),
		.reset(reset),
		.O(config_reg_15_O),
		.config_addr(config_reg_15_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_16_config_addr;
	assign config_reg_16_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4:0]};
	ConfigRegister_32_8_32_16 config_reg_16(
		.clk(clk),
		.reset(reset),
		.O(config_reg_16_O),
		.config_addr(config_reg_16_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_17_config_addr;
	assign config_reg_17_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4:0]};
	ConfigRegister_1_8_32_17 config_reg_17(
		.clk(clk),
		.reset(reset),
		.O(config_reg_17_O),
		.config_addr(config_reg_17_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_2_config_addr;
	assign config_reg_2_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4:0]};
	ConfigRegister_32_8_32_2 config_reg_2(
		.clk(clk),
		.reset(reset),
		.O(config_reg_2_O),
		.config_addr(config_reg_2_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_3_config_addr;
	assign config_reg_3_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4:0]};
	ConfigRegister_32_8_32_3 config_reg_3(
		.clk(clk),
		.reset(reset),
		.O(config_reg_3_O),
		.config_addr(config_reg_3_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_4_config_addr;
	assign config_reg_4_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4:0]};
	ConfigRegister_32_8_32_4 config_reg_4(
		.clk(clk),
		.reset(reset),
		.O(config_reg_4_O),
		.config_addr(config_reg_4_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_5_config_addr;
	assign config_reg_5_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4:0]};
	ConfigRegister_32_8_32_5 config_reg_5(
		.clk(clk),
		.reset(reset),
		.O(config_reg_5_O),
		.config_addr(config_reg_5_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_6_config_addr;
	assign config_reg_6_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4:0]};
	ConfigRegister_32_8_32_6 config_reg_6(
		.clk(clk),
		.reset(reset),
		.O(config_reg_6_O),
		.config_addr(config_reg_6_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_7_config_addr;
	assign config_reg_7_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4:0]};
	ConfigRegister_32_8_32_7 config_reg_7(
		.clk(clk),
		.reset(reset),
		.O(config_reg_7_O),
		.config_addr(config_reg_7_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_8_config_addr;
	assign config_reg_8_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4:0]};
	ConfigRegister_30_8_32_8 config_reg_8(
		.clk(clk),
		.reset(reset),
		.O(config_reg_8_O),
		.config_addr(config_reg_8_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_9_config_addr;
	assign config_reg_9_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5], self_config_config_addr_out[4:0]};
	ConfigRegister_32_8_32_9 config_reg_9(
		.clk(clk),
		.reset(reset),
		.O(config_reg_9_O),
		.config_addr(config_reg_9_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	coreir_wrap coreir_wrapInAsyncReset_inst0(
		.in(reset),
		.out(coreir_wrapInAsyncReset_inst0_out)
	);
	coreir_wrap coreir_wrapOutAsyncReset_inst0(
		.in(Invert1_inst0_out[0]),
		.out(coreir_wrapOutAsyncReset_inst0_out)
	);
	wire [575:0] mux_aoi_18_32_inst0_I;
	assign mux_aoi_18_32_inst0_I[544+:32] = {ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, config_reg_17_O[0]};
	assign mux_aoi_18_32_inst0_I[512+:32] = config_reg_16_O;
	assign mux_aoi_18_32_inst0_I[480+:32] = config_reg_15_O;
	assign mux_aoi_18_32_inst0_I[448+:32] = config_reg_14_O;
	assign mux_aoi_18_32_inst0_I[416+:32] = config_reg_13_O;
	assign mux_aoi_18_32_inst0_I[384+:32] = config_reg_12_O;
	assign mux_aoi_18_32_inst0_I[352+:32] = config_reg_11_O;
	assign mux_aoi_18_32_inst0_I[320+:32] = config_reg_10_O;
	assign mux_aoi_18_32_inst0_I[288+:32] = config_reg_9_O;
	assign mux_aoi_18_32_inst0_I[256+:32] = ZextWrapper_30_32_inst0$self_O_in;
	assign mux_aoi_18_32_inst0_I[224+:32] = config_reg_7_O;
	assign mux_aoi_18_32_inst0_I[192+:32] = config_reg_6_O;
	assign mux_aoi_18_32_inst0_I[160+:32] = config_reg_5_O;
	assign mux_aoi_18_32_inst0_I[128+:32] = config_reg_4_O;
	assign mux_aoi_18_32_inst0_I[96+:32] = config_reg_3_O;
	assign mux_aoi_18_32_inst0_I[64+:32] = config_reg_2_O;
	assign mux_aoi_18_32_inst0_I[32+:32] = config_reg_1_O;
	assign mux_aoi_18_32_inst0_I[0+:32] = config_reg_0_O;
	mux_aoi_18_32 mux_aoi_18_32_inst0(
		.I(mux_aoi_18_32_inst0_I),
		.O(mux_aoi_18_32_inst0_O),
		.S(self_config_config_addr_out[4:0]),
		.out_sel(mux_aoi_18_32_inst0_out_sel)
	);
	coreir_or #(.width(1)) or1_inst0(
		.in0(flush_core),
		.in1(flush),
		.out(or1_inst0_out)
	);
	mantle_wire__typeBit8 self_config_config_addr(
		.in(config_config_addr),
		.out(self_config_config_addr_out)
	);
	SliceWrapper_1_0_1 tile_en_value(
		.I(config_reg_17_O),
		.O(tile_en_value_O)
	);
	assign PondTop_input_width_17_num_0_ready = bit_const_1_None_out;
	assign PondTop_input_width_17_num_1_ready = bit_const_1_None_out;
	assign PondTop_output_width_17_num_0 = PondTop_W_inst0_PondTop_output_width_17_num_0;
	assign PondTop_output_width_17_num_0_valid = bit_const_1_None_out;
	assign PondTop_output_width_17_num_1 = PondTop_W_inst0_PondTop_output_width_17_num_1;
	assign PondTop_output_width_17_num_1_valid = bit_const_1_None_out;
	assign PondTop_output_width_1_num_0 = PondTop_W_inst0_PondTop_output_width_1_num_0;
	assign PondTop_output_width_1_num_0_valid = bit_const_1_None_out;
	assign PondTop_output_width_1_num_1 = PondTop_W_inst0_PondTop_output_width_1_num_1;
	assign PondTop_output_width_1_num_1_valid = bit_const_1_None_out;
	assign read_config_data = mux_aoi_18_32_inst0_O;
	assign read_config_data_1 = PondTop_W_inst0_config_data_out;
endmodule
module ConfigRegister_1_8_32_0 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [0:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [0:0] Register_inst0_O;
	wire [7:0] const_0_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq4 Register_inst0(
		.I(config_data[0:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h00),
		.width(8)
	) const_0_8(.out(const_0_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_0_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module PowerDomainConfigReg (
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	ps_en_out,
	read_config_data,
	reset
);
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output wire [0:0] ps_en_out;
	output wire [31:0] read_config_data;
	input reset;
	wire ZextWrapper_1_32_inst0$bit_const_0_None_out;
	wire [0:0] config_reg_0_O;
	wire [0:0] ps_en_value_O;
	corebit_const #(.value(1'b0)) ZextWrapper_1_32_inst0$bit_const_0_None(.out(ZextWrapper_1_32_inst0$bit_const_0_None_out));
	ConfigRegister_1_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	SliceWrapper_1_0_1 ps_en_value(
		.I(config_reg_0_O),
		.O(ps_en_value_O)
	);
	assign ps_en_out = ps_en_value_O;
	assign read_config_data = {ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, ZextWrapper_1_32_inst0$bit_const_0_None_out, config_reg_0_O[0]};
endmodule
module ConfigRegister_19_8_32_40 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output wire [18:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [18:0] Register_inst0_O;
	wire [7:0] const_40_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq7 Register_inst0(
		.I(config_data[18:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h28),
		.width(8)
	) const_40_8(.out(const_40_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_40_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module MemCore (
	MEM_input_width_17_num_0,
	MEM_input_width_17_num_0_ready,
	MEM_input_width_17_num_0_valid,
	MEM_input_width_17_num_1,
	MEM_input_width_17_num_1_ready,
	MEM_input_width_17_num_1_valid,
	MEM_input_width_17_num_2,
	MEM_input_width_17_num_2_ready,
	MEM_input_width_17_num_2_valid,
	MEM_input_width_17_num_3,
	MEM_input_width_17_num_3_ready,
	MEM_input_width_17_num_3_valid,
	MEM_input_width_1_num_0,
	MEM_input_width_1_num_0_ready,
	MEM_input_width_1_num_0_valid,
	MEM_input_width_1_num_1,
	MEM_input_width_1_num_1_ready,
	MEM_input_width_1_num_1_valid,
	MEM_output_width_17_num_0,
	MEM_output_width_17_num_0_ready,
	MEM_output_width_17_num_0_valid,
	MEM_output_width_17_num_1,
	MEM_output_width_17_num_1_ready,
	MEM_output_width_17_num_1_valid,
	MEM_output_width_17_num_2,
	MEM_output_width_17_num_2_ready,
	MEM_output_width_17_num_2_valid,
	MEM_output_width_1_num_0,
	MEM_output_width_1_num_0_ready,
	MEM_output_width_1_num_0_valid,
	MEM_output_width_1_num_1,
	MEM_output_width_1_num_1_ready,
	MEM_output_width_1_num_1_valid,
	MEM_output_width_1_num_2,
	MEM_output_width_1_num_2_ready,
	MEM_output_width_1_num_2_valid,
	clk,
	config_1_config_addr,
	config_1_config_data,
	config_1_read,
	config_1_write,
	config_2_config_addr,
	config_2_config_data,
	config_2_read,
	config_2_write,
	config_config_addr,
	config_config_data,
	config_en_0,
	config_en_1,
	config_read,
	config_write,
	flush,
	flush_core,
	read_config_data,
	read_config_data_1,
	read_config_data_2,
	reset,
	stall
);
	input [16:0] MEM_input_width_17_num_0;
	output wire [0:0] MEM_input_width_17_num_0_ready;
	input [0:0] MEM_input_width_17_num_0_valid;
	input [16:0] MEM_input_width_17_num_1;
	output wire [0:0] MEM_input_width_17_num_1_ready;
	input [0:0] MEM_input_width_17_num_1_valid;
	input [16:0] MEM_input_width_17_num_2;
	output wire [0:0] MEM_input_width_17_num_2_ready;
	input [0:0] MEM_input_width_17_num_2_valid;
	input [16:0] MEM_input_width_17_num_3;
	output wire [0:0] MEM_input_width_17_num_3_ready;
	input [0:0] MEM_input_width_17_num_3_valid;
	input [0:0] MEM_input_width_1_num_0;
	output wire MEM_input_width_1_num_0_ready;
	input MEM_input_width_1_num_0_valid;
	input [0:0] MEM_input_width_1_num_1;
	output wire MEM_input_width_1_num_1_ready;
	input MEM_input_width_1_num_1_valid;
	output wire [16:0] MEM_output_width_17_num_0;
	input [0:0] MEM_output_width_17_num_0_ready;
	output wire [0:0] MEM_output_width_17_num_0_valid;
	output wire [16:0] MEM_output_width_17_num_1;
	input [0:0] MEM_output_width_17_num_1_ready;
	output wire [0:0] MEM_output_width_17_num_1_valid;
	output wire [16:0] MEM_output_width_17_num_2;
	input [0:0] MEM_output_width_17_num_2_ready;
	output wire [0:0] MEM_output_width_17_num_2_valid;
	output wire [0:0] MEM_output_width_1_num_0;
	input MEM_output_width_1_num_0_ready;
	output wire MEM_output_width_1_num_0_valid;
	output wire [0:0] MEM_output_width_1_num_1;
	input MEM_output_width_1_num_1_ready;
	output wire MEM_output_width_1_num_1_valid;
	output wire [0:0] MEM_output_width_1_num_2;
	input MEM_output_width_1_num_2_ready;
	output wire MEM_output_width_1_num_2_valid;
	input clk;
	input [7:0] config_1_config_addr;
	input [31:0] config_1_config_data;
	input [0:0] config_1_read;
	input [0:0] config_1_write;
	input [7:0] config_2_config_addr;
	input [31:0] config_2_config_data;
	input [0:0] config_2_read;
	input [0:0] config_2_write;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input config_en_0;
	input config_en_1;
	input [0:0] config_read;
	input [0:0] config_write;
	input [0:0] flush;
	input [0:0] flush_core;
	output wire [31:0] read_config_data;
	output wire [31:0] read_config_data_1;
	output wire [31:0] read_config_data_2;
	input reset;
	input [0:0] stall;
	wire [0:0] AND_CONFIG_EN_SRAM_0_out;
	wire [0:0] AND_CONFIG_EN_SRAM_1_out;
	wire [31:0] CONFIG_SPACE_0_value_O;
	wire [31:0] CONFIG_SPACE_10_value_O;
	wire [31:0] CONFIG_SPACE_11_value_O;
	wire [31:0] CONFIG_SPACE_12_value_O;
	wire [31:0] CONFIG_SPACE_13_value_O;
	wire [31:0] CONFIG_SPACE_14_value_O;
	wire [31:0] CONFIG_SPACE_15_value_O;
	wire [31:0] CONFIG_SPACE_16_value_O;
	wire [31:0] CONFIG_SPACE_17_value_O;
	wire [31:0] CONFIG_SPACE_18_value_O;
	wire [31:0] CONFIG_SPACE_19_value_O;
	wire [31:0] CONFIG_SPACE_1_value_O;
	wire [31:0] CONFIG_SPACE_20_value_O;
	wire [31:0] CONFIG_SPACE_21_value_O;
	wire [31:0] CONFIG_SPACE_22_value_O;
	wire [31:0] CONFIG_SPACE_23_value_O;
	wire [31:0] CONFIG_SPACE_24_value_O;
	wire [31:0] CONFIG_SPACE_25_value_O;
	wire [31:0] CONFIG_SPACE_26_value_O;
	wire [31:0] CONFIG_SPACE_27_value_O;
	wire [31:0] CONFIG_SPACE_28_value_O;
	wire [31:0] CONFIG_SPACE_29_value_O;
	wire [31:0] CONFIG_SPACE_2_value_O;
	wire [31:0] CONFIG_SPACE_30_value_O;
	wire [31:0] CONFIG_SPACE_31_value_O;
	wire [31:0] CONFIG_SPACE_32_value_O;
	wire [31:0] CONFIG_SPACE_33_value_O;
	wire [31:0] CONFIG_SPACE_34_value_O;
	wire [31:0] CONFIG_SPACE_35_value_O;
	wire [31:0] CONFIG_SPACE_36_value_O;
	wire [31:0] CONFIG_SPACE_37_value_O;
	wire [31:0] CONFIG_SPACE_38_value_O;
	wire [31:0] CONFIG_SPACE_39_value_O;
	wire [31:0] CONFIG_SPACE_3_value_O;
	wire [31:0] CONFIG_SPACE_40_value_O;
	wire [31:0] CONFIG_SPACE_41_value_O;
	wire [31:0] CONFIG_SPACE_42_value_O;
	wire [31:0] CONFIG_SPACE_43_value_O;
	wire [31:0] CONFIG_SPACE_44_value_O;
	wire [18:0] CONFIG_SPACE_45_value_O;
	wire [31:0] CONFIG_SPACE_4_value_O;
	wire [31:0] CONFIG_SPACE_5_value_O;
	wire [31:0] CONFIG_SPACE_6_value_O;
	wire [31:0] CONFIG_SPACE_7_value_O;
	wire [31:0] CONFIG_SPACE_8_value_O;
	wire [31:0] CONFIG_SPACE_9_value_O;
	wire [0:0] Invert1_inst0_out;
	wire [0:0] Invert1_inst1_out;
	wire [0:0] MEM_input_width_17_num_0_valid_reg_sel_value_O;
	wire [0:0] MEM_input_width_17_num_0_valid_reg_value_value_O;
	wire [0:0] MEM_input_width_17_num_0_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] MEM_input_width_17_num_1_valid_reg_sel_value_O;
	wire [0:0] MEM_input_width_17_num_1_valid_reg_value_value_O;
	wire [0:0] MEM_input_width_17_num_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] MEM_input_width_17_num_2_valid_reg_sel_value_O;
	wire [0:0] MEM_input_width_17_num_2_valid_reg_value_value_O;
	wire [0:0] MEM_input_width_17_num_2_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] MEM_input_width_17_num_3_valid_reg_sel_value_O;
	wire [0:0] MEM_input_width_17_num_3_valid_reg_value_value_O;
	wire [0:0] MEM_input_width_17_num_3_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] MEM_input_width_1_num_0_reg_sel_value_O;
	wire [0:0] MEM_input_width_1_num_0_reg_value_value_O;
	wire [0:0] MEM_input_width_1_num_0_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] MEM_input_width_1_num_1_reg_sel_value_O;
	wire [0:0] MEM_input_width_1_num_1_reg_value_value_O;
	wire [0:0] MEM_input_width_1_num_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] MEM_output_width_17_num_0_ready_reg_sel_value_O;
	wire [0:0] MEM_output_width_17_num_0_ready_reg_value_value_O;
	wire [0:0] MEM_output_width_17_num_0_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] MEM_output_width_17_num_1_ready_reg_sel_value_O;
	wire [0:0] MEM_output_width_17_num_1_ready_reg_value_value_O;
	wire [0:0] MEM_output_width_17_num_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] MEM_output_width_17_num_2_ready_reg_sel_value_O;
	wire [0:0] MEM_output_width_17_num_2_ready_reg_value_value_O;
	wire [0:0] MEM_output_width_17_num_2_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [31:0] MemCore_inner_W_inst0_config_data_out_1;
	wire [31:0] MemCore_inner_W_inst0_config_data_out_0;
	wire [0:0] MemCore_inner_W_inst0_MEM_input_width_17_num_3_ready;
	wire [0:0] MemCore_inner_W_inst0_MEM_output_width_1_num_2;
	wire [0:0] MemCore_inner_W_inst0_MEM_output_width_1_num_1;
	wire [0:0] MemCore_inner_W_inst0_MEM_output_width_17_num_1_valid;
	wire [16:0] MemCore_inner_W_inst0_MEM_output_width_17_num_2;
	wire [0:0] MemCore_inner_W_inst0_MEM_input_width_17_num_2_ready;
	wire [16:0] MemCore_inner_W_inst0_MEM_output_width_17_num_1;
	wire [0:0] MemCore_inner_W_inst0_MEM_output_width_1_num_0;
	wire [0:0] MemCore_inner_W_inst0_MEM_output_width_17_num_2_valid;
	wire [0:0] MemCore_inner_W_inst0_MEM_input_width_17_num_1_ready;
	wire [0:0] MemCore_inner_W_inst0_MEM_input_width_17_num_0_ready;
	wire [0:0] MemCore_inner_W_inst0_MEM_output_width_17_num_0_valid;
	wire [16:0] MemCore_inner_W_inst0_MEM_output_width_17_num_0;
	wire [0:0] OR_CONFIG_EN_SRAM_0_out;
	wire [0:0] OR_CONFIG_EN_SRAM_1_out;
	wire [0:0] OR_CONFIG_RD_SRAM_out;
	wire [0:0] OR_CONFIG_WR_SRAM_out;
	wire [7:0] OR_config_addr_FEATURE_O;
	wire [31:0] OR_config_data_FEATURE_O;
	wire ZextWrapper_19_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_19_32_inst0$self_O_in;
	wire ZextWrapper_25_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_25_32_inst0$self_O_in;
	wire bit_const_1_None_out;
	wire [31:0] config_reg_0_O;
	wire [31:0] config_reg_1_O;
	wire [31:0] config_reg_10_O;
	wire [31:0] config_reg_11_O;
	wire [31:0] config_reg_12_O;
	wire [31:0] config_reg_13_O;
	wire [31:0] config_reg_14_O;
	wire [31:0] config_reg_15_O;
	wire [31:0] config_reg_16_O;
	wire [31:0] config_reg_17_O;
	wire [31:0] config_reg_18_O;
	wire [31:0] config_reg_19_O;
	wire [31:0] config_reg_2_O;
	wire [31:0] config_reg_20_O;
	wire [31:0] config_reg_21_O;
	wire [31:0] config_reg_22_O;
	wire [31:0] config_reg_23_O;
	wire [31:0] config_reg_24_O;
	wire [31:0] config_reg_25_O;
	wire [31:0] config_reg_26_O;
	wire [31:0] config_reg_27_O;
	wire [31:0] config_reg_28_O;
	wire [31:0] config_reg_29_O;
	wire [31:0] config_reg_3_O;
	wire [31:0] config_reg_30_O;
	wire [31:0] config_reg_31_O;
	wire [31:0] config_reg_32_O;
	wire [31:0] config_reg_33_O;
	wire [31:0] config_reg_34_O;
	wire [31:0] config_reg_35_O;
	wire [31:0] config_reg_36_O;
	wire [31:0] config_reg_37_O;
	wire [31:0] config_reg_38_O;
	wire [31:0] config_reg_39_O;
	wire [31:0] config_reg_4_O;
	wire [18:0] config_reg_40_O;
	wire [31:0] config_reg_41_O;
	wire [31:0] config_reg_42_O;
	wire [31:0] config_reg_43_O;
	wire [31:0] config_reg_44_O;
	wire [31:0] config_reg_45_O;
	wire [24:0] config_reg_46_O;
	wire [31:0] config_reg_5_O;
	wire [31:0] config_reg_6_O;
	wire [31:0] config_reg_7_O;
	wire [31:0] config_reg_8_O;
	wire [31:0] config_reg_9_O;
	wire coreir_wrapInAsyncReset_inst0_out;
	wire coreir_wrapOutAsyncReset_inst0_out;
	wire [0:0] flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] flush_mux_sel_value_O;
	wire [0:0] flush_reg_sel_value_O;
	wire [0:0] flush_reg_value_value_O;
	wire [0:0] flush_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] mode_excl_value_O;
	wire [1:0] mode_value_O;
	wire [31:0] mux_aoi_47_32_inst0_O;
	wire [63:0] mux_aoi_47_32_inst0_out_sel;
	wire [7:0] self_config_config_addr_out;
	wire [0:0] tile_en_value_O;
	coreir_and #(.width(1)) AND_CONFIG_EN_SRAM_0(
		.in0(OR_CONFIG_EN_SRAM_0_out),
		.in1(config_en_0),
		.out(AND_CONFIG_EN_SRAM_0_out)
	);
	coreir_and #(.width(1)) AND_CONFIG_EN_SRAM_1(
		.in0(OR_CONFIG_EN_SRAM_1_out),
		.in1(config_en_1),
		.out(AND_CONFIG_EN_SRAM_1_out)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_0_value(
		.I(config_reg_0_O),
		.O(CONFIG_SPACE_0_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_10_value(
		.I(config_reg_2_O),
		.O(CONFIG_SPACE_10_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_11_value(
		.I(config_reg_3_O),
		.O(CONFIG_SPACE_11_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_12_value(
		.I(config_reg_4_O),
		.O(CONFIG_SPACE_12_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_13_value(
		.I(config_reg_5_O),
		.O(CONFIG_SPACE_13_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_14_value(
		.I(config_reg_6_O),
		.O(CONFIG_SPACE_14_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_15_value(
		.I(config_reg_7_O),
		.O(CONFIG_SPACE_15_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_16_value(
		.I(config_reg_8_O),
		.O(CONFIG_SPACE_16_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_17_value(
		.I(config_reg_9_O),
		.O(CONFIG_SPACE_17_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_18_value(
		.I(config_reg_10_O),
		.O(CONFIG_SPACE_18_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_19_value(
		.I(config_reg_11_O),
		.O(CONFIG_SPACE_19_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_1_value(
		.I(config_reg_1_O),
		.O(CONFIG_SPACE_1_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_20_value(
		.I(config_reg_13_O),
		.O(CONFIG_SPACE_20_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_21_value(
		.I(config_reg_14_O),
		.O(CONFIG_SPACE_21_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_22_value(
		.I(config_reg_15_O),
		.O(CONFIG_SPACE_22_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_23_value(
		.I(config_reg_16_O),
		.O(CONFIG_SPACE_23_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_24_value(
		.I(config_reg_17_O),
		.O(CONFIG_SPACE_24_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_25_value(
		.I(config_reg_18_O),
		.O(CONFIG_SPACE_25_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_26_value(
		.I(config_reg_19_O),
		.O(CONFIG_SPACE_26_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_27_value(
		.I(config_reg_20_O),
		.O(CONFIG_SPACE_27_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_28_value(
		.I(config_reg_21_O),
		.O(CONFIG_SPACE_28_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_29_value(
		.I(config_reg_22_O),
		.O(CONFIG_SPACE_29_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_2_value(
		.I(config_reg_12_O),
		.O(CONFIG_SPACE_2_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_30_value(
		.I(config_reg_24_O),
		.O(CONFIG_SPACE_30_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_31_value(
		.I(config_reg_25_O),
		.O(CONFIG_SPACE_31_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_32_value(
		.I(config_reg_26_O),
		.O(CONFIG_SPACE_32_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_33_value(
		.I(config_reg_27_O),
		.O(CONFIG_SPACE_33_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_34_value(
		.I(config_reg_28_O),
		.O(CONFIG_SPACE_34_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_35_value(
		.I(config_reg_29_O),
		.O(CONFIG_SPACE_35_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_36_value(
		.I(config_reg_30_O),
		.O(CONFIG_SPACE_36_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_37_value(
		.I(config_reg_31_O),
		.O(CONFIG_SPACE_37_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_38_value(
		.I(config_reg_32_O),
		.O(CONFIG_SPACE_38_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_39_value(
		.I(config_reg_33_O),
		.O(CONFIG_SPACE_39_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_3_value(
		.I(config_reg_23_O),
		.O(CONFIG_SPACE_3_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_40_value(
		.I(config_reg_35_O),
		.O(CONFIG_SPACE_40_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_41_value(
		.I(config_reg_36_O),
		.O(CONFIG_SPACE_41_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_42_value(
		.I(config_reg_37_O),
		.O(CONFIG_SPACE_42_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_43_value(
		.I(config_reg_38_O),
		.O(CONFIG_SPACE_43_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_44_value(
		.I(config_reg_39_O),
		.O(CONFIG_SPACE_44_value_O)
	);
	SliceWrapper_19_0_19 CONFIG_SPACE_45_value(
		.I(config_reg_40_O),
		.O(CONFIG_SPACE_45_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_4_value(
		.I(config_reg_34_O),
		.O(CONFIG_SPACE_4_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_5_value(
		.I(config_reg_41_O),
		.O(CONFIG_SPACE_5_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_6_value(
		.I(config_reg_42_O),
		.O(CONFIG_SPACE_6_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_7_value(
		.I(config_reg_43_O),
		.O(CONFIG_SPACE_7_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_8_value(
		.I(config_reg_44_O),
		.O(CONFIG_SPACE_8_value_O)
	);
	SliceWrapper_32_0_32 CONFIG_SPACE_9_value(
		.I(config_reg_45_O),
		.O(CONFIG_SPACE_9_value_O)
	);
	coreir_not #(.width(1)) Invert1_inst0(
		.in(coreir_wrapInAsyncReset_inst0_out),
		.out(Invert1_inst0_out)
	);
	coreir_not #(.width(1)) Invert1_inst1(
		.in(stall),
		.out(Invert1_inst1_out)
	);
	SliceWrapper_25_0_1 MEM_input_width_17_num_0_valid_reg_sel_value(
		.I(config_reg_46_O),
		.O(MEM_input_width_17_num_0_valid_reg_sel_value_O)
	);
	SliceWrapper_25_1_2 MEM_input_width_17_num_0_valid_reg_value_value(
		.I(config_reg_46_O),
		.O(MEM_input_width_17_num_0_valid_reg_value_value_O)
	);
	coreir_mux #(.width(1)) MEM_input_width_17_num_0_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MEM_input_width_17_num_0_valid),
		.in1(MEM_input_width_17_num_0_valid_reg_value_value_O),
		.sel(MEM_input_width_17_num_0_valid_reg_sel_value_O[0]),
		.out(MEM_input_width_17_num_0_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_25_2_3 MEM_input_width_17_num_1_valid_reg_sel_value(
		.I(config_reg_46_O),
		.O(MEM_input_width_17_num_1_valid_reg_sel_value_O)
	);
	SliceWrapper_25_3_4 MEM_input_width_17_num_1_valid_reg_value_value(
		.I(config_reg_46_O),
		.O(MEM_input_width_17_num_1_valid_reg_value_value_O)
	);
	coreir_mux #(.width(1)) MEM_input_width_17_num_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MEM_input_width_17_num_1_valid),
		.in1(MEM_input_width_17_num_1_valid_reg_value_value_O),
		.sel(MEM_input_width_17_num_1_valid_reg_sel_value_O[0]),
		.out(MEM_input_width_17_num_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_25_4_5 MEM_input_width_17_num_2_valid_reg_sel_value(
		.I(config_reg_46_O),
		.O(MEM_input_width_17_num_2_valid_reg_sel_value_O)
	);
	SliceWrapper_25_5_6 MEM_input_width_17_num_2_valid_reg_value_value(
		.I(config_reg_46_O),
		.O(MEM_input_width_17_num_2_valid_reg_value_value_O)
	);
	coreir_mux #(.width(1)) MEM_input_width_17_num_2_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MEM_input_width_17_num_2_valid),
		.in1(MEM_input_width_17_num_2_valid_reg_value_value_O),
		.sel(MEM_input_width_17_num_2_valid_reg_sel_value_O[0]),
		.out(MEM_input_width_17_num_2_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_25_6_7 MEM_input_width_17_num_3_valid_reg_sel_value(
		.I(config_reg_46_O),
		.O(MEM_input_width_17_num_3_valid_reg_sel_value_O)
	);
	SliceWrapper_25_7_8 MEM_input_width_17_num_3_valid_reg_value_value(
		.I(config_reg_46_O),
		.O(MEM_input_width_17_num_3_valid_reg_value_value_O)
	);
	coreir_mux #(.width(1)) MEM_input_width_17_num_3_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MEM_input_width_17_num_3_valid),
		.in1(MEM_input_width_17_num_3_valid_reg_value_value_O),
		.sel(MEM_input_width_17_num_3_valid_reg_sel_value_O[0]),
		.out(MEM_input_width_17_num_3_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_25_8_9 MEM_input_width_1_num_0_reg_sel_value(
		.I(config_reg_46_O),
		.O(MEM_input_width_1_num_0_reg_sel_value_O)
	);
	SliceWrapper_25_9_10 MEM_input_width_1_num_0_reg_value_value(
		.I(config_reg_46_O),
		.O(MEM_input_width_1_num_0_reg_value_value_O)
	);
	coreir_mux #(.width(1)) MEM_input_width_1_num_0_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MEM_input_width_1_num_0),
		.in1(MEM_input_width_1_num_0_reg_value_value_O),
		.sel(MEM_input_width_1_num_0_reg_sel_value_O[0]),
		.out(MEM_input_width_1_num_0_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_25_10_11 MEM_input_width_1_num_1_reg_sel_value(
		.I(config_reg_46_O),
		.O(MEM_input_width_1_num_1_reg_sel_value_O)
	);
	SliceWrapper_25_11_12 MEM_input_width_1_num_1_reg_value_value(
		.I(config_reg_46_O),
		.O(MEM_input_width_1_num_1_reg_value_value_O)
	);
	coreir_mux #(.width(1)) MEM_input_width_1_num_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MEM_input_width_1_num_1),
		.in1(MEM_input_width_1_num_1_reg_value_value_O),
		.sel(MEM_input_width_1_num_1_reg_sel_value_O[0]),
		.out(MEM_input_width_1_num_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_25_12_13 MEM_output_width_17_num_0_ready_reg_sel_value(
		.I(config_reg_46_O),
		.O(MEM_output_width_17_num_0_ready_reg_sel_value_O)
	);
	SliceWrapper_25_13_14 MEM_output_width_17_num_0_ready_reg_value_value(
		.I(config_reg_46_O),
		.O(MEM_output_width_17_num_0_ready_reg_value_value_O)
	);
	coreir_mux #(.width(1)) MEM_output_width_17_num_0_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MEM_output_width_17_num_0_ready),
		.in1(MEM_output_width_17_num_0_ready_reg_value_value_O),
		.sel(MEM_output_width_17_num_0_ready_reg_sel_value_O[0]),
		.out(MEM_output_width_17_num_0_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_25_14_15 MEM_output_width_17_num_1_ready_reg_sel_value(
		.I(config_reg_46_O),
		.O(MEM_output_width_17_num_1_ready_reg_sel_value_O)
	);
	SliceWrapper_25_15_16 MEM_output_width_17_num_1_ready_reg_value_value(
		.I(config_reg_46_O),
		.O(MEM_output_width_17_num_1_ready_reg_value_value_O)
	);
	coreir_mux #(.width(1)) MEM_output_width_17_num_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MEM_output_width_17_num_1_ready),
		.in1(MEM_output_width_17_num_1_ready_reg_value_value_O),
		.sel(MEM_output_width_17_num_1_ready_reg_sel_value_O[0]),
		.out(MEM_output_width_17_num_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_25_16_17 MEM_output_width_17_num_2_ready_reg_sel_value(
		.I(config_reg_46_O),
		.O(MEM_output_width_17_num_2_ready_reg_sel_value_O)
	);
	SliceWrapper_25_17_18 MEM_output_width_17_num_2_ready_reg_value_value(
		.I(config_reg_46_O),
		.O(MEM_output_width_17_num_2_ready_reg_value_value_O)
	);
	coreir_mux #(.width(1)) MEM_output_width_17_num_2_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MEM_output_width_17_num_2_ready),
		.in1(MEM_output_width_17_num_2_ready_reg_value_value_O),
		.sel(MEM_output_width_17_num_2_ready_reg_sel_value_O[0]),
		.out(MEM_output_width_17_num_2_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	wire [1:0] MemCore_inner_W_inst0_config_en;
	assign MemCore_inner_W_inst0_config_en = {AND_CONFIG_EN_SRAM_1_out[0], AND_CONFIG_EN_SRAM_0_out[0]};
	MemCore_inner_W MemCore_inner_W_inst0(
		.config_data_out_1(MemCore_inner_W_inst0_config_data_out_1),
		.CONFIG_SPACE_24(CONFIG_SPACE_24_value_O),
		.CONFIG_SPACE_38(CONFIG_SPACE_38_value_O),
		.CONFIG_SPACE_11(CONFIG_SPACE_11_value_O),
		.MEM_input_width_17_num_2_valid(MEM_input_width_17_num_2_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.config_data_in(OR_config_data_FEATURE_O),
		.CONFIG_SPACE_0(CONFIG_SPACE_0_value_O),
		.CONFIG_SPACE_42(CONFIG_SPACE_42_value_O),
		.CONFIG_SPACE_43(CONFIG_SPACE_43_value_O),
		.CONFIG_SPACE_8(CONFIG_SPACE_8_value_O),
		.config_data_out_0(MemCore_inner_W_inst0_config_data_out_0),
		.MEM_input_width_17_num_3_valid(MEM_input_width_17_num_3_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.CONFIG_SPACE_6(CONFIG_SPACE_6_value_O),
		.CONFIG_SPACE_13(CONFIG_SPACE_13_value_O),
		.CONFIG_SPACE_3(CONFIG_SPACE_3_value_O),
		.CONFIG_SPACE_30(CONFIG_SPACE_30_value_O),
		.CONFIG_SPACE_29(CONFIG_SPACE_29_value_O),
		.CONFIG_SPACE_1(CONFIG_SPACE_1_value_O),
		.CONFIG_SPACE_33(CONFIG_SPACE_33_value_O),
		.CONFIG_SPACE_44(CONFIG_SPACE_44_value_O),
		.MEM_input_width_17_num_0(MEM_input_width_17_num_0),
		.MEM_input_width_17_num_2(MEM_input_width_17_num_2),
		.CONFIG_SPACE_20(CONFIG_SPACE_20_value_O),
		.MEM_output_width_17_num_2_ready(MEM_output_width_17_num_2_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.MEM_input_width_17_num_3_ready(MemCore_inner_W_inst0_MEM_input_width_17_num_3_ready),
		.CONFIG_SPACE_37(CONFIG_SPACE_37_value_O),
		.tile_en(tile_en_value_O),
		.MEM_output_width_1_num_2(MemCore_inner_W_inst0_MEM_output_width_1_num_2),
		.MEM_output_width_1_num_1(MemCore_inner_W_inst0_MEM_output_width_1_num_1),
		.CONFIG_SPACE_9(CONFIG_SPACE_9_value_O),
		.clk(clk),
		.CONFIG_SPACE_35(CONFIG_SPACE_35_value_O),
		.CONFIG_SPACE_40(CONFIG_SPACE_40_value_O),
		.MEM_output_width_17_num_1_ready(MEM_output_width_17_num_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.CONFIG_SPACE_36(CONFIG_SPACE_36_value_O),
		.CONFIG_SPACE_2(CONFIG_SPACE_2_value_O),
		.CONFIG_SPACE_28(CONFIG_SPACE_28_value_O),
		.MEM_output_width_17_num_1_valid(MemCore_inner_W_inst0_MEM_output_width_17_num_1_valid),
		.MEM_output_width_17_num_2(MemCore_inner_W_inst0_MEM_output_width_17_num_2),
		.rst_n(coreir_wrapOutAsyncReset_inst0_out),
		.MEM_input_width_17_num_0_valid(MEM_input_width_17_num_0_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.MEM_input_width_17_num_2_ready(MemCore_inner_W_inst0_MEM_input_width_17_num_2_ready),
		.MEM_output_width_17_num_1(MemCore_inner_W_inst0_MEM_output_width_17_num_1),
		.MEM_output_width_1_num_0(MemCore_inner_W_inst0_MEM_output_width_1_num_0),
		.CONFIG_SPACE_34(CONFIG_SPACE_34_value_O),
		.CONFIG_SPACE_39(CONFIG_SPACE_39_value_O),
		.clk_en(Invert1_inst1_out),
		.CONFIG_SPACE_14(CONFIG_SPACE_14_value_O),
		.CONFIG_SPACE_32(CONFIG_SPACE_32_value_O),
		.MEM_output_width_17_num_2_valid(MemCore_inner_W_inst0_MEM_output_width_17_num_2_valid),
		.CONFIG_SPACE_31(CONFIG_SPACE_31_value_O),
		.MEM_input_width_1_num_1(MEM_input_width_1_num_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.CONFIG_SPACE_41(CONFIG_SPACE_41_value_O),
		.MEM_output_width_17_num_0_ready(MEM_output_width_17_num_0_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.MEM_input_width_17_num_1(MEM_input_width_17_num_1),
		.mode(mode_value_O),
		.MEM_input_width_1_num_0(MEM_input_width_1_num_0_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.CONFIG_SPACE_19(CONFIG_SPACE_19_value_O),
		.CONFIG_SPACE_22(CONFIG_SPACE_22_value_O),
		.CONFIG_SPACE_16(CONFIG_SPACE_16_value_O),
		.MEM_input_width_17_num_1_ready(MemCore_inner_W_inst0_MEM_input_width_17_num_1_ready),
		.CONFIG_SPACE_12(CONFIG_SPACE_12_value_O),
		.config_addr_in(OR_config_addr_FEATURE_O),
		.CONFIG_SPACE_7(CONFIG_SPACE_7_value_O),
		.CONFIG_SPACE_27(CONFIG_SPACE_27_value_O),
		.MEM_input_width_17_num_0_ready(MemCore_inner_W_inst0_MEM_input_width_17_num_0_ready),
		.CONFIG_SPACE_5(CONFIG_SPACE_5_value_O),
		.MEM_input_width_17_num_1_valid(MEM_input_width_17_num_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.CONFIG_SPACE_25(CONFIG_SPACE_25_value_O),
		.config_write(OR_CONFIG_RD_SRAM_out),
		.CONFIG_SPACE_45(CONFIG_SPACE_45_value_O),
		.CONFIG_SPACE_17(CONFIG_SPACE_17_value_O),
		.MEM_input_width_17_num_3(MEM_input_width_17_num_3),
		.config_en(MemCore_inner_W_inst0_config_en),
		.CONFIG_SPACE_23(CONFIG_SPACE_23_value_O),
		.CONFIG_SPACE_18(CONFIG_SPACE_18_value_O),
		.CONFIG_SPACE_10(CONFIG_SPACE_10_value_O),
		.CONFIG_SPACE_21(CONFIG_SPACE_21_value_O),
		.flush(flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.mode_excl(mode_excl_value_O),
		.MEM_output_width_17_num_0_valid(MemCore_inner_W_inst0_MEM_output_width_17_num_0_valid),
		.CONFIG_SPACE_4(CONFIG_SPACE_4_value_O),
		.MEM_output_width_17_num_0(MemCore_inner_W_inst0_MEM_output_width_17_num_0),
		.CONFIG_SPACE_26(CONFIG_SPACE_26_value_O),
		.CONFIG_SPACE_15(CONFIG_SPACE_15_value_O),
		.config_read(OR_CONFIG_WR_SRAM_out)
	);
	coreir_or #(.width(1)) OR_CONFIG_EN_SRAM_0(
		.in0(config_1_write),
		.in1(config_1_read),
		.out(OR_CONFIG_EN_SRAM_0_out)
	);
	coreir_or #(.width(1)) OR_CONFIG_EN_SRAM_1(
		.in0(config_2_write),
		.in1(config_2_read),
		.out(OR_CONFIG_EN_SRAM_1_out)
	);
	coreir_or #(.width(1)) OR_CONFIG_RD_SRAM(
		.in0(config_1_write),
		.in1(config_2_write),
		.out(OR_CONFIG_RD_SRAM_out)
	);
	coreir_or #(.width(1)) OR_CONFIG_WR_SRAM(
		.in0(config_1_read),
		.in1(config_2_read),
		.out(OR_CONFIG_WR_SRAM_out)
	);
	wire [7:0] OR_config_addr_FEATURE_I0;
	assign OR_config_addr_FEATURE_I0 = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	Or3x8 OR_config_addr_FEATURE(
		.I0(OR_config_addr_FEATURE_I0),
		.I1(config_1_config_addr),
		.I2(config_2_config_addr),
		.O(OR_config_addr_FEATURE_O)
	);
	Or3x32 OR_config_data_FEATURE(
		.I0(config_config_data),
		.I1(config_1_config_data),
		.I2(config_2_config_data),
		.O(OR_config_data_FEATURE_O)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_19_32_inst0$bit_const_0_None(.out(ZextWrapper_19_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_19_32_inst0$self_O_out;
	assign ZextWrapper_19_32_inst0$self_O_out = {ZextWrapper_19_32_inst0$bit_const_0_None_out, ZextWrapper_19_32_inst0$bit_const_0_None_out, ZextWrapper_19_32_inst0$bit_const_0_None_out, ZextWrapper_19_32_inst0$bit_const_0_None_out, ZextWrapper_19_32_inst0$bit_const_0_None_out, ZextWrapper_19_32_inst0$bit_const_0_None_out, ZextWrapper_19_32_inst0$bit_const_0_None_out, ZextWrapper_19_32_inst0$bit_const_0_None_out, ZextWrapper_19_32_inst0$bit_const_0_None_out, ZextWrapper_19_32_inst0$bit_const_0_None_out, ZextWrapper_19_32_inst0$bit_const_0_None_out, ZextWrapper_19_32_inst0$bit_const_0_None_out, ZextWrapper_19_32_inst0$bit_const_0_None_out, config_reg_40_O};
	mantle_wire__typeBitIn32 ZextWrapper_19_32_inst0$self_O(
		.in(ZextWrapper_19_32_inst0$self_O_in),
		.out(ZextWrapper_19_32_inst0$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_25_32_inst0$bit_const_0_None(.out(ZextWrapper_25_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_25_32_inst0$self_O_out;
	assign ZextWrapper_25_32_inst0$self_O_out = {ZextWrapper_25_32_inst0$bit_const_0_None_out, ZextWrapper_25_32_inst0$bit_const_0_None_out, ZextWrapper_25_32_inst0$bit_const_0_None_out, ZextWrapper_25_32_inst0$bit_const_0_None_out, ZextWrapper_25_32_inst0$bit_const_0_None_out, ZextWrapper_25_32_inst0$bit_const_0_None_out, ZextWrapper_25_32_inst0$bit_const_0_None_out, config_reg_46_O};
	mantle_wire__typeBitIn32 ZextWrapper_25_32_inst0$self_O(
		.in(ZextWrapper_25_32_inst0$self_O_in),
		.out(ZextWrapper_25_32_inst0$self_O_out)
	);
	corebit_const #(.value(1'b1)) bit_const_1_None(.out(bit_const_1_None_out));
	wire [7:0] config_reg_0_config_addr;
	assign config_reg_0_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_reg_0_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_1_config_addr;
	assign config_reg_1_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_1 config_reg_1(
		.clk(clk),
		.reset(reset),
		.O(config_reg_1_O),
		.config_addr(config_reg_1_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_10_config_addr;
	assign config_reg_10_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_10 config_reg_10(
		.clk(clk),
		.reset(reset),
		.O(config_reg_10_O),
		.config_addr(config_reg_10_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_11_config_addr;
	assign config_reg_11_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_11 config_reg_11(
		.clk(clk),
		.reset(reset),
		.O(config_reg_11_O),
		.config_addr(config_reg_11_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_12_config_addr;
	assign config_reg_12_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_12 config_reg_12(
		.clk(clk),
		.reset(reset),
		.O(config_reg_12_O),
		.config_addr(config_reg_12_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_13_config_addr;
	assign config_reg_13_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_13 config_reg_13(
		.clk(clk),
		.reset(reset),
		.O(config_reg_13_O),
		.config_addr(config_reg_13_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_14_config_addr;
	assign config_reg_14_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_14 config_reg_14(
		.clk(clk),
		.reset(reset),
		.O(config_reg_14_O),
		.config_addr(config_reg_14_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_15_config_addr;
	assign config_reg_15_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_15 config_reg_15(
		.clk(clk),
		.reset(reset),
		.O(config_reg_15_O),
		.config_addr(config_reg_15_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_16_config_addr;
	assign config_reg_16_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_16 config_reg_16(
		.clk(clk),
		.reset(reset),
		.O(config_reg_16_O),
		.config_addr(config_reg_16_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_17_config_addr;
	assign config_reg_17_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_17 config_reg_17(
		.clk(clk),
		.reset(reset),
		.O(config_reg_17_O),
		.config_addr(config_reg_17_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_18_config_addr;
	assign config_reg_18_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_18 config_reg_18(
		.clk(clk),
		.reset(reset),
		.O(config_reg_18_O),
		.config_addr(config_reg_18_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_19_config_addr;
	assign config_reg_19_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_19 config_reg_19(
		.clk(clk),
		.reset(reset),
		.O(config_reg_19_O),
		.config_addr(config_reg_19_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_2_config_addr;
	assign config_reg_2_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_2 config_reg_2(
		.clk(clk),
		.reset(reset),
		.O(config_reg_2_O),
		.config_addr(config_reg_2_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_20_config_addr;
	assign config_reg_20_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_20 config_reg_20(
		.clk(clk),
		.reset(reset),
		.O(config_reg_20_O),
		.config_addr(config_reg_20_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_21_config_addr;
	assign config_reg_21_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_21 config_reg_21(
		.clk(clk),
		.reset(reset),
		.O(config_reg_21_O),
		.config_addr(config_reg_21_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_22_config_addr;
	assign config_reg_22_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_22 config_reg_22(
		.clk(clk),
		.reset(reset),
		.O(config_reg_22_O),
		.config_addr(config_reg_22_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_23_config_addr;
	assign config_reg_23_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_23 config_reg_23(
		.clk(clk),
		.reset(reset),
		.O(config_reg_23_O),
		.config_addr(config_reg_23_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_24_config_addr;
	assign config_reg_24_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_24 config_reg_24(
		.clk(clk),
		.reset(reset),
		.O(config_reg_24_O),
		.config_addr(config_reg_24_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_25_config_addr;
	assign config_reg_25_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_25 config_reg_25(
		.clk(clk),
		.reset(reset),
		.O(config_reg_25_O),
		.config_addr(config_reg_25_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_26_config_addr;
	assign config_reg_26_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_26 config_reg_26(
		.clk(clk),
		.reset(reset),
		.O(config_reg_26_O),
		.config_addr(config_reg_26_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_27_config_addr;
	assign config_reg_27_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_27 config_reg_27(
		.clk(clk),
		.reset(reset),
		.O(config_reg_27_O),
		.config_addr(config_reg_27_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_28_config_addr;
	assign config_reg_28_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_28 config_reg_28(
		.clk(clk),
		.reset(reset),
		.O(config_reg_28_O),
		.config_addr(config_reg_28_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_29_config_addr;
	assign config_reg_29_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_29 config_reg_29(
		.clk(clk),
		.reset(reset),
		.O(config_reg_29_O),
		.config_addr(config_reg_29_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_3_config_addr;
	assign config_reg_3_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_3 config_reg_3(
		.clk(clk),
		.reset(reset),
		.O(config_reg_3_O),
		.config_addr(config_reg_3_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_30_config_addr;
	assign config_reg_30_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_30 config_reg_30(
		.clk(clk),
		.reset(reset),
		.O(config_reg_30_O),
		.config_addr(config_reg_30_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_31_config_addr;
	assign config_reg_31_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_31 config_reg_31(
		.clk(clk),
		.reset(reset),
		.O(config_reg_31_O),
		.config_addr(config_reg_31_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_32_config_addr;
	assign config_reg_32_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_32 config_reg_32(
		.clk(clk),
		.reset(reset),
		.O(config_reg_32_O),
		.config_addr(config_reg_32_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_33_config_addr;
	assign config_reg_33_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_33 config_reg_33(
		.clk(clk),
		.reset(reset),
		.O(config_reg_33_O),
		.config_addr(config_reg_33_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_34_config_addr;
	assign config_reg_34_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_34 config_reg_34(
		.clk(clk),
		.reset(reset),
		.O(config_reg_34_O),
		.config_addr(config_reg_34_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_35_config_addr;
	assign config_reg_35_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_35 config_reg_35(
		.clk(clk),
		.reset(reset),
		.O(config_reg_35_O),
		.config_addr(config_reg_35_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_36_config_addr;
	assign config_reg_36_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_36 config_reg_36(
		.clk(clk),
		.reset(reset),
		.O(config_reg_36_O),
		.config_addr(config_reg_36_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_37_config_addr;
	assign config_reg_37_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_37 config_reg_37(
		.clk(clk),
		.reset(reset),
		.O(config_reg_37_O),
		.config_addr(config_reg_37_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_38_config_addr;
	assign config_reg_38_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_38 config_reg_38(
		.clk(clk),
		.reset(reset),
		.O(config_reg_38_O),
		.config_addr(config_reg_38_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_39_config_addr;
	assign config_reg_39_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_39 config_reg_39(
		.clk(clk),
		.reset(reset),
		.O(config_reg_39_O),
		.config_addr(config_reg_39_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_4_config_addr;
	assign config_reg_4_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_4 config_reg_4(
		.clk(clk),
		.reset(reset),
		.O(config_reg_4_O),
		.config_addr(config_reg_4_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_40_config_addr;
	assign config_reg_40_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_19_8_32_40 config_reg_40(
		.clk(clk),
		.reset(reset),
		.O(config_reg_40_O),
		.config_addr(config_reg_40_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_41_config_addr;
	assign config_reg_41_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_41 config_reg_41(
		.clk(clk),
		.reset(reset),
		.O(config_reg_41_O),
		.config_addr(config_reg_41_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_42_config_addr;
	assign config_reg_42_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_42 config_reg_42(
		.clk(clk),
		.reset(reset),
		.O(config_reg_42_O),
		.config_addr(config_reg_42_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_43_config_addr;
	assign config_reg_43_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_43 config_reg_43(
		.clk(clk),
		.reset(reset),
		.O(config_reg_43_O),
		.config_addr(config_reg_43_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_44_config_addr;
	assign config_reg_44_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_44 config_reg_44(
		.clk(clk),
		.reset(reset),
		.O(config_reg_44_O),
		.config_addr(config_reg_44_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_45_config_addr;
	assign config_reg_45_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_45 config_reg_45(
		.clk(clk),
		.reset(reset),
		.O(config_reg_45_O),
		.config_addr(config_reg_45_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_46_config_addr;
	assign config_reg_46_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_25_8_32_46 config_reg_46(
		.clk(clk),
		.reset(reset),
		.O(config_reg_46_O),
		.config_addr(config_reg_46_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_5_config_addr;
	assign config_reg_5_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_5 config_reg_5(
		.clk(clk),
		.reset(reset),
		.O(config_reg_5_O),
		.config_addr(config_reg_5_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_6_config_addr;
	assign config_reg_6_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_6 config_reg_6(
		.clk(clk),
		.reset(reset),
		.O(config_reg_6_O),
		.config_addr(config_reg_6_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_7_config_addr;
	assign config_reg_7_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_7 config_reg_7(
		.clk(clk),
		.reset(reset),
		.O(config_reg_7_O),
		.config_addr(config_reg_7_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_8_config_addr;
	assign config_reg_8_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_8 config_reg_8(
		.clk(clk),
		.reset(reset),
		.O(config_reg_8_O),
		.config_addr(config_reg_8_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	wire [7:0] config_reg_9_config_addr;
	assign config_reg_9_config_addr = {self_config_config_addr_out[7], self_config_config_addr_out[6], self_config_config_addr_out[5:0]};
	ConfigRegister_32_8_32_9 config_reg_9(
		.clk(clk),
		.reset(reset),
		.O(config_reg_9_O),
		.config_addr(config_reg_9_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	coreir_wrap coreir_wrapInAsyncReset_inst0(
		.in(reset),
		.out(coreir_wrapInAsyncReset_inst0_out)
	);
	coreir_wrap coreir_wrapOutAsyncReset_inst0(
		.in(Invert1_inst0_out[0]),
		.out(coreir_wrapOutAsyncReset_inst0_out)
	);
	coreir_mux #(.width(1)) flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(flush_core),
		.in1(flush),
		.sel(flush_mux_sel_value_O[0]),
		.out(flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_25_18_19 flush_mux_sel_value(
		.I(config_reg_46_O),
		.O(flush_mux_sel_value_O)
	);
	SliceWrapper_25_19_20 flush_reg_sel_value(
		.I(config_reg_46_O),
		.O(flush_reg_sel_value_O)
	);
	SliceWrapper_25_20_21 flush_reg_value_value(
		.I(config_reg_46_O),
		.O(flush_reg_value_value_O)
	);
	coreir_mux #(.width(1)) flush_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(flush),
		.in1(flush_reg_value_value_O),
		.sel(flush_reg_sel_value_O[0]),
		.out(flush_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	SliceWrapper_25_23_24 mode_excl_value(
		.I(config_reg_46_O),
		.O(mode_excl_value_O)
	);
	SliceWrapper_25_21_23 mode_value(
		.I(config_reg_46_O),
		.O(mode_value_O)
	);
	wire [1503:0] mux_aoi_47_32_inst0_I;
	assign mux_aoi_47_32_inst0_I[1472+:32] = ZextWrapper_25_32_inst0$self_O_in;
	assign mux_aoi_47_32_inst0_I[1440+:32] = config_reg_45_O;
	assign mux_aoi_47_32_inst0_I[1408+:32] = config_reg_44_O;
	assign mux_aoi_47_32_inst0_I[1376+:32] = config_reg_43_O;
	assign mux_aoi_47_32_inst0_I[1344+:32] = config_reg_42_O;
	assign mux_aoi_47_32_inst0_I[1312+:32] = config_reg_41_O;
	assign mux_aoi_47_32_inst0_I[1280+:32] = ZextWrapper_19_32_inst0$self_O_in;
	assign mux_aoi_47_32_inst0_I[1248+:32] = config_reg_39_O;
	assign mux_aoi_47_32_inst0_I[1216+:32] = config_reg_38_O;
	assign mux_aoi_47_32_inst0_I[1184+:32] = config_reg_37_O;
	assign mux_aoi_47_32_inst0_I[1152+:32] = config_reg_36_O;
	assign mux_aoi_47_32_inst0_I[1120+:32] = config_reg_35_O;
	assign mux_aoi_47_32_inst0_I[1088+:32] = config_reg_34_O;
	assign mux_aoi_47_32_inst0_I[1056+:32] = config_reg_33_O;
	assign mux_aoi_47_32_inst0_I[1024+:32] = config_reg_32_O;
	assign mux_aoi_47_32_inst0_I[992+:32] = config_reg_31_O;
	assign mux_aoi_47_32_inst0_I[960+:32] = config_reg_30_O;
	assign mux_aoi_47_32_inst0_I[928+:32] = config_reg_29_O;
	assign mux_aoi_47_32_inst0_I[896+:32] = config_reg_28_O;
	assign mux_aoi_47_32_inst0_I[864+:32] = config_reg_27_O;
	assign mux_aoi_47_32_inst0_I[832+:32] = config_reg_26_O;
	assign mux_aoi_47_32_inst0_I[800+:32] = config_reg_25_O;
	assign mux_aoi_47_32_inst0_I[768+:32] = config_reg_24_O;
	assign mux_aoi_47_32_inst0_I[736+:32] = config_reg_23_O;
	assign mux_aoi_47_32_inst0_I[704+:32] = config_reg_22_O;
	assign mux_aoi_47_32_inst0_I[672+:32] = config_reg_21_O;
	assign mux_aoi_47_32_inst0_I[640+:32] = config_reg_20_O;
	assign mux_aoi_47_32_inst0_I[608+:32] = config_reg_19_O;
	assign mux_aoi_47_32_inst0_I[576+:32] = config_reg_18_O;
	assign mux_aoi_47_32_inst0_I[544+:32] = config_reg_17_O;
	assign mux_aoi_47_32_inst0_I[512+:32] = config_reg_16_O;
	assign mux_aoi_47_32_inst0_I[480+:32] = config_reg_15_O;
	assign mux_aoi_47_32_inst0_I[448+:32] = config_reg_14_O;
	assign mux_aoi_47_32_inst0_I[416+:32] = config_reg_13_O;
	assign mux_aoi_47_32_inst0_I[384+:32] = config_reg_12_O;
	assign mux_aoi_47_32_inst0_I[352+:32] = config_reg_11_O;
	assign mux_aoi_47_32_inst0_I[320+:32] = config_reg_10_O;
	assign mux_aoi_47_32_inst0_I[288+:32] = config_reg_9_O;
	assign mux_aoi_47_32_inst0_I[256+:32] = config_reg_8_O;
	assign mux_aoi_47_32_inst0_I[224+:32] = config_reg_7_O;
	assign mux_aoi_47_32_inst0_I[192+:32] = config_reg_6_O;
	assign mux_aoi_47_32_inst0_I[160+:32] = config_reg_5_O;
	assign mux_aoi_47_32_inst0_I[128+:32] = config_reg_4_O;
	assign mux_aoi_47_32_inst0_I[96+:32] = config_reg_3_O;
	assign mux_aoi_47_32_inst0_I[64+:32] = config_reg_2_O;
	assign mux_aoi_47_32_inst0_I[32+:32] = config_reg_1_O;
	assign mux_aoi_47_32_inst0_I[0+:32] = config_reg_0_O;
	mux_aoi_47_32 mux_aoi_47_32_inst0(
		.I(mux_aoi_47_32_inst0_I),
		.O(mux_aoi_47_32_inst0_O),
		.S(self_config_config_addr_out[5:0]),
		.out_sel(mux_aoi_47_32_inst0_out_sel)
	);
	mantle_wire__typeBit8 self_config_config_addr(
		.in(config_config_addr),
		.out(self_config_config_addr_out)
	);
	SliceWrapper_25_24_25 tile_en_value(
		.I(config_reg_46_O),
		.O(tile_en_value_O)
	);
	assign MEM_input_width_17_num_0_ready = MemCore_inner_W_inst0_MEM_input_width_17_num_0_ready;
	assign MEM_input_width_17_num_1_ready = MemCore_inner_W_inst0_MEM_input_width_17_num_1_ready;
	assign MEM_input_width_17_num_2_ready = MemCore_inner_W_inst0_MEM_input_width_17_num_2_ready;
	assign MEM_input_width_17_num_3_ready = MemCore_inner_W_inst0_MEM_input_width_17_num_3_ready;
	assign MEM_input_width_1_num_0_ready = bit_const_1_None_out;
	assign MEM_input_width_1_num_1_ready = bit_const_1_None_out;
	assign MEM_output_width_17_num_0 = MemCore_inner_W_inst0_MEM_output_width_17_num_0;
	assign MEM_output_width_17_num_0_valid = MemCore_inner_W_inst0_MEM_output_width_17_num_0_valid;
	assign MEM_output_width_17_num_1 = MemCore_inner_W_inst0_MEM_output_width_17_num_1;
	assign MEM_output_width_17_num_1_valid = MemCore_inner_W_inst0_MEM_output_width_17_num_1_valid;
	assign MEM_output_width_17_num_2 = MemCore_inner_W_inst0_MEM_output_width_17_num_2;
	assign MEM_output_width_17_num_2_valid = MemCore_inner_W_inst0_MEM_output_width_17_num_2_valid;
	assign MEM_output_width_1_num_0 = MemCore_inner_W_inst0_MEM_output_width_1_num_0;
	assign MEM_output_width_1_num_0_valid = bit_const_1_None_out;
	assign MEM_output_width_1_num_1 = MemCore_inner_W_inst0_MEM_output_width_1_num_1;
	assign MEM_output_width_1_num_1_valid = bit_const_1_None_out;
	assign MEM_output_width_1_num_2 = MemCore_inner_W_inst0_MEM_output_width_1_num_2;
	assign MEM_output_width_1_num_2_valid = bit_const_1_None_out;
	assign read_config_data = mux_aoi_47_32_inst0_O;
	assign read_config_data_1 = MemCore_inner_W_inst0_config_data_out_0;
	assign read_config_data_2 = MemCore_inner_W_inst0_config_data_out_1;
endmodule
module CB_flush (
	I,
	O,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	enable,
	out_sel,
	read_config_data,
	ready_in,
	ready_out,
	reset,
	valid_in,
	valid_out
);
	input [19:0] I;
	output wire [0:0] O;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output wire enable;
	output wire [31:0] out_sel;
	output wire [31:0] read_config_data;
	input ready_in;
	output wire ready_out;
	input reset;
	input [19:0] valid_in;
	output wire valid_out;
	wire [0:0] CB_flush_O;
	wire CB_flush_ready_out;
	wire CB_flush_valid_out;
	wire [31:0] CB_flush_out_sel;
	wire [0:0] CB_flush_enable_value_O;
	wire [4:0] CB_flush_sel_value_O;
	wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
	wire [5:0] config_reg_0_O;
	wire [19:0] CB_flush_I;
	assign CB_flush_I[19+:1] = I[19+:1];
	assign CB_flush_I[18+:1] = I[18+:1];
	assign CB_flush_I[17+:1] = I[17+:1];
	assign CB_flush_I[16+:1] = I[16+:1];
	assign CB_flush_I[15+:1] = I[15+:1];
	assign CB_flush_I[14+:1] = I[14+:1];
	assign CB_flush_I[13+:1] = I[13+:1];
	assign CB_flush_I[12+:1] = I[12+:1];
	assign CB_flush_I[11+:1] = I[11+:1];
	assign CB_flush_I[10+:1] = I[10+:1];
	assign CB_flush_I[9+:1] = I[9+:1];
	assign CB_flush_I[8+:1] = I[8+:1];
	assign CB_flush_I[7+:1] = I[7+:1];
	assign CB_flush_I[6+:1] = I[6+:1];
	assign CB_flush_I[5+:1] = I[5+:1];
	assign CB_flush_I[4+:1] = I[4+:1];
	assign CB_flush_I[3+:1] = I[3+:1];
	assign CB_flush_I[2+:1] = I[2+:1];
	assign CB_flush_I[1+:1] = I[1+:1];
	assign CB_flush_I[0+:1] = I[0+:1];
	mux_aoi_ready_valid_const_20_1 CB_flush(
		.I(CB_flush_I),
		.O(CB_flush_O),
		.ready_in(ready_in),
		.ready_out(CB_flush_ready_out),
		.valid_in(valid_in),
		.valid_out(CB_flush_valid_out),
		.S(CB_flush_sel_value_O),
		.out_sel(CB_flush_out_sel)
	);
	SliceWrapper_6_0_1 CB_flush_enable_value(
		.I(config_reg_0_O),
		.O(CB_flush_enable_value_O)
	);
	SliceWrapper_6_1_6 CB_flush_sel_value(
		.I(config_reg_0_O),
		.O(CB_flush_sel_value_O)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_6_32_inst0$bit_const_0_None(.out(ZextWrapper_6_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
	assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, config_reg_0_O};
	mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O(
		.in(ZextWrapper_6_32_inst0$self_O_in),
		.out(ZextWrapper_6_32_inst0$self_O_out)
	);
	ConfigRegister_6_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	assign O = CB_flush_O;
	assign enable = CB_flush_enable_value_O[0];
	assign out_sel = CB_flush_out_sel;
	assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
	assign ready_out = CB_flush_ready_out;
	assign valid_out = CB_flush_valid_out;
endmodule
module CB_f2io_17 (
	O,
	I,
	ready_in,
	ready_out,
	valid_in,
	valid_out,
	out_sel
);
	output wire [16:0] O;
	input [16:0] I;
	input ready_in;
	output wire ready_out;
	input [0:0] valid_in;
	output wire valid_out;
	output wire [0:0] out_sel;
	wire [16:0] CB_f2io_17_O;
	wire CB_f2io_17_ready_out;
	wire CB_f2io_17_valid_out;
	wire [0:0] const_0_1_out;
	MuxWrapperAOI_1_17_ConstReadyValid CB_f2io_17(
		.I(I),
		.O(CB_f2io_17_O),
		.ready_in(ready_in),
		.ready_out(CB_f2io_17_ready_out),
		.valid_in(valid_in[0]),
		.valid_out(CB_f2io_17_valid_out)
	);
	coreir_const #(
		.value(1'h0),
		.width(1)
	) const_0_1(.out(const_0_1_out));
	assign O = CB_f2io_17_O;
	assign ready_out = CB_f2io_17_ready_out;
	assign valid_out = CB_f2io_17_valid_out;
	assign out_sel = const_0_1_out;
endmodule
module CB_f2io_1 (
	O,
	I,
	ready_in,
	ready_out,
	valid_in,
	valid_out,
	out_sel
);
	output wire [0:0] O;
	input [0:0] I;
	input ready_in;
	output wire ready_out;
	input [0:0] valid_in;
	output wire valid_out;
	output wire [0:0] out_sel;
	wire [0:0] CB_f2io_1_O;
	wire CB_f2io_1_ready_out;
	wire CB_f2io_1_valid_out;
	wire [0:0] const_0_1_out;
	MuxWrapperAOI_1_1_ConstReadyValid CB_f2io_1(
		.I(I),
		.O(CB_f2io_1_O),
		.ready_in(ready_in),
		.ready_out(CB_f2io_1_ready_out),
		.valid_in(valid_in[0]),
		.valid_out(CB_f2io_1_valid_out)
	);
	coreir_const #(
		.value(1'h0),
		.width(1)
	) const_0_1(.out(const_0_1_out));
	assign O = CB_f2io_1_O;
	assign ready_out = CB_f2io_1_ready_out;
	assign valid_out = CB_f2io_1_valid_out;
	assign out_sel = const_0_1_out;
endmodule
module Tile_IOCoreReadyValid (
	clk,
	clk_out,
	config_config_addr,
	config_config_data,
	config_out_config_addr,
	config_out_config_data,
	config_out_read,
	config_out_write,
	config_read,
	config_write,
	f2io_1,
	f2io_17,
	f2io_17_ready,
	f2io_17_valid,
	f2io_1_ready,
	f2io_1_valid,
	flush,
	flush_out,
	glb2io_1,
	glb2io_17,
	glb2io_17_ready,
	glb2io_17_valid,
	glb2io_1_ready,
	glb2io_1_valid,
	hi,
	io2f_1,
	io2f_17,
	io2f_17_ready,
	io2f_17_valid,
	io2f_1_ready,
	io2f_1_valid,
	io2glb_1,
	io2glb_17,
	io2glb_17_ready,
	io2glb_17_valid,
	io2glb_1_ready,
	io2glb_1_valid,
	lo,
	read_config_data,
	read_config_data_in,
	reset,
	reset_out,
	stall,
	stall_out,
	tile_id
);
	input clk;
	output wire clk_out;
	input [31:0] config_config_addr;
	input [31:0] config_config_data;
	output wire [31:0] config_out_config_addr;
	output wire [31:0] config_out_config_data;
	output wire [0:0] config_out_read;
	output wire [0:0] config_out_write;
	input [0:0] config_read;
	input [0:0] config_write;
	input [0:0] f2io_1;
	input [16:0] f2io_17;
	output wire f2io_17_ready;
	input f2io_17_valid;
	output wire f2io_1_ready;
	input f2io_1_valid;
	input [0:0] flush;
	output wire [0:0] flush_out;
	input [0:0] glb2io_1;
	input [16:0] glb2io_17;
	output wire glb2io_17_ready;
	input glb2io_17_valid;
	output wire glb2io_1_ready;
	input glb2io_1_valid;
	output wire [8:0] hi;
	output wire [0:0] io2f_1;
	output wire [16:0] io2f_17;
	input [4:0] io2f_17_ready;
	output wire io2f_17_valid;
	input [4:0] io2f_1_ready;
	output wire io2f_1_valid;
	output wire [0:0] io2glb_1;
	output wire [16:0] io2glb_17;
	input io2glb_17_ready;
	output wire io2glb_17_valid;
	input io2glb_1_ready;
	output wire io2glb_1_valid;
	output wire [7:0] lo;
	output wire [31:0] read_config_data;
	input [31:0] read_config_data_in;
	input reset;
	output wire reset_out;
	input [0:0] stall;
	output wire [0:0] stall_out;
	input [15:0] tile_id;
	wire [0:0] CB_f2io_1_O;
	wire CB_f2io_1_ready_out;
	wire CB_f2io_1_valid_out;
	wire [0:0] CB_f2io_1_out_sel;
	wire [16:0] CB_f2io_17_O;
	wire CB_f2io_17_ready_out;
	wire CB_f2io_17_valid_out;
	wire [0:0] CB_f2io_17_out_sel;
	wire DECODE_FEATURE_0_O;
	wire DECODE_FEATURE_1_O;
	wire DECODE_FEATURE_2_O;
	wire DECODE_FEATURE_3_O;
	wire DECODE_FEATURE_4_O;
	wire DECODE_FEATURE_5_O;
	wire FEATURE_AND_0_out;
	wire FEATURE_AND_1_out;
	wire FEATURE_AND_2_out;
	wire FEATURE_AND_3_out;
	wire FEATURE_AND_4_out;
	wire FEATURE_AND_5_out;
	wire [0:0] IOCoreReadyValid_inst0_f2io_17_ready;
	wire [0:0] IOCoreReadyValid_inst0_f2io_1_ready;
	wire [0:0] IOCoreReadyValid_inst0_glb2io_17_ready;
	wire [0:0] IOCoreReadyValid_inst0_glb2io_1_ready;
	wire [0:0] IOCoreReadyValid_inst0_io2f_1;
	wire [16:0] IOCoreReadyValid_inst0_io2f_17;
	wire [0:0] IOCoreReadyValid_inst0_io2f_17_valid;
	wire [0:0] IOCoreReadyValid_inst0_io2f_1_valid;
	wire [0:0] IOCoreReadyValid_inst0_io2glb_1;
	wire [16:0] IOCoreReadyValid_inst0_io2glb_17;
	wire [0:0] IOCoreReadyValid_inst0_io2glb_17_valid;
	wire [0:0] IOCoreReadyValid_inst0_io2glb_1_valid;
	wire [31:0] IOCoreReadyValid_inst0_read_config_data;
	wire [0:0] PowerDomainConfigReg_inst0_ps_en_out;
	wire [31:0] PowerDomainConfigReg_inst0_read_config_data;
	wire [31:0] PowerDomainOR_O;
	wire and_inst0_out;
	wire and_inst1_out;
	wire [31:0] const_0_32_out;
	wire [7:0] const_0_8_out;
	wire [8:0] const_511_9_out;
	wire coreir_eq_16_inst0_out;
	wire io2f_17_ready_merge$andr_inst0_out;
	wire io2f_1_ready_merge$andr_inst0_out;
	wire [31:0] read_data_mux_O;
	wire [31:0] self_config_config_addr_out;
	CB_f2io_1 CB_f2io_1(
		.O(CB_f2io_1_O),
		.I(f2io_1),
		.ready_in(IOCoreReadyValid_inst0_f2io_1_ready[0]),
		.ready_out(CB_f2io_1_ready_out),
		.valid_in(f2io_1_valid),
		.valid_out(CB_f2io_1_valid_out),
		.out_sel(CB_f2io_1_out_sel)
	);
	CB_f2io_17 CB_f2io_17(
		.O(CB_f2io_17_O),
		.I(f2io_17),
		.ready_in(IOCoreReadyValid_inst0_f2io_17_ready[0]),
		.ready_out(CB_f2io_17_ready_out),
		.valid_in(f2io_17_valid),
		.valid_out(CB_f2io_17_valid_out),
		.out_sel(CB_f2io_17_out_sel)
	);
	Decode08 DECODE_FEATURE_0(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_0_O)
	);
	Decode18 DECODE_FEATURE_1(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_1_O)
	);
	Decode28 DECODE_FEATURE_2(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_2_O)
	);
	Decode38 DECODE_FEATURE_3(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_3_O)
	);
	Decode48 DECODE_FEATURE_4(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_4_O)
	);
	Decode58 DECODE_FEATURE_5(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_5_O)
	);
	corebit_and FEATURE_AND_0(
		.in0(DECODE_FEATURE_0_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_0_out)
	);
	corebit_and FEATURE_AND_1(
		.in0(DECODE_FEATURE_1_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_1_out)
	);
	corebit_and FEATURE_AND_2(
		.in0(DECODE_FEATURE_2_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_2_out)
	);
	corebit_and FEATURE_AND_3(
		.in0(DECODE_FEATURE_3_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_3_out)
	);
	corebit_and FEATURE_AND_4(
		.in0(DECODE_FEATURE_4_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_4_out)
	);
	corebit_and FEATURE_AND_5(
		.in0(DECODE_FEATURE_5_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_5_out)
	);
	IOCoreReadyValid IOCoreReadyValid_inst0(
		.clk(clk),
		.config_config_addr(self_config_config_addr_out[31:24]),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_0_out),
		.f2io_1(CB_f2io_1_O),
		.f2io_17(CB_f2io_17_O),
		.f2io_17_ready(IOCoreReadyValid_inst0_f2io_17_ready),
		.f2io_17_valid(CB_f2io_17_valid_out),
		.f2io_1_ready(IOCoreReadyValid_inst0_f2io_1_ready),
		.f2io_1_valid(CB_f2io_1_valid_out),
		.flush(flush),
		.flush_core(flush),
		.glb2io_1(glb2io_1),
		.glb2io_17(glb2io_17),
		.glb2io_17_ready(IOCoreReadyValid_inst0_glb2io_17_ready),
		.glb2io_17_valid(glb2io_17_valid),
		.glb2io_1_ready(IOCoreReadyValid_inst0_glb2io_1_ready),
		.glb2io_1_valid(glb2io_1_valid),
		.io2f_1(IOCoreReadyValid_inst0_io2f_1),
		.io2f_17(IOCoreReadyValid_inst0_io2f_17),
		.io2f_17_ready(io2f_17_ready_merge$andr_inst0_out),
		.io2f_17_valid(IOCoreReadyValid_inst0_io2f_17_valid),
		.io2f_1_ready(io2f_1_ready_merge$andr_inst0_out),
		.io2f_1_valid(IOCoreReadyValid_inst0_io2f_1_valid),
		.io2glb_1(IOCoreReadyValid_inst0_io2glb_1),
		.io2glb_17(IOCoreReadyValid_inst0_io2glb_17),
		.io2glb_17_ready(io2glb_17_ready),
		.io2glb_17_valid(IOCoreReadyValid_inst0_io2glb_17_valid),
		.io2glb_1_ready(io2glb_1_ready),
		.io2glb_1_valid(IOCoreReadyValid_inst0_io2glb_1_valid),
		.read_config_data(IOCoreReadyValid_inst0_read_config_data),
		.reset(reset),
		.stall(stall)
	);
	PowerDomainConfigReg PowerDomainConfigReg_inst0(
		.clk(clk),
		.config_config_addr(self_config_config_addr_out[31:24]),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_5_out),
		.ps_en_out(PowerDomainConfigReg_inst0_ps_en_out),
		.read_config_data(PowerDomainConfigReg_inst0_read_config_data),
		.reset(reset)
	);
	PowerDomainOR PowerDomainOR(
		.I0(read_data_mux_O),
		.I1(read_config_data_in),
		.O(PowerDomainOR_O),
		.I_not(PowerDomainConfigReg_inst0_ps_en_out)
	);
	corebit_and and_inst0(
		.in0(coreir_eq_16_inst0_out),
		.in1(config_read[0]),
		.out(and_inst0_out)
	);
	corebit_and and_inst1(
		.in0(coreir_eq_16_inst0_out),
		.in1(config_write[0]),
		.out(and_inst1_out)
	);
	coreir_const #(
		.value(32'h00000000),
		.width(32)
	) const_0_32(.out(const_0_32_out));
	coreir_const #(
		.value(8'h00),
		.width(8)
	) const_0_8(.out(const_0_8_out));
	coreir_const #(
		.value(9'h1ff),
		.width(9)
	) const_511_9(.out(const_511_9_out));
	coreir_eq #(.width(16)) coreir_eq_16_inst0(
		.in0(tile_id),
		.in1(self_config_config_addr_out[15:0]),
		.out(coreir_eq_16_inst0_out)
	);
	wire [4:0] io2f_17_ready_merge$andr_inst0_in;
	assign io2f_17_ready_merge$andr_inst0_in = {io2f_17_ready[4], io2f_17_ready[3], io2f_17_ready[2], io2f_17_ready[1], io2f_17_ready[0]};
	coreir_andr #(.width(5)) io2f_17_ready_merge$andr_inst0(
		.in(io2f_17_ready_merge$andr_inst0_in),
		.out(io2f_17_ready_merge$andr_inst0_out)
	);
	wire [4:0] io2f_1_ready_merge$andr_inst0_in;
	assign io2f_1_ready_merge$andr_inst0_in = {io2f_1_ready[4], io2f_1_ready[3], io2f_1_ready[2], io2f_1_ready[1], io2f_1_ready[0]};
	coreir_andr #(.width(5)) io2f_1_ready_merge$andr_inst0(
		.in(io2f_1_ready_merge$andr_inst0_in),
		.out(io2f_1_ready_merge$andr_inst0_out)
	);
	wire [191:0] read_data_mux_I;
	assign read_data_mux_I[160+:32] = PowerDomainConfigReg_inst0_read_config_data;
	assign read_data_mux_I[128+:32] = const_0_32_out;
	assign read_data_mux_I[96+:32] = const_0_32_out;
	assign read_data_mux_I[64+:32] = const_0_32_out;
	assign read_data_mux_I[32+:32] = const_0_32_out;
	assign read_data_mux_I[0+:32] = IOCoreReadyValid_inst0_read_config_data;
	MuxWithDefaultWrapper_6_32_8_0 read_data_mux(
		.I(read_data_mux_I),
		.S(self_config_config_addr_out[23:16]),
		.EN(and_inst0_out),
		.O(read_data_mux_O)
	);
	mantle_wire__typeBit32 self_config_config_addr(
		.in(config_config_addr),
		.out(self_config_config_addr_out)
	);
	assign clk_out = clk;
	assign config_out_config_addr = config_config_addr;
	assign config_out_config_data = config_config_data;
	assign config_out_read = config_read;
	assign config_out_write = config_write;
	assign f2io_17_ready = CB_f2io_17_ready_out;
	assign f2io_1_ready = CB_f2io_1_ready_out;
	assign flush_out = flush;
	assign glb2io_17_ready = IOCoreReadyValid_inst0_glb2io_17_ready[0];
	assign glb2io_1_ready = IOCoreReadyValid_inst0_glb2io_1_ready[0];
	assign hi = const_511_9_out;
	assign io2f_1 = IOCoreReadyValid_inst0_io2f_1;
	assign io2f_17 = IOCoreReadyValid_inst0_io2f_17;
	assign io2f_17_valid = IOCoreReadyValid_inst0_io2f_17_valid[0];
	assign io2f_1_valid = IOCoreReadyValid_inst0_io2f_1_valid[0];
	assign io2glb_1 = IOCoreReadyValid_inst0_io2glb_1;
	assign io2glb_17 = IOCoreReadyValid_inst0_io2glb_17;
	assign io2glb_17_valid = IOCoreReadyValid_inst0_io2glb_17_valid[0];
	assign io2glb_1_valid = IOCoreReadyValid_inst0_io2glb_1_valid[0];
	assign lo = const_0_8_out;
	assign read_config_data = PowerDomainOR_O;
	assign reset_out = reset;
	assign stall_out = stall;
endmodule
module CB_PondTop_input_width_17_num_1 (
	I,
	O,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	enable,
	out_sel,
	read_config_data,
	ready_in,
	ready_out,
	reset,
	valid_in,
	valid_out
);
	input [356:0] I;
	output wire [16:0] O;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output wire enable;
	output wire [31:0] out_sel;
	output wire [31:0] read_config_data;
	input ready_in;
	output wire ready_out;
	input reset;
	input [20:0] valid_in;
	output wire valid_out;
	wire [16:0] CB_PondTop_input_width_17_num_1_O;
	wire CB_PondTop_input_width_17_num_1_ready_out;
	wire CB_PondTop_input_width_17_num_1_valid_out;
	wire [31:0] CB_PondTop_input_width_17_num_1_out_sel;
	wire [0:0] CB_PondTop_input_width_17_num_1_enable_value_O;
	wire [4:0] CB_PondTop_input_width_17_num_1_sel_value_O;
	wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
	wire [5:0] config_reg_0_O;
	wire [356:0] CB_PondTop_input_width_17_num_1_I;
	assign CB_PondTop_input_width_17_num_1_I[340+:17] = I[340+:17];
	assign CB_PondTop_input_width_17_num_1_I[323+:17] = I[323+:17];
	assign CB_PondTop_input_width_17_num_1_I[306+:17] = I[306+:17];
	assign CB_PondTop_input_width_17_num_1_I[289+:17] = I[289+:17];
	assign CB_PondTop_input_width_17_num_1_I[272+:17] = I[272+:17];
	assign CB_PondTop_input_width_17_num_1_I[255+:17] = I[255+:17];
	assign CB_PondTop_input_width_17_num_1_I[238+:17] = I[238+:17];
	assign CB_PondTop_input_width_17_num_1_I[221+:17] = I[221+:17];
	assign CB_PondTop_input_width_17_num_1_I[204+:17] = I[204+:17];
	assign CB_PondTop_input_width_17_num_1_I[187+:17] = I[187+:17];
	assign CB_PondTop_input_width_17_num_1_I[170+:17] = I[170+:17];
	assign CB_PondTop_input_width_17_num_1_I[153+:17] = I[153+:17];
	assign CB_PondTop_input_width_17_num_1_I[136+:17] = I[136+:17];
	assign CB_PondTop_input_width_17_num_1_I[119+:17] = I[119+:17];
	assign CB_PondTop_input_width_17_num_1_I[102+:17] = I[102+:17];
	assign CB_PondTop_input_width_17_num_1_I[85+:17] = I[85+:17];
	assign CB_PondTop_input_width_17_num_1_I[68+:17] = I[68+:17];
	assign CB_PondTop_input_width_17_num_1_I[51+:17] = I[51+:17];
	assign CB_PondTop_input_width_17_num_1_I[34+:17] = I[34+:17];
	assign CB_PondTop_input_width_17_num_1_I[17+:17] = I[17+:17];
	assign CB_PondTop_input_width_17_num_1_I[0+:17] = I[0+:17];
	mux_aoi_ready_valid_const_21_17 CB_PondTop_input_width_17_num_1(
		.I(CB_PondTop_input_width_17_num_1_I),
		.O(CB_PondTop_input_width_17_num_1_O),
		.ready_in(ready_in),
		.ready_out(CB_PondTop_input_width_17_num_1_ready_out),
		.valid_in(valid_in),
		.valid_out(CB_PondTop_input_width_17_num_1_valid_out),
		.S(CB_PondTop_input_width_17_num_1_sel_value_O),
		.out_sel(CB_PondTop_input_width_17_num_1_out_sel)
	);
	SliceWrapper_6_0_1 CB_PondTop_input_width_17_num_1_enable_value(
		.I(config_reg_0_O),
		.O(CB_PondTop_input_width_17_num_1_enable_value_O)
	);
	SliceWrapper_6_1_6 CB_PondTop_input_width_17_num_1_sel_value(
		.I(config_reg_0_O),
		.O(CB_PondTop_input_width_17_num_1_sel_value_O)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_6_32_inst0$bit_const_0_None(.out(ZextWrapper_6_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
	assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, config_reg_0_O};
	mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O(
		.in(ZextWrapper_6_32_inst0$self_O_in),
		.out(ZextWrapper_6_32_inst0$self_O_out)
	);
	ConfigRegister_6_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	assign O = CB_PondTop_input_width_17_num_1_O;
	assign enable = CB_PondTop_input_width_17_num_1_enable_value_O[0];
	assign out_sel = CB_PondTop_input_width_17_num_1_out_sel;
	assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
	assign ready_out = CB_PondTop_input_width_17_num_1_ready_out;
	assign valid_out = CB_PondTop_input_width_17_num_1_valid_out;
endmodule
module CB_PondTop_input_width_17_num_0 (
	I,
	O,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	enable,
	out_sel,
	read_config_data,
	ready_in,
	ready_out,
	reset,
	valid_in,
	valid_out
);
	input [356:0] I;
	output wire [16:0] O;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output wire enable;
	output wire [31:0] out_sel;
	output wire [31:0] read_config_data;
	input ready_in;
	output wire ready_out;
	input reset;
	input [20:0] valid_in;
	output wire valid_out;
	wire [16:0] CB_PondTop_input_width_17_num_0_O;
	wire CB_PondTop_input_width_17_num_0_ready_out;
	wire CB_PondTop_input_width_17_num_0_valid_out;
	wire [31:0] CB_PondTop_input_width_17_num_0_out_sel;
	wire [0:0] CB_PondTop_input_width_17_num_0_enable_value_O;
	wire [4:0] CB_PondTop_input_width_17_num_0_sel_value_O;
	wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
	wire [5:0] config_reg_0_O;
	wire [356:0] CB_PondTop_input_width_17_num_0_I;
	assign CB_PondTop_input_width_17_num_0_I[340+:17] = I[340+:17];
	assign CB_PondTop_input_width_17_num_0_I[323+:17] = I[323+:17];
	assign CB_PondTop_input_width_17_num_0_I[306+:17] = I[306+:17];
	assign CB_PondTop_input_width_17_num_0_I[289+:17] = I[289+:17];
	assign CB_PondTop_input_width_17_num_0_I[272+:17] = I[272+:17];
	assign CB_PondTop_input_width_17_num_0_I[255+:17] = I[255+:17];
	assign CB_PondTop_input_width_17_num_0_I[238+:17] = I[238+:17];
	assign CB_PondTop_input_width_17_num_0_I[221+:17] = I[221+:17];
	assign CB_PondTop_input_width_17_num_0_I[204+:17] = I[204+:17];
	assign CB_PondTop_input_width_17_num_0_I[187+:17] = I[187+:17];
	assign CB_PondTop_input_width_17_num_0_I[170+:17] = I[170+:17];
	assign CB_PondTop_input_width_17_num_0_I[153+:17] = I[153+:17];
	assign CB_PondTop_input_width_17_num_0_I[136+:17] = I[136+:17];
	assign CB_PondTop_input_width_17_num_0_I[119+:17] = I[119+:17];
	assign CB_PondTop_input_width_17_num_0_I[102+:17] = I[102+:17];
	assign CB_PondTop_input_width_17_num_0_I[85+:17] = I[85+:17];
	assign CB_PondTop_input_width_17_num_0_I[68+:17] = I[68+:17];
	assign CB_PondTop_input_width_17_num_0_I[51+:17] = I[51+:17];
	assign CB_PondTop_input_width_17_num_0_I[34+:17] = I[34+:17];
	assign CB_PondTop_input_width_17_num_0_I[17+:17] = I[17+:17];
	assign CB_PondTop_input_width_17_num_0_I[0+:17] = I[0+:17];
	mux_aoi_ready_valid_const_21_17 CB_PondTop_input_width_17_num_0(
		.I(CB_PondTop_input_width_17_num_0_I),
		.O(CB_PondTop_input_width_17_num_0_O),
		.ready_in(ready_in),
		.ready_out(CB_PondTop_input_width_17_num_0_ready_out),
		.valid_in(valid_in),
		.valid_out(CB_PondTop_input_width_17_num_0_valid_out),
		.S(CB_PondTop_input_width_17_num_0_sel_value_O),
		.out_sel(CB_PondTop_input_width_17_num_0_out_sel)
	);
	SliceWrapper_6_0_1 CB_PondTop_input_width_17_num_0_enable_value(
		.I(config_reg_0_O),
		.O(CB_PondTop_input_width_17_num_0_enable_value_O)
	);
	SliceWrapper_6_1_6 CB_PondTop_input_width_17_num_0_sel_value(
		.I(config_reg_0_O),
		.O(CB_PondTop_input_width_17_num_0_sel_value_O)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_6_32_inst0$bit_const_0_None(.out(ZextWrapper_6_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
	assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, config_reg_0_O};
	mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O(
		.in(ZextWrapper_6_32_inst0$self_O_in),
		.out(ZextWrapper_6_32_inst0$self_O_out)
	);
	ConfigRegister_6_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	assign O = CB_PondTop_input_width_17_num_0_O;
	assign enable = CB_PondTop_input_width_17_num_0_enable_value_O[0];
	assign out_sel = CB_PondTop_input_width_17_num_0_out_sel;
	assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
	assign ready_out = CB_PondTop_input_width_17_num_0_ready_out;
	assign valid_out = CB_PondTop_input_width_17_num_0_valid_out;
endmodule
module CB_PE_input_width_1_num_2 (
	I,
	O,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	enable,
	out_sel,
	read_config_data,
	ready_in,
	ready_out,
	reset,
	valid_in,
	valid_out
);
	input [19:0] I;
	output wire [0:0] O;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output wire enable;
	output wire [31:0] out_sel;
	output wire [31:0] read_config_data;
	input ready_in;
	output wire ready_out;
	input reset;
	input [19:0] valid_in;
	output wire valid_out;
	wire [0:0] CB_PE_input_width_1_num_2_O;
	wire CB_PE_input_width_1_num_2_ready_out;
	wire CB_PE_input_width_1_num_2_valid_out;
	wire [31:0] CB_PE_input_width_1_num_2_out_sel;
	wire [0:0] CB_PE_input_width_1_num_2_enable_value_O;
	wire [4:0] CB_PE_input_width_1_num_2_sel_value_O;
	wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
	wire [5:0] config_reg_0_O;
	wire [19:0] CB_PE_input_width_1_num_2_I;
	assign CB_PE_input_width_1_num_2_I[19+:1] = I[19+:1];
	assign CB_PE_input_width_1_num_2_I[18+:1] = I[18+:1];
	assign CB_PE_input_width_1_num_2_I[17+:1] = I[17+:1];
	assign CB_PE_input_width_1_num_2_I[16+:1] = I[16+:1];
	assign CB_PE_input_width_1_num_2_I[15+:1] = I[15+:1];
	assign CB_PE_input_width_1_num_2_I[14+:1] = I[14+:1];
	assign CB_PE_input_width_1_num_2_I[13+:1] = I[13+:1];
	assign CB_PE_input_width_1_num_2_I[12+:1] = I[12+:1];
	assign CB_PE_input_width_1_num_2_I[11+:1] = I[11+:1];
	assign CB_PE_input_width_1_num_2_I[10+:1] = I[10+:1];
	assign CB_PE_input_width_1_num_2_I[9+:1] = I[9+:1];
	assign CB_PE_input_width_1_num_2_I[8+:1] = I[8+:1];
	assign CB_PE_input_width_1_num_2_I[7+:1] = I[7+:1];
	assign CB_PE_input_width_1_num_2_I[6+:1] = I[6+:1];
	assign CB_PE_input_width_1_num_2_I[5+:1] = I[5+:1];
	assign CB_PE_input_width_1_num_2_I[4+:1] = I[4+:1];
	assign CB_PE_input_width_1_num_2_I[3+:1] = I[3+:1];
	assign CB_PE_input_width_1_num_2_I[2+:1] = I[2+:1];
	assign CB_PE_input_width_1_num_2_I[1+:1] = I[1+:1];
	assign CB_PE_input_width_1_num_2_I[0+:1] = I[0+:1];
	mux_aoi_ready_valid_const_20_1 CB_PE_input_width_1_num_2(
		.I(CB_PE_input_width_1_num_2_I),
		.O(CB_PE_input_width_1_num_2_O),
		.ready_in(ready_in),
		.ready_out(CB_PE_input_width_1_num_2_ready_out),
		.valid_in(valid_in),
		.valid_out(CB_PE_input_width_1_num_2_valid_out),
		.S(CB_PE_input_width_1_num_2_sel_value_O),
		.out_sel(CB_PE_input_width_1_num_2_out_sel)
	);
	SliceWrapper_6_0_1 CB_PE_input_width_1_num_2_enable_value(
		.I(config_reg_0_O),
		.O(CB_PE_input_width_1_num_2_enable_value_O)
	);
	SliceWrapper_6_1_6 CB_PE_input_width_1_num_2_sel_value(
		.I(config_reg_0_O),
		.O(CB_PE_input_width_1_num_2_sel_value_O)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_6_32_inst0$bit_const_0_None(.out(ZextWrapper_6_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
	assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, config_reg_0_O};
	mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O(
		.in(ZextWrapper_6_32_inst0$self_O_in),
		.out(ZextWrapper_6_32_inst0$self_O_out)
	);
	ConfigRegister_6_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	assign O = CB_PE_input_width_1_num_2_O;
	assign enable = CB_PE_input_width_1_num_2_enable_value_O[0];
	assign out_sel = CB_PE_input_width_1_num_2_out_sel;
	assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
	assign ready_out = CB_PE_input_width_1_num_2_ready_out;
	assign valid_out = CB_PE_input_width_1_num_2_valid_out;
endmodule
module CB_PE_input_width_1_num_1 (
	I,
	O,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	enable,
	out_sel,
	read_config_data,
	ready_in,
	ready_out,
	reset,
	valid_in,
	valid_out
);
	input [19:0] I;
	output wire [0:0] O;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output wire enable;
	output wire [31:0] out_sel;
	output wire [31:0] read_config_data;
	input ready_in;
	output wire ready_out;
	input reset;
	input [19:0] valid_in;
	output wire valid_out;
	wire [0:0] CB_PE_input_width_1_num_1_O;
	wire CB_PE_input_width_1_num_1_ready_out;
	wire CB_PE_input_width_1_num_1_valid_out;
	wire [31:0] CB_PE_input_width_1_num_1_out_sel;
	wire [0:0] CB_PE_input_width_1_num_1_enable_value_O;
	wire [4:0] CB_PE_input_width_1_num_1_sel_value_O;
	wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
	wire [5:0] config_reg_0_O;
	wire [19:0] CB_PE_input_width_1_num_1_I;
	assign CB_PE_input_width_1_num_1_I[19+:1] = I[19+:1];
	assign CB_PE_input_width_1_num_1_I[18+:1] = I[18+:1];
	assign CB_PE_input_width_1_num_1_I[17+:1] = I[17+:1];
	assign CB_PE_input_width_1_num_1_I[16+:1] = I[16+:1];
	assign CB_PE_input_width_1_num_1_I[15+:1] = I[15+:1];
	assign CB_PE_input_width_1_num_1_I[14+:1] = I[14+:1];
	assign CB_PE_input_width_1_num_1_I[13+:1] = I[13+:1];
	assign CB_PE_input_width_1_num_1_I[12+:1] = I[12+:1];
	assign CB_PE_input_width_1_num_1_I[11+:1] = I[11+:1];
	assign CB_PE_input_width_1_num_1_I[10+:1] = I[10+:1];
	assign CB_PE_input_width_1_num_1_I[9+:1] = I[9+:1];
	assign CB_PE_input_width_1_num_1_I[8+:1] = I[8+:1];
	assign CB_PE_input_width_1_num_1_I[7+:1] = I[7+:1];
	assign CB_PE_input_width_1_num_1_I[6+:1] = I[6+:1];
	assign CB_PE_input_width_1_num_1_I[5+:1] = I[5+:1];
	assign CB_PE_input_width_1_num_1_I[4+:1] = I[4+:1];
	assign CB_PE_input_width_1_num_1_I[3+:1] = I[3+:1];
	assign CB_PE_input_width_1_num_1_I[2+:1] = I[2+:1];
	assign CB_PE_input_width_1_num_1_I[1+:1] = I[1+:1];
	assign CB_PE_input_width_1_num_1_I[0+:1] = I[0+:1];
	mux_aoi_ready_valid_const_20_1 CB_PE_input_width_1_num_1(
		.I(CB_PE_input_width_1_num_1_I),
		.O(CB_PE_input_width_1_num_1_O),
		.ready_in(ready_in),
		.ready_out(CB_PE_input_width_1_num_1_ready_out),
		.valid_in(valid_in),
		.valid_out(CB_PE_input_width_1_num_1_valid_out),
		.S(CB_PE_input_width_1_num_1_sel_value_O),
		.out_sel(CB_PE_input_width_1_num_1_out_sel)
	);
	SliceWrapper_6_0_1 CB_PE_input_width_1_num_1_enable_value(
		.I(config_reg_0_O),
		.O(CB_PE_input_width_1_num_1_enable_value_O)
	);
	SliceWrapper_6_1_6 CB_PE_input_width_1_num_1_sel_value(
		.I(config_reg_0_O),
		.O(CB_PE_input_width_1_num_1_sel_value_O)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_6_32_inst0$bit_const_0_None(.out(ZextWrapper_6_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
	assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, config_reg_0_O};
	mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O(
		.in(ZextWrapper_6_32_inst0$self_O_in),
		.out(ZextWrapper_6_32_inst0$self_O_out)
	);
	ConfigRegister_6_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	assign O = CB_PE_input_width_1_num_1_O;
	assign enable = CB_PE_input_width_1_num_1_enable_value_O[0];
	assign out_sel = CB_PE_input_width_1_num_1_out_sel;
	assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
	assign ready_out = CB_PE_input_width_1_num_1_ready_out;
	assign valid_out = CB_PE_input_width_1_num_1_valid_out;
endmodule
module CB_PE_input_width_1_num_0 (
	I,
	O,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	enable,
	out_sel,
	read_config_data,
	ready_in,
	ready_out,
	reset,
	valid_in,
	valid_out
);
	input [20:0] I;
	output wire [0:0] O;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output wire enable;
	output wire [31:0] out_sel;
	output wire [31:0] read_config_data;
	input ready_in;
	output wire ready_out;
	input reset;
	input [20:0] valid_in;
	output wire valid_out;
	wire [0:0] CB_PE_input_width_1_num_0_O;
	wire CB_PE_input_width_1_num_0_ready_out;
	wire CB_PE_input_width_1_num_0_valid_out;
	wire [31:0] CB_PE_input_width_1_num_0_out_sel;
	wire [0:0] CB_PE_input_width_1_num_0_enable_value_O;
	wire [4:0] CB_PE_input_width_1_num_0_sel_value_O;
	wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
	wire [5:0] config_reg_0_O;
	wire [20:0] CB_PE_input_width_1_num_0_I;
	assign CB_PE_input_width_1_num_0_I[20+:1] = I[20+:1];
	assign CB_PE_input_width_1_num_0_I[19+:1] = I[19+:1];
	assign CB_PE_input_width_1_num_0_I[18+:1] = I[18+:1];
	assign CB_PE_input_width_1_num_0_I[17+:1] = I[17+:1];
	assign CB_PE_input_width_1_num_0_I[16+:1] = I[16+:1];
	assign CB_PE_input_width_1_num_0_I[15+:1] = I[15+:1];
	assign CB_PE_input_width_1_num_0_I[14+:1] = I[14+:1];
	assign CB_PE_input_width_1_num_0_I[13+:1] = I[13+:1];
	assign CB_PE_input_width_1_num_0_I[12+:1] = I[12+:1];
	assign CB_PE_input_width_1_num_0_I[11+:1] = I[11+:1];
	assign CB_PE_input_width_1_num_0_I[10+:1] = I[10+:1];
	assign CB_PE_input_width_1_num_0_I[9+:1] = I[9+:1];
	assign CB_PE_input_width_1_num_0_I[8+:1] = I[8+:1];
	assign CB_PE_input_width_1_num_0_I[7+:1] = I[7+:1];
	assign CB_PE_input_width_1_num_0_I[6+:1] = I[6+:1];
	assign CB_PE_input_width_1_num_0_I[5+:1] = I[5+:1];
	assign CB_PE_input_width_1_num_0_I[4+:1] = I[4+:1];
	assign CB_PE_input_width_1_num_0_I[3+:1] = I[3+:1];
	assign CB_PE_input_width_1_num_0_I[2+:1] = I[2+:1];
	assign CB_PE_input_width_1_num_0_I[1+:1] = I[1+:1];
	assign CB_PE_input_width_1_num_0_I[0+:1] = I[0+:1];
	mux_aoi_ready_valid_const_21_1 CB_PE_input_width_1_num_0(
		.I(CB_PE_input_width_1_num_0_I),
		.O(CB_PE_input_width_1_num_0_O),
		.ready_in(ready_in),
		.ready_out(CB_PE_input_width_1_num_0_ready_out),
		.valid_in(valid_in),
		.valid_out(CB_PE_input_width_1_num_0_valid_out),
		.S(CB_PE_input_width_1_num_0_sel_value_O),
		.out_sel(CB_PE_input_width_1_num_0_out_sel)
	);
	SliceWrapper_6_0_1 CB_PE_input_width_1_num_0_enable_value(
		.I(config_reg_0_O),
		.O(CB_PE_input_width_1_num_0_enable_value_O)
	);
	SliceWrapper_6_1_6 CB_PE_input_width_1_num_0_sel_value(
		.I(config_reg_0_O),
		.O(CB_PE_input_width_1_num_0_sel_value_O)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_6_32_inst0$bit_const_0_None(.out(ZextWrapper_6_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
	assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, config_reg_0_O};
	mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O(
		.in(ZextWrapper_6_32_inst0$self_O_in),
		.out(ZextWrapper_6_32_inst0$self_O_out)
	);
	ConfigRegister_6_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	assign O = CB_PE_input_width_1_num_0_O;
	assign enable = CB_PE_input_width_1_num_0_enable_value_O[0];
	assign out_sel = CB_PE_input_width_1_num_0_out_sel;
	assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
	assign ready_out = CB_PE_input_width_1_num_0_ready_out;
	assign valid_out = CB_PE_input_width_1_num_0_valid_out;
endmodule
module CB_PE_input_width_17_num_3 (
	I,
	O,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	enable,
	out_sel,
	read_config_data,
	ready_in,
	ready_out,
	reset,
	valid_in,
	valid_out
);
	input [339:0] I;
	output wire [16:0] O;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output wire enable;
	output wire [31:0] out_sel;
	output wire [31:0] read_config_data;
	input ready_in;
	output wire ready_out;
	input reset;
	input [19:0] valid_in;
	output wire valid_out;
	wire [16:0] CB_PE_input_width_17_num_3_O;
	wire CB_PE_input_width_17_num_3_ready_out;
	wire CB_PE_input_width_17_num_3_valid_out;
	wire [31:0] CB_PE_input_width_17_num_3_out_sel;
	wire [0:0] CB_PE_input_width_17_num_3_enable_value_O;
	wire [4:0] CB_PE_input_width_17_num_3_sel_value_O;
	wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
	wire [5:0] config_reg_0_O;
	wire [339:0] CB_PE_input_width_17_num_3_I;
	assign CB_PE_input_width_17_num_3_I[323+:17] = I[323+:17];
	assign CB_PE_input_width_17_num_3_I[306+:17] = I[306+:17];
	assign CB_PE_input_width_17_num_3_I[289+:17] = I[289+:17];
	assign CB_PE_input_width_17_num_3_I[272+:17] = I[272+:17];
	assign CB_PE_input_width_17_num_3_I[255+:17] = I[255+:17];
	assign CB_PE_input_width_17_num_3_I[238+:17] = I[238+:17];
	assign CB_PE_input_width_17_num_3_I[221+:17] = I[221+:17];
	assign CB_PE_input_width_17_num_3_I[204+:17] = I[204+:17];
	assign CB_PE_input_width_17_num_3_I[187+:17] = I[187+:17];
	assign CB_PE_input_width_17_num_3_I[170+:17] = I[170+:17];
	assign CB_PE_input_width_17_num_3_I[153+:17] = I[153+:17];
	assign CB_PE_input_width_17_num_3_I[136+:17] = I[136+:17];
	assign CB_PE_input_width_17_num_3_I[119+:17] = I[119+:17];
	assign CB_PE_input_width_17_num_3_I[102+:17] = I[102+:17];
	assign CB_PE_input_width_17_num_3_I[85+:17] = I[85+:17];
	assign CB_PE_input_width_17_num_3_I[68+:17] = I[68+:17];
	assign CB_PE_input_width_17_num_3_I[51+:17] = I[51+:17];
	assign CB_PE_input_width_17_num_3_I[34+:17] = I[34+:17];
	assign CB_PE_input_width_17_num_3_I[17+:17] = I[17+:17];
	assign CB_PE_input_width_17_num_3_I[0+:17] = I[0+:17];
	mux_aoi_ready_valid_const_20_17 CB_PE_input_width_17_num_3(
		.I(CB_PE_input_width_17_num_3_I),
		.O(CB_PE_input_width_17_num_3_O),
		.ready_in(ready_in),
		.ready_out(CB_PE_input_width_17_num_3_ready_out),
		.valid_in(valid_in),
		.valid_out(CB_PE_input_width_17_num_3_valid_out),
		.S(CB_PE_input_width_17_num_3_sel_value_O),
		.out_sel(CB_PE_input_width_17_num_3_out_sel)
	);
	SliceWrapper_6_0_1 CB_PE_input_width_17_num_3_enable_value(
		.I(config_reg_0_O),
		.O(CB_PE_input_width_17_num_3_enable_value_O)
	);
	SliceWrapper_6_1_6 CB_PE_input_width_17_num_3_sel_value(
		.I(config_reg_0_O),
		.O(CB_PE_input_width_17_num_3_sel_value_O)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_6_32_inst0$bit_const_0_None(.out(ZextWrapper_6_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
	assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, config_reg_0_O};
	mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O(
		.in(ZextWrapper_6_32_inst0$self_O_in),
		.out(ZextWrapper_6_32_inst0$self_O_out)
	);
	ConfigRegister_6_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	assign O = CB_PE_input_width_17_num_3_O;
	assign enable = CB_PE_input_width_17_num_3_enable_value_O[0];
	assign out_sel = CB_PE_input_width_17_num_3_out_sel;
	assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
	assign ready_out = CB_PE_input_width_17_num_3_ready_out;
	assign valid_out = CB_PE_input_width_17_num_3_valid_out;
endmodule
module CB_PE_input_width_17_num_2 (
	I,
	O,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	enable,
	out_sel,
	read_config_data,
	ready_in,
	ready_out,
	reset,
	valid_in,
	valid_out
);
	input [356:0] I;
	output wire [16:0] O;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output wire enable;
	output wire [31:0] out_sel;
	output wire [31:0] read_config_data;
	input ready_in;
	output wire ready_out;
	input reset;
	input [20:0] valid_in;
	output wire valid_out;
	wire [16:0] CB_PE_input_width_17_num_2_O;
	wire CB_PE_input_width_17_num_2_ready_out;
	wire CB_PE_input_width_17_num_2_valid_out;
	wire [31:0] CB_PE_input_width_17_num_2_out_sel;
	wire [0:0] CB_PE_input_width_17_num_2_enable_value_O;
	wire [4:0] CB_PE_input_width_17_num_2_sel_value_O;
	wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
	wire [5:0] config_reg_0_O;
	wire [356:0] CB_PE_input_width_17_num_2_I;
	assign CB_PE_input_width_17_num_2_I[340+:17] = I[340+:17];
	assign CB_PE_input_width_17_num_2_I[323+:17] = I[323+:17];
	assign CB_PE_input_width_17_num_2_I[306+:17] = I[306+:17];
	assign CB_PE_input_width_17_num_2_I[289+:17] = I[289+:17];
	assign CB_PE_input_width_17_num_2_I[272+:17] = I[272+:17];
	assign CB_PE_input_width_17_num_2_I[255+:17] = I[255+:17];
	assign CB_PE_input_width_17_num_2_I[238+:17] = I[238+:17];
	assign CB_PE_input_width_17_num_2_I[221+:17] = I[221+:17];
	assign CB_PE_input_width_17_num_2_I[204+:17] = I[204+:17];
	assign CB_PE_input_width_17_num_2_I[187+:17] = I[187+:17];
	assign CB_PE_input_width_17_num_2_I[170+:17] = I[170+:17];
	assign CB_PE_input_width_17_num_2_I[153+:17] = I[153+:17];
	assign CB_PE_input_width_17_num_2_I[136+:17] = I[136+:17];
	assign CB_PE_input_width_17_num_2_I[119+:17] = I[119+:17];
	assign CB_PE_input_width_17_num_2_I[102+:17] = I[102+:17];
	assign CB_PE_input_width_17_num_2_I[85+:17] = I[85+:17];
	assign CB_PE_input_width_17_num_2_I[68+:17] = I[68+:17];
	assign CB_PE_input_width_17_num_2_I[51+:17] = I[51+:17];
	assign CB_PE_input_width_17_num_2_I[34+:17] = I[34+:17];
	assign CB_PE_input_width_17_num_2_I[17+:17] = I[17+:17];
	assign CB_PE_input_width_17_num_2_I[0+:17] = I[0+:17];
	mux_aoi_ready_valid_const_21_17 CB_PE_input_width_17_num_2(
		.I(CB_PE_input_width_17_num_2_I),
		.O(CB_PE_input_width_17_num_2_O),
		.ready_in(ready_in),
		.ready_out(CB_PE_input_width_17_num_2_ready_out),
		.valid_in(valid_in),
		.valid_out(CB_PE_input_width_17_num_2_valid_out),
		.S(CB_PE_input_width_17_num_2_sel_value_O),
		.out_sel(CB_PE_input_width_17_num_2_out_sel)
	);
	SliceWrapper_6_0_1 CB_PE_input_width_17_num_2_enable_value(
		.I(config_reg_0_O),
		.O(CB_PE_input_width_17_num_2_enable_value_O)
	);
	SliceWrapper_6_1_6 CB_PE_input_width_17_num_2_sel_value(
		.I(config_reg_0_O),
		.O(CB_PE_input_width_17_num_2_sel_value_O)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_6_32_inst0$bit_const_0_None(.out(ZextWrapper_6_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
	assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, config_reg_0_O};
	mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O(
		.in(ZextWrapper_6_32_inst0$self_O_in),
		.out(ZextWrapper_6_32_inst0$self_O_out)
	);
	ConfigRegister_6_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	assign O = CB_PE_input_width_17_num_2_O;
	assign enable = CB_PE_input_width_17_num_2_enable_value_O[0];
	assign out_sel = CB_PE_input_width_17_num_2_out_sel;
	assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
	assign ready_out = CB_PE_input_width_17_num_2_ready_out;
	assign valid_out = CB_PE_input_width_17_num_2_valid_out;
endmodule
module CB_PE_input_width_17_num_1 (
	I,
	O,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	enable,
	out_sel,
	read_config_data,
	ready_in,
	ready_out,
	reset,
	valid_in,
	valid_out
);
	input [356:0] I;
	output wire [16:0] O;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output wire enable;
	output wire [31:0] out_sel;
	output wire [31:0] read_config_data;
	input ready_in;
	output wire ready_out;
	input reset;
	input [20:0] valid_in;
	output wire valid_out;
	wire [16:0] CB_PE_input_width_17_num_1_O;
	wire CB_PE_input_width_17_num_1_ready_out;
	wire CB_PE_input_width_17_num_1_valid_out;
	wire [31:0] CB_PE_input_width_17_num_1_out_sel;
	wire [0:0] CB_PE_input_width_17_num_1_enable_value_O;
	wire [4:0] CB_PE_input_width_17_num_1_sel_value_O;
	wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
	wire [5:0] config_reg_0_O;
	wire [356:0] CB_PE_input_width_17_num_1_I;
	assign CB_PE_input_width_17_num_1_I[340+:17] = I[340+:17];
	assign CB_PE_input_width_17_num_1_I[323+:17] = I[323+:17];
	assign CB_PE_input_width_17_num_1_I[306+:17] = I[306+:17];
	assign CB_PE_input_width_17_num_1_I[289+:17] = I[289+:17];
	assign CB_PE_input_width_17_num_1_I[272+:17] = I[272+:17];
	assign CB_PE_input_width_17_num_1_I[255+:17] = I[255+:17];
	assign CB_PE_input_width_17_num_1_I[238+:17] = I[238+:17];
	assign CB_PE_input_width_17_num_1_I[221+:17] = I[221+:17];
	assign CB_PE_input_width_17_num_1_I[204+:17] = I[204+:17];
	assign CB_PE_input_width_17_num_1_I[187+:17] = I[187+:17];
	assign CB_PE_input_width_17_num_1_I[170+:17] = I[170+:17];
	assign CB_PE_input_width_17_num_1_I[153+:17] = I[153+:17];
	assign CB_PE_input_width_17_num_1_I[136+:17] = I[136+:17];
	assign CB_PE_input_width_17_num_1_I[119+:17] = I[119+:17];
	assign CB_PE_input_width_17_num_1_I[102+:17] = I[102+:17];
	assign CB_PE_input_width_17_num_1_I[85+:17] = I[85+:17];
	assign CB_PE_input_width_17_num_1_I[68+:17] = I[68+:17];
	assign CB_PE_input_width_17_num_1_I[51+:17] = I[51+:17];
	assign CB_PE_input_width_17_num_1_I[34+:17] = I[34+:17];
	assign CB_PE_input_width_17_num_1_I[17+:17] = I[17+:17];
	assign CB_PE_input_width_17_num_1_I[0+:17] = I[0+:17];
	mux_aoi_ready_valid_const_21_17 CB_PE_input_width_17_num_1(
		.I(CB_PE_input_width_17_num_1_I),
		.O(CB_PE_input_width_17_num_1_O),
		.ready_in(ready_in),
		.ready_out(CB_PE_input_width_17_num_1_ready_out),
		.valid_in(valid_in),
		.valid_out(CB_PE_input_width_17_num_1_valid_out),
		.S(CB_PE_input_width_17_num_1_sel_value_O),
		.out_sel(CB_PE_input_width_17_num_1_out_sel)
	);
	SliceWrapper_6_0_1 CB_PE_input_width_17_num_1_enable_value(
		.I(config_reg_0_O),
		.O(CB_PE_input_width_17_num_1_enable_value_O)
	);
	SliceWrapper_6_1_6 CB_PE_input_width_17_num_1_sel_value(
		.I(config_reg_0_O),
		.O(CB_PE_input_width_17_num_1_sel_value_O)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_6_32_inst0$bit_const_0_None(.out(ZextWrapper_6_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
	assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, config_reg_0_O};
	mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O(
		.in(ZextWrapper_6_32_inst0$self_O_in),
		.out(ZextWrapper_6_32_inst0$self_O_out)
	);
	ConfigRegister_6_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	assign O = CB_PE_input_width_17_num_1_O;
	assign enable = CB_PE_input_width_17_num_1_enable_value_O[0];
	assign out_sel = CB_PE_input_width_17_num_1_out_sel;
	assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
	assign ready_out = CB_PE_input_width_17_num_1_ready_out;
	assign valid_out = CB_PE_input_width_17_num_1_valid_out;
endmodule
module CB_PE_input_width_17_num_0 (
	I,
	O,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	enable,
	out_sel,
	read_config_data,
	ready_in,
	ready_out,
	reset,
	valid_in,
	valid_out
);
	input [356:0] I;
	output wire [16:0] O;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output wire enable;
	output wire [31:0] out_sel;
	output wire [31:0] read_config_data;
	input ready_in;
	output wire ready_out;
	input reset;
	input [20:0] valid_in;
	output wire valid_out;
	wire [16:0] CB_PE_input_width_17_num_0_O;
	wire CB_PE_input_width_17_num_0_ready_out;
	wire CB_PE_input_width_17_num_0_valid_out;
	wire [31:0] CB_PE_input_width_17_num_0_out_sel;
	wire [0:0] CB_PE_input_width_17_num_0_enable_value_O;
	wire [4:0] CB_PE_input_width_17_num_0_sel_value_O;
	wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
	wire [5:0] config_reg_0_O;
	wire [356:0] CB_PE_input_width_17_num_0_I;
	assign CB_PE_input_width_17_num_0_I[340+:17] = I[340+:17];
	assign CB_PE_input_width_17_num_0_I[323+:17] = I[323+:17];
	assign CB_PE_input_width_17_num_0_I[306+:17] = I[306+:17];
	assign CB_PE_input_width_17_num_0_I[289+:17] = I[289+:17];
	assign CB_PE_input_width_17_num_0_I[272+:17] = I[272+:17];
	assign CB_PE_input_width_17_num_0_I[255+:17] = I[255+:17];
	assign CB_PE_input_width_17_num_0_I[238+:17] = I[238+:17];
	assign CB_PE_input_width_17_num_0_I[221+:17] = I[221+:17];
	assign CB_PE_input_width_17_num_0_I[204+:17] = I[204+:17];
	assign CB_PE_input_width_17_num_0_I[187+:17] = I[187+:17];
	assign CB_PE_input_width_17_num_0_I[170+:17] = I[170+:17];
	assign CB_PE_input_width_17_num_0_I[153+:17] = I[153+:17];
	assign CB_PE_input_width_17_num_0_I[136+:17] = I[136+:17];
	assign CB_PE_input_width_17_num_0_I[119+:17] = I[119+:17];
	assign CB_PE_input_width_17_num_0_I[102+:17] = I[102+:17];
	assign CB_PE_input_width_17_num_0_I[85+:17] = I[85+:17];
	assign CB_PE_input_width_17_num_0_I[68+:17] = I[68+:17];
	assign CB_PE_input_width_17_num_0_I[51+:17] = I[51+:17];
	assign CB_PE_input_width_17_num_0_I[34+:17] = I[34+:17];
	assign CB_PE_input_width_17_num_0_I[17+:17] = I[17+:17];
	assign CB_PE_input_width_17_num_0_I[0+:17] = I[0+:17];
	mux_aoi_ready_valid_const_21_17 CB_PE_input_width_17_num_0(
		.I(CB_PE_input_width_17_num_0_I),
		.O(CB_PE_input_width_17_num_0_O),
		.ready_in(ready_in),
		.ready_out(CB_PE_input_width_17_num_0_ready_out),
		.valid_in(valid_in),
		.valid_out(CB_PE_input_width_17_num_0_valid_out),
		.S(CB_PE_input_width_17_num_0_sel_value_O),
		.out_sel(CB_PE_input_width_17_num_0_out_sel)
	);
	SliceWrapper_6_0_1 CB_PE_input_width_17_num_0_enable_value(
		.I(config_reg_0_O),
		.O(CB_PE_input_width_17_num_0_enable_value_O)
	);
	SliceWrapper_6_1_6 CB_PE_input_width_17_num_0_sel_value(
		.I(config_reg_0_O),
		.O(CB_PE_input_width_17_num_0_sel_value_O)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_6_32_inst0$bit_const_0_None(.out(ZextWrapper_6_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
	assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, config_reg_0_O};
	mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O(
		.in(ZextWrapper_6_32_inst0$self_O_in),
		.out(ZextWrapper_6_32_inst0$self_O_out)
	);
	ConfigRegister_6_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	assign O = CB_PE_input_width_17_num_0_O;
	assign enable = CB_PE_input_width_17_num_0_enable_value_O[0];
	assign out_sel = CB_PE_input_width_17_num_0_out_sel;
	assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
	assign ready_out = CB_PE_input_width_17_num_0_ready_out;
	assign valid_out = CB_PE_input_width_17_num_0_valid_out;
endmodule
module Tile_PE (
	SB_T0_EAST_SB_IN_B1,
	SB_T0_EAST_SB_IN_B17,
	SB_T0_EAST_SB_IN_B17_ready,
	SB_T0_EAST_SB_IN_B17_valid,
	SB_T0_EAST_SB_IN_B1_ready,
	SB_T0_EAST_SB_IN_B1_valid,
	SB_T0_EAST_SB_OUT_B1,
	SB_T0_EAST_SB_OUT_B17,
	SB_T0_EAST_SB_OUT_B17_ready,
	SB_T0_EAST_SB_OUT_B17_valid,
	SB_T0_EAST_SB_OUT_B1_ready,
	SB_T0_EAST_SB_OUT_B1_valid,
	SB_T0_NORTH_SB_IN_B1,
	SB_T0_NORTH_SB_IN_B17,
	SB_T0_NORTH_SB_IN_B17_ready,
	SB_T0_NORTH_SB_IN_B17_valid,
	SB_T0_NORTH_SB_IN_B1_ready,
	SB_T0_NORTH_SB_IN_B1_valid,
	SB_T0_NORTH_SB_OUT_B1,
	SB_T0_NORTH_SB_OUT_B17,
	SB_T0_NORTH_SB_OUT_B17_ready,
	SB_T0_NORTH_SB_OUT_B17_valid,
	SB_T0_NORTH_SB_OUT_B1_ready,
	SB_T0_NORTH_SB_OUT_B1_valid,
	SB_T0_SOUTH_SB_IN_B1,
	SB_T0_SOUTH_SB_IN_B17,
	SB_T0_SOUTH_SB_IN_B17_ready,
	SB_T0_SOUTH_SB_IN_B17_valid,
	SB_T0_SOUTH_SB_IN_B1_ready,
	SB_T0_SOUTH_SB_IN_B1_valid,
	SB_T0_SOUTH_SB_OUT_B1,
	SB_T0_SOUTH_SB_OUT_B17,
	SB_T0_SOUTH_SB_OUT_B17_ready,
	SB_T0_SOUTH_SB_OUT_B17_valid,
	SB_T0_SOUTH_SB_OUT_B1_ready,
	SB_T0_SOUTH_SB_OUT_B1_valid,
	SB_T0_WEST_SB_IN_B1,
	SB_T0_WEST_SB_IN_B17,
	SB_T0_WEST_SB_IN_B17_ready,
	SB_T0_WEST_SB_IN_B17_valid,
	SB_T0_WEST_SB_IN_B1_ready,
	SB_T0_WEST_SB_IN_B1_valid,
	SB_T0_WEST_SB_OUT_B1,
	SB_T0_WEST_SB_OUT_B17,
	SB_T0_WEST_SB_OUT_B17_ready,
	SB_T0_WEST_SB_OUT_B17_valid,
	SB_T0_WEST_SB_OUT_B1_ready,
	SB_T0_WEST_SB_OUT_B1_valid,
	SB_T1_EAST_SB_IN_B1,
	SB_T1_EAST_SB_IN_B17,
	SB_T1_EAST_SB_IN_B17_ready,
	SB_T1_EAST_SB_IN_B17_valid,
	SB_T1_EAST_SB_IN_B1_ready,
	SB_T1_EAST_SB_IN_B1_valid,
	SB_T1_EAST_SB_OUT_B1,
	SB_T1_EAST_SB_OUT_B17,
	SB_T1_EAST_SB_OUT_B17_ready,
	SB_T1_EAST_SB_OUT_B17_valid,
	SB_T1_EAST_SB_OUT_B1_ready,
	SB_T1_EAST_SB_OUT_B1_valid,
	SB_T1_NORTH_SB_IN_B1,
	SB_T1_NORTH_SB_IN_B17,
	SB_T1_NORTH_SB_IN_B17_ready,
	SB_T1_NORTH_SB_IN_B17_valid,
	SB_T1_NORTH_SB_IN_B1_ready,
	SB_T1_NORTH_SB_IN_B1_valid,
	SB_T1_NORTH_SB_OUT_B1,
	SB_T1_NORTH_SB_OUT_B17,
	SB_T1_NORTH_SB_OUT_B17_ready,
	SB_T1_NORTH_SB_OUT_B17_valid,
	SB_T1_NORTH_SB_OUT_B1_ready,
	SB_T1_NORTH_SB_OUT_B1_valid,
	SB_T1_SOUTH_SB_IN_B1,
	SB_T1_SOUTH_SB_IN_B17,
	SB_T1_SOUTH_SB_IN_B17_ready,
	SB_T1_SOUTH_SB_IN_B17_valid,
	SB_T1_SOUTH_SB_IN_B1_ready,
	SB_T1_SOUTH_SB_IN_B1_valid,
	SB_T1_SOUTH_SB_OUT_B1,
	SB_T1_SOUTH_SB_OUT_B17,
	SB_T1_SOUTH_SB_OUT_B17_ready,
	SB_T1_SOUTH_SB_OUT_B17_valid,
	SB_T1_SOUTH_SB_OUT_B1_ready,
	SB_T1_SOUTH_SB_OUT_B1_valid,
	SB_T1_WEST_SB_IN_B1,
	SB_T1_WEST_SB_IN_B17,
	SB_T1_WEST_SB_IN_B17_ready,
	SB_T1_WEST_SB_IN_B17_valid,
	SB_T1_WEST_SB_IN_B1_ready,
	SB_T1_WEST_SB_IN_B1_valid,
	SB_T1_WEST_SB_OUT_B1,
	SB_T1_WEST_SB_OUT_B17,
	SB_T1_WEST_SB_OUT_B17_ready,
	SB_T1_WEST_SB_OUT_B17_valid,
	SB_T1_WEST_SB_OUT_B1_ready,
	SB_T1_WEST_SB_OUT_B1_valid,
	SB_T2_EAST_SB_IN_B1,
	SB_T2_EAST_SB_IN_B17,
	SB_T2_EAST_SB_IN_B17_ready,
	SB_T2_EAST_SB_IN_B17_valid,
	SB_T2_EAST_SB_IN_B1_ready,
	SB_T2_EAST_SB_IN_B1_valid,
	SB_T2_EAST_SB_OUT_B1,
	SB_T2_EAST_SB_OUT_B17,
	SB_T2_EAST_SB_OUT_B17_ready,
	SB_T2_EAST_SB_OUT_B17_valid,
	SB_T2_EAST_SB_OUT_B1_ready,
	SB_T2_EAST_SB_OUT_B1_valid,
	SB_T2_NORTH_SB_IN_B1,
	SB_T2_NORTH_SB_IN_B17,
	SB_T2_NORTH_SB_IN_B17_ready,
	SB_T2_NORTH_SB_IN_B17_valid,
	SB_T2_NORTH_SB_IN_B1_ready,
	SB_T2_NORTH_SB_IN_B1_valid,
	SB_T2_NORTH_SB_OUT_B1,
	SB_T2_NORTH_SB_OUT_B17,
	SB_T2_NORTH_SB_OUT_B17_ready,
	SB_T2_NORTH_SB_OUT_B17_valid,
	SB_T2_NORTH_SB_OUT_B1_ready,
	SB_T2_NORTH_SB_OUT_B1_valid,
	SB_T2_SOUTH_SB_IN_B1,
	SB_T2_SOUTH_SB_IN_B17,
	SB_T2_SOUTH_SB_IN_B17_ready,
	SB_T2_SOUTH_SB_IN_B17_valid,
	SB_T2_SOUTH_SB_IN_B1_ready,
	SB_T2_SOUTH_SB_IN_B1_valid,
	SB_T2_SOUTH_SB_OUT_B1,
	SB_T2_SOUTH_SB_OUT_B17,
	SB_T2_SOUTH_SB_OUT_B17_ready,
	SB_T2_SOUTH_SB_OUT_B17_valid,
	SB_T2_SOUTH_SB_OUT_B1_ready,
	SB_T2_SOUTH_SB_OUT_B1_valid,
	SB_T2_WEST_SB_IN_B1,
	SB_T2_WEST_SB_IN_B17,
	SB_T2_WEST_SB_IN_B17_ready,
	SB_T2_WEST_SB_IN_B17_valid,
	SB_T2_WEST_SB_IN_B1_ready,
	SB_T2_WEST_SB_IN_B1_valid,
	SB_T2_WEST_SB_OUT_B1,
	SB_T2_WEST_SB_OUT_B17,
	SB_T2_WEST_SB_OUT_B17_ready,
	SB_T2_WEST_SB_OUT_B17_valid,
	SB_T2_WEST_SB_OUT_B1_ready,
	SB_T2_WEST_SB_OUT_B1_valid,
	SB_T3_EAST_SB_IN_B1,
	SB_T3_EAST_SB_IN_B17,
	SB_T3_EAST_SB_IN_B17_ready,
	SB_T3_EAST_SB_IN_B17_valid,
	SB_T3_EAST_SB_IN_B1_ready,
	SB_T3_EAST_SB_IN_B1_valid,
	SB_T3_EAST_SB_OUT_B1,
	SB_T3_EAST_SB_OUT_B17,
	SB_T3_EAST_SB_OUT_B17_ready,
	SB_T3_EAST_SB_OUT_B17_valid,
	SB_T3_EAST_SB_OUT_B1_ready,
	SB_T3_EAST_SB_OUT_B1_valid,
	SB_T3_NORTH_SB_IN_B1,
	SB_T3_NORTH_SB_IN_B17,
	SB_T3_NORTH_SB_IN_B17_ready,
	SB_T3_NORTH_SB_IN_B17_valid,
	SB_T3_NORTH_SB_IN_B1_ready,
	SB_T3_NORTH_SB_IN_B1_valid,
	SB_T3_NORTH_SB_OUT_B1,
	SB_T3_NORTH_SB_OUT_B17,
	SB_T3_NORTH_SB_OUT_B17_ready,
	SB_T3_NORTH_SB_OUT_B17_valid,
	SB_T3_NORTH_SB_OUT_B1_ready,
	SB_T3_NORTH_SB_OUT_B1_valid,
	SB_T3_SOUTH_SB_IN_B1,
	SB_T3_SOUTH_SB_IN_B17,
	SB_T3_SOUTH_SB_IN_B17_ready,
	SB_T3_SOUTH_SB_IN_B17_valid,
	SB_T3_SOUTH_SB_IN_B1_ready,
	SB_T3_SOUTH_SB_IN_B1_valid,
	SB_T3_SOUTH_SB_OUT_B1,
	SB_T3_SOUTH_SB_OUT_B17,
	SB_T3_SOUTH_SB_OUT_B17_ready,
	SB_T3_SOUTH_SB_OUT_B17_valid,
	SB_T3_SOUTH_SB_OUT_B1_ready,
	SB_T3_SOUTH_SB_OUT_B1_valid,
	SB_T3_WEST_SB_IN_B1,
	SB_T3_WEST_SB_IN_B17,
	SB_T3_WEST_SB_IN_B17_ready,
	SB_T3_WEST_SB_IN_B17_valid,
	SB_T3_WEST_SB_IN_B1_ready,
	SB_T3_WEST_SB_IN_B1_valid,
	SB_T3_WEST_SB_OUT_B1,
	SB_T3_WEST_SB_OUT_B17,
	SB_T3_WEST_SB_OUT_B17_ready,
	SB_T3_WEST_SB_OUT_B17_valid,
	SB_T3_WEST_SB_OUT_B1_ready,
	SB_T3_WEST_SB_OUT_B1_valid,
	SB_T4_EAST_SB_IN_B1,
	SB_T4_EAST_SB_IN_B17,
	SB_T4_EAST_SB_IN_B17_ready,
	SB_T4_EAST_SB_IN_B17_valid,
	SB_T4_EAST_SB_IN_B1_ready,
	SB_T4_EAST_SB_IN_B1_valid,
	SB_T4_EAST_SB_OUT_B1,
	SB_T4_EAST_SB_OUT_B17,
	SB_T4_EAST_SB_OUT_B17_ready,
	SB_T4_EAST_SB_OUT_B17_valid,
	SB_T4_EAST_SB_OUT_B1_ready,
	SB_T4_EAST_SB_OUT_B1_valid,
	SB_T4_NORTH_SB_IN_B1,
	SB_T4_NORTH_SB_IN_B17,
	SB_T4_NORTH_SB_IN_B17_ready,
	SB_T4_NORTH_SB_IN_B17_valid,
	SB_T4_NORTH_SB_IN_B1_ready,
	SB_T4_NORTH_SB_IN_B1_valid,
	SB_T4_NORTH_SB_OUT_B1,
	SB_T4_NORTH_SB_OUT_B17,
	SB_T4_NORTH_SB_OUT_B17_ready,
	SB_T4_NORTH_SB_OUT_B17_valid,
	SB_T4_NORTH_SB_OUT_B1_ready,
	SB_T4_NORTH_SB_OUT_B1_valid,
	SB_T4_SOUTH_SB_IN_B1,
	SB_T4_SOUTH_SB_IN_B17,
	SB_T4_SOUTH_SB_IN_B17_ready,
	SB_T4_SOUTH_SB_IN_B17_valid,
	SB_T4_SOUTH_SB_IN_B1_ready,
	SB_T4_SOUTH_SB_IN_B1_valid,
	SB_T4_SOUTH_SB_OUT_B1,
	SB_T4_SOUTH_SB_OUT_B17,
	SB_T4_SOUTH_SB_OUT_B17_ready,
	SB_T4_SOUTH_SB_OUT_B17_valid,
	SB_T4_SOUTH_SB_OUT_B1_ready,
	SB_T4_SOUTH_SB_OUT_B1_valid,
	SB_T4_WEST_SB_IN_B1,
	SB_T4_WEST_SB_IN_B17,
	SB_T4_WEST_SB_IN_B17_ready,
	SB_T4_WEST_SB_IN_B17_valid,
	SB_T4_WEST_SB_IN_B1_ready,
	SB_T4_WEST_SB_IN_B1_valid,
	SB_T4_WEST_SB_OUT_B1,
	SB_T4_WEST_SB_OUT_B17,
	SB_T4_WEST_SB_OUT_B17_ready,
	SB_T4_WEST_SB_OUT_B17_valid,
	SB_T4_WEST_SB_OUT_B1_ready,
	SB_T4_WEST_SB_OUT_B1_valid,
	clk,
	clk_out,
	clk_pass_through,
	clk_pass_through_out_bot,
	clk_pass_through_out_right,
	config_config_addr,
	config_config_data,
	config_out_config_addr,
	config_out_config_data,
	config_out_read,
	config_out_write,
	config_read,
	config_write,
	flush,
	flush_out,
	hi,
	lo,
	read_config_data,
	read_config_data_in,
	reset,
	reset_out,
	stall,
	stall_out,
	tile_id
);
	input [0:0] SB_T0_EAST_SB_IN_B1;
	input [16:0] SB_T0_EAST_SB_IN_B17;
	output wire SB_T0_EAST_SB_IN_B17_ready;
	input SB_T0_EAST_SB_IN_B17_valid;
	output wire SB_T0_EAST_SB_IN_B1_ready;
	input SB_T0_EAST_SB_IN_B1_valid;
	output wire [0:0] SB_T0_EAST_SB_OUT_B1;
	output wire [16:0] SB_T0_EAST_SB_OUT_B17;
	input SB_T0_EAST_SB_OUT_B17_ready;
	output wire SB_T0_EAST_SB_OUT_B17_valid;
	input SB_T0_EAST_SB_OUT_B1_ready;
	output wire SB_T0_EAST_SB_OUT_B1_valid;
	input [0:0] SB_T0_NORTH_SB_IN_B1;
	input [16:0] SB_T0_NORTH_SB_IN_B17;
	output wire SB_T0_NORTH_SB_IN_B17_ready;
	input SB_T0_NORTH_SB_IN_B17_valid;
	output wire SB_T0_NORTH_SB_IN_B1_ready;
	input SB_T0_NORTH_SB_IN_B1_valid;
	output wire [0:0] SB_T0_NORTH_SB_OUT_B1;
	output wire [16:0] SB_T0_NORTH_SB_OUT_B17;
	input SB_T0_NORTH_SB_OUT_B17_ready;
	output wire SB_T0_NORTH_SB_OUT_B17_valid;
	input SB_T0_NORTH_SB_OUT_B1_ready;
	output wire SB_T0_NORTH_SB_OUT_B1_valid;
	input [0:0] SB_T0_SOUTH_SB_IN_B1;
	input [16:0] SB_T0_SOUTH_SB_IN_B17;
	output wire SB_T0_SOUTH_SB_IN_B17_ready;
	input SB_T0_SOUTH_SB_IN_B17_valid;
	output wire SB_T0_SOUTH_SB_IN_B1_ready;
	input SB_T0_SOUTH_SB_IN_B1_valid;
	output wire [0:0] SB_T0_SOUTH_SB_OUT_B1;
	output wire [16:0] SB_T0_SOUTH_SB_OUT_B17;
	input SB_T0_SOUTH_SB_OUT_B17_ready;
	output wire SB_T0_SOUTH_SB_OUT_B17_valid;
	input SB_T0_SOUTH_SB_OUT_B1_ready;
	output wire SB_T0_SOUTH_SB_OUT_B1_valid;
	input [0:0] SB_T0_WEST_SB_IN_B1;
	input [16:0] SB_T0_WEST_SB_IN_B17;
	output wire SB_T0_WEST_SB_IN_B17_ready;
	input SB_T0_WEST_SB_IN_B17_valid;
	output wire SB_T0_WEST_SB_IN_B1_ready;
	input SB_T0_WEST_SB_IN_B1_valid;
	output wire [0:0] SB_T0_WEST_SB_OUT_B1;
	output wire [16:0] SB_T0_WEST_SB_OUT_B17;
	input SB_T0_WEST_SB_OUT_B17_ready;
	output wire SB_T0_WEST_SB_OUT_B17_valid;
	input SB_T0_WEST_SB_OUT_B1_ready;
	output wire SB_T0_WEST_SB_OUT_B1_valid;
	input [0:0] SB_T1_EAST_SB_IN_B1;
	input [16:0] SB_T1_EAST_SB_IN_B17;
	output wire SB_T1_EAST_SB_IN_B17_ready;
	input SB_T1_EAST_SB_IN_B17_valid;
	output wire SB_T1_EAST_SB_IN_B1_ready;
	input SB_T1_EAST_SB_IN_B1_valid;
	output wire [0:0] SB_T1_EAST_SB_OUT_B1;
	output wire [16:0] SB_T1_EAST_SB_OUT_B17;
	input SB_T1_EAST_SB_OUT_B17_ready;
	output wire SB_T1_EAST_SB_OUT_B17_valid;
	input SB_T1_EAST_SB_OUT_B1_ready;
	output wire SB_T1_EAST_SB_OUT_B1_valid;
	input [0:0] SB_T1_NORTH_SB_IN_B1;
	input [16:0] SB_T1_NORTH_SB_IN_B17;
	output wire SB_T1_NORTH_SB_IN_B17_ready;
	input SB_T1_NORTH_SB_IN_B17_valid;
	output wire SB_T1_NORTH_SB_IN_B1_ready;
	input SB_T1_NORTH_SB_IN_B1_valid;
	output wire [0:0] SB_T1_NORTH_SB_OUT_B1;
	output wire [16:0] SB_T1_NORTH_SB_OUT_B17;
	input SB_T1_NORTH_SB_OUT_B17_ready;
	output wire SB_T1_NORTH_SB_OUT_B17_valid;
	input SB_T1_NORTH_SB_OUT_B1_ready;
	output wire SB_T1_NORTH_SB_OUT_B1_valid;
	input [0:0] SB_T1_SOUTH_SB_IN_B1;
	input [16:0] SB_T1_SOUTH_SB_IN_B17;
	output wire SB_T1_SOUTH_SB_IN_B17_ready;
	input SB_T1_SOUTH_SB_IN_B17_valid;
	output wire SB_T1_SOUTH_SB_IN_B1_ready;
	input SB_T1_SOUTH_SB_IN_B1_valid;
	output wire [0:0] SB_T1_SOUTH_SB_OUT_B1;
	output wire [16:0] SB_T1_SOUTH_SB_OUT_B17;
	input SB_T1_SOUTH_SB_OUT_B17_ready;
	output wire SB_T1_SOUTH_SB_OUT_B17_valid;
	input SB_T1_SOUTH_SB_OUT_B1_ready;
	output wire SB_T1_SOUTH_SB_OUT_B1_valid;
	input [0:0] SB_T1_WEST_SB_IN_B1;
	input [16:0] SB_T1_WEST_SB_IN_B17;
	output wire SB_T1_WEST_SB_IN_B17_ready;
	input SB_T1_WEST_SB_IN_B17_valid;
	output wire SB_T1_WEST_SB_IN_B1_ready;
	input SB_T1_WEST_SB_IN_B1_valid;
	output wire [0:0] SB_T1_WEST_SB_OUT_B1;
	output wire [16:0] SB_T1_WEST_SB_OUT_B17;
	input SB_T1_WEST_SB_OUT_B17_ready;
	output wire SB_T1_WEST_SB_OUT_B17_valid;
	input SB_T1_WEST_SB_OUT_B1_ready;
	output wire SB_T1_WEST_SB_OUT_B1_valid;
	input [0:0] SB_T2_EAST_SB_IN_B1;
	input [16:0] SB_T2_EAST_SB_IN_B17;
	output wire SB_T2_EAST_SB_IN_B17_ready;
	input SB_T2_EAST_SB_IN_B17_valid;
	output wire SB_T2_EAST_SB_IN_B1_ready;
	input SB_T2_EAST_SB_IN_B1_valid;
	output wire [0:0] SB_T2_EAST_SB_OUT_B1;
	output wire [16:0] SB_T2_EAST_SB_OUT_B17;
	input SB_T2_EAST_SB_OUT_B17_ready;
	output wire SB_T2_EAST_SB_OUT_B17_valid;
	input SB_T2_EAST_SB_OUT_B1_ready;
	output wire SB_T2_EAST_SB_OUT_B1_valid;
	input [0:0] SB_T2_NORTH_SB_IN_B1;
	input [16:0] SB_T2_NORTH_SB_IN_B17;
	output wire SB_T2_NORTH_SB_IN_B17_ready;
	input SB_T2_NORTH_SB_IN_B17_valid;
	output wire SB_T2_NORTH_SB_IN_B1_ready;
	input SB_T2_NORTH_SB_IN_B1_valid;
	output wire [0:0] SB_T2_NORTH_SB_OUT_B1;
	output wire [16:0] SB_T2_NORTH_SB_OUT_B17;
	input SB_T2_NORTH_SB_OUT_B17_ready;
	output wire SB_T2_NORTH_SB_OUT_B17_valid;
	input SB_T2_NORTH_SB_OUT_B1_ready;
	output wire SB_T2_NORTH_SB_OUT_B1_valid;
	input [0:0] SB_T2_SOUTH_SB_IN_B1;
	input [16:0] SB_T2_SOUTH_SB_IN_B17;
	output wire SB_T2_SOUTH_SB_IN_B17_ready;
	input SB_T2_SOUTH_SB_IN_B17_valid;
	output wire SB_T2_SOUTH_SB_IN_B1_ready;
	input SB_T2_SOUTH_SB_IN_B1_valid;
	output wire [0:0] SB_T2_SOUTH_SB_OUT_B1;
	output wire [16:0] SB_T2_SOUTH_SB_OUT_B17;
	input SB_T2_SOUTH_SB_OUT_B17_ready;
	output wire SB_T2_SOUTH_SB_OUT_B17_valid;
	input SB_T2_SOUTH_SB_OUT_B1_ready;
	output wire SB_T2_SOUTH_SB_OUT_B1_valid;
	input [0:0] SB_T2_WEST_SB_IN_B1;
	input [16:0] SB_T2_WEST_SB_IN_B17;
	output wire SB_T2_WEST_SB_IN_B17_ready;
	input SB_T2_WEST_SB_IN_B17_valid;
	output wire SB_T2_WEST_SB_IN_B1_ready;
	input SB_T2_WEST_SB_IN_B1_valid;
	output wire [0:0] SB_T2_WEST_SB_OUT_B1;
	output wire [16:0] SB_T2_WEST_SB_OUT_B17;
	input SB_T2_WEST_SB_OUT_B17_ready;
	output wire SB_T2_WEST_SB_OUT_B17_valid;
	input SB_T2_WEST_SB_OUT_B1_ready;
	output wire SB_T2_WEST_SB_OUT_B1_valid;
	input [0:0] SB_T3_EAST_SB_IN_B1;
	input [16:0] SB_T3_EAST_SB_IN_B17;
	output wire SB_T3_EAST_SB_IN_B17_ready;
	input SB_T3_EAST_SB_IN_B17_valid;
	output wire SB_T3_EAST_SB_IN_B1_ready;
	input SB_T3_EAST_SB_IN_B1_valid;
	output wire [0:0] SB_T3_EAST_SB_OUT_B1;
	output wire [16:0] SB_T3_EAST_SB_OUT_B17;
	input SB_T3_EAST_SB_OUT_B17_ready;
	output wire SB_T3_EAST_SB_OUT_B17_valid;
	input SB_T3_EAST_SB_OUT_B1_ready;
	output wire SB_T3_EAST_SB_OUT_B1_valid;
	input [0:0] SB_T3_NORTH_SB_IN_B1;
	input [16:0] SB_T3_NORTH_SB_IN_B17;
	output wire SB_T3_NORTH_SB_IN_B17_ready;
	input SB_T3_NORTH_SB_IN_B17_valid;
	output wire SB_T3_NORTH_SB_IN_B1_ready;
	input SB_T3_NORTH_SB_IN_B1_valid;
	output wire [0:0] SB_T3_NORTH_SB_OUT_B1;
	output wire [16:0] SB_T3_NORTH_SB_OUT_B17;
	input SB_T3_NORTH_SB_OUT_B17_ready;
	output wire SB_T3_NORTH_SB_OUT_B17_valid;
	input SB_T3_NORTH_SB_OUT_B1_ready;
	output wire SB_T3_NORTH_SB_OUT_B1_valid;
	input [0:0] SB_T3_SOUTH_SB_IN_B1;
	input [16:0] SB_T3_SOUTH_SB_IN_B17;
	output wire SB_T3_SOUTH_SB_IN_B17_ready;
	input SB_T3_SOUTH_SB_IN_B17_valid;
	output wire SB_T3_SOUTH_SB_IN_B1_ready;
	input SB_T3_SOUTH_SB_IN_B1_valid;
	output wire [0:0] SB_T3_SOUTH_SB_OUT_B1;
	output wire [16:0] SB_T3_SOUTH_SB_OUT_B17;
	input SB_T3_SOUTH_SB_OUT_B17_ready;
	output wire SB_T3_SOUTH_SB_OUT_B17_valid;
	input SB_T3_SOUTH_SB_OUT_B1_ready;
	output wire SB_T3_SOUTH_SB_OUT_B1_valid;
	input [0:0] SB_T3_WEST_SB_IN_B1;
	input [16:0] SB_T3_WEST_SB_IN_B17;
	output wire SB_T3_WEST_SB_IN_B17_ready;
	input SB_T3_WEST_SB_IN_B17_valid;
	output wire SB_T3_WEST_SB_IN_B1_ready;
	input SB_T3_WEST_SB_IN_B1_valid;
	output wire [0:0] SB_T3_WEST_SB_OUT_B1;
	output wire [16:0] SB_T3_WEST_SB_OUT_B17;
	input SB_T3_WEST_SB_OUT_B17_ready;
	output wire SB_T3_WEST_SB_OUT_B17_valid;
	input SB_T3_WEST_SB_OUT_B1_ready;
	output wire SB_T3_WEST_SB_OUT_B1_valid;
	input [0:0] SB_T4_EAST_SB_IN_B1;
	input [16:0] SB_T4_EAST_SB_IN_B17;
	output wire SB_T4_EAST_SB_IN_B17_ready;
	input SB_T4_EAST_SB_IN_B17_valid;
	output wire SB_T4_EAST_SB_IN_B1_ready;
	input SB_T4_EAST_SB_IN_B1_valid;
	output wire [0:0] SB_T4_EAST_SB_OUT_B1;
	output wire [16:0] SB_T4_EAST_SB_OUT_B17;
	input SB_T4_EAST_SB_OUT_B17_ready;
	output wire SB_T4_EAST_SB_OUT_B17_valid;
	input SB_T4_EAST_SB_OUT_B1_ready;
	output wire SB_T4_EAST_SB_OUT_B1_valid;
	input [0:0] SB_T4_NORTH_SB_IN_B1;
	input [16:0] SB_T4_NORTH_SB_IN_B17;
	output wire SB_T4_NORTH_SB_IN_B17_ready;
	input SB_T4_NORTH_SB_IN_B17_valid;
	output wire SB_T4_NORTH_SB_IN_B1_ready;
	input SB_T4_NORTH_SB_IN_B1_valid;
	output wire [0:0] SB_T4_NORTH_SB_OUT_B1;
	output wire [16:0] SB_T4_NORTH_SB_OUT_B17;
	input SB_T4_NORTH_SB_OUT_B17_ready;
	output wire SB_T4_NORTH_SB_OUT_B17_valid;
	input SB_T4_NORTH_SB_OUT_B1_ready;
	output wire SB_T4_NORTH_SB_OUT_B1_valid;
	input [0:0] SB_T4_SOUTH_SB_IN_B1;
	input [16:0] SB_T4_SOUTH_SB_IN_B17;
	output wire SB_T4_SOUTH_SB_IN_B17_ready;
	input SB_T4_SOUTH_SB_IN_B17_valid;
	output wire SB_T4_SOUTH_SB_IN_B1_ready;
	input SB_T4_SOUTH_SB_IN_B1_valid;
	output wire [0:0] SB_T4_SOUTH_SB_OUT_B1;
	output wire [16:0] SB_T4_SOUTH_SB_OUT_B17;
	input SB_T4_SOUTH_SB_OUT_B17_ready;
	output wire SB_T4_SOUTH_SB_OUT_B17_valid;
	input SB_T4_SOUTH_SB_OUT_B1_ready;
	output wire SB_T4_SOUTH_SB_OUT_B1_valid;
	input [0:0] SB_T4_WEST_SB_IN_B1;
	input [16:0] SB_T4_WEST_SB_IN_B17;
	output wire SB_T4_WEST_SB_IN_B17_ready;
	input SB_T4_WEST_SB_IN_B17_valid;
	output wire SB_T4_WEST_SB_IN_B1_ready;
	input SB_T4_WEST_SB_IN_B1_valid;
	output wire [0:0] SB_T4_WEST_SB_OUT_B1;
	output wire [16:0] SB_T4_WEST_SB_OUT_B17;
	input SB_T4_WEST_SB_OUT_B17_ready;
	output wire SB_T4_WEST_SB_OUT_B17_valid;
	input SB_T4_WEST_SB_OUT_B1_ready;
	output wire SB_T4_WEST_SB_OUT_B1_valid;
	input clk;
	output wire clk_out;
	input clk_pass_through;
	output wire clk_pass_through_out_bot;
	output wire clk_pass_through_out_right;
	input [31:0] config_config_addr;
	input [31:0] config_config_data;
	output wire [31:0] config_out_config_addr;
	output wire [31:0] config_out_config_data;
	output wire [0:0] config_out_read;
	output wire [0:0] config_out_write;
	input [0:0] config_read;
	input [0:0] config_write;
	input [0:0] flush;
	output wire [0:0] flush_out;
	output wire [8:0] hi;
	output wire [7:0] lo;
	output wire [31:0] read_config_data;
	input [31:0] read_config_data_in;
	input reset;
	output wire reset_out;
	input [0:0] stall;
	output wire [0:0] stall_out;
	input [15:0] tile_id;
	wire [16:0] CB_PE_input_width_17_num_0_O;
	wire CB_PE_input_width_17_num_0_enable;
	wire [31:0] CB_PE_input_width_17_num_0_out_sel;
	wire [31:0] CB_PE_input_width_17_num_0_read_config_data;
	wire CB_PE_input_width_17_num_0_ready_out;
	wire CB_PE_input_width_17_num_0_valid_out;
	wire [16:0] CB_PE_input_width_17_num_1_O;
	wire CB_PE_input_width_17_num_1_enable;
	wire [31:0] CB_PE_input_width_17_num_1_out_sel;
	wire [31:0] CB_PE_input_width_17_num_1_read_config_data;
	wire CB_PE_input_width_17_num_1_ready_out;
	wire CB_PE_input_width_17_num_1_valid_out;
	wire [16:0] CB_PE_input_width_17_num_2_O;
	wire CB_PE_input_width_17_num_2_enable;
	wire [31:0] CB_PE_input_width_17_num_2_out_sel;
	wire [31:0] CB_PE_input_width_17_num_2_read_config_data;
	wire CB_PE_input_width_17_num_2_ready_out;
	wire CB_PE_input_width_17_num_2_valid_out;
	wire [16:0] CB_PE_input_width_17_num_3_O;
	wire CB_PE_input_width_17_num_3_enable;
	wire [31:0] CB_PE_input_width_17_num_3_out_sel;
	wire [31:0] CB_PE_input_width_17_num_3_read_config_data;
	wire CB_PE_input_width_17_num_3_ready_out;
	wire CB_PE_input_width_17_num_3_valid_out;
	wire [0:0] CB_PE_input_width_1_num_0_O;
	wire CB_PE_input_width_1_num_0_enable;
	wire [31:0] CB_PE_input_width_1_num_0_out_sel;
	wire [31:0] CB_PE_input_width_1_num_0_read_config_data;
	wire CB_PE_input_width_1_num_0_ready_out;
	wire CB_PE_input_width_1_num_0_valid_out;
	wire [0:0] CB_PE_input_width_1_num_1_O;
	wire CB_PE_input_width_1_num_1_enable;
	wire [31:0] CB_PE_input_width_1_num_1_out_sel;
	wire [31:0] CB_PE_input_width_1_num_1_read_config_data;
	wire CB_PE_input_width_1_num_1_ready_out;
	wire CB_PE_input_width_1_num_1_valid_out;
	wire [0:0] CB_PE_input_width_1_num_2_O;
	wire CB_PE_input_width_1_num_2_enable;
	wire [31:0] CB_PE_input_width_1_num_2_out_sel;
	wire [31:0] CB_PE_input_width_1_num_2_read_config_data;
	wire CB_PE_input_width_1_num_2_ready_out;
	wire CB_PE_input_width_1_num_2_valid_out;
	wire [16:0] CB_PondTop_input_width_17_num_0_O;
	wire CB_PondTop_input_width_17_num_0_enable;
	wire [31:0] CB_PondTop_input_width_17_num_0_out_sel;
	wire [31:0] CB_PondTop_input_width_17_num_0_read_config_data;
	wire CB_PondTop_input_width_17_num_0_ready_out;
	wire CB_PondTop_input_width_17_num_0_valid_out;
	wire [16:0] CB_PondTop_input_width_17_num_1_O;
	wire CB_PondTop_input_width_17_num_1_enable;
	wire [31:0] CB_PondTop_input_width_17_num_1_out_sel;
	wire [31:0] CB_PondTop_input_width_17_num_1_read_config_data;
	wire CB_PondTop_input_width_17_num_1_ready_out;
	wire CB_PondTop_input_width_17_num_1_valid_out;
	wire [0:0] CB_flush_O;
	wire CB_flush_enable;
	wire [31:0] CB_flush_out_sel;
	wire [31:0] CB_flush_read_config_data;
	wire CB_flush_ready_out;
	wire CB_flush_valid_out;
	wire DECODE_FEATURE_0_O;
	wire DECODE_FEATURE_1_O;
	wire DECODE_FEATURE_10_O;
	wire DECODE_FEATURE_11_O;
	wire DECODE_FEATURE_12_O;
	wire DECODE_FEATURE_13_O;
	wire DECODE_FEATURE_14_O;
	wire DECODE_FEATURE_15_O;
	wire DECODE_FEATURE_2_O;
	wire DECODE_FEATURE_3_O;
	wire DECODE_FEATURE_4_O;
	wire DECODE_FEATURE_5_O;
	wire DECODE_FEATURE_6_O;
	wire DECODE_FEATURE_7_O;
	wire DECODE_FEATURE_8_O;
	wire DECODE_FEATURE_9_O;
	wire FEATURE_AND_0_out;
	wire FEATURE_AND_1_out;
	wire FEATURE_AND_10_out;
	wire FEATURE_AND_11_out;
	wire FEATURE_AND_12_out;
	wire FEATURE_AND_13_out;
	wire FEATURE_AND_14_out;
	wire FEATURE_AND_15_out;
	wire FEATURE_AND_2_out;
	wire FEATURE_AND_3_out;
	wire FEATURE_AND_4_out;
	wire FEATURE_AND_5_out;
	wire FEATURE_AND_6_out;
	wire FEATURE_AND_7_out;
	wire FEATURE_AND_8_out;
	wire FEATURE_AND_9_out;
	wire [0:0] PE_inst0_PE_input_width_17_num_0_ready;
	wire [0:0] PE_inst0_PE_input_width_17_num_1_ready;
	wire [0:0] PE_inst0_PE_input_width_17_num_2_ready;
	wire [0:0] PE_inst0_PE_input_width_17_num_3_ready;
	wire PE_inst0_PE_input_width_1_num_0_ready;
	wire PE_inst0_PE_input_width_1_num_1_ready;
	wire PE_inst0_PE_input_width_1_num_2_ready;
	wire [16:0] PE_inst0_PE_output_width_17_num_0;
	wire [0:0] PE_inst0_PE_output_width_17_num_0_valid;
	wire [16:0] PE_inst0_PE_output_width_17_num_1;
	wire [0:0] PE_inst0_PE_output_width_17_num_1_valid;
	wire [16:0] PE_inst0_PE_output_width_17_num_2;
	wire [0:0] PE_inst0_PE_output_width_17_num_2_valid;
	wire [0:0] PE_inst0_PE_output_width_1_num_0;
	wire PE_inst0_PE_output_width_1_num_0_valid;
	wire [31:0] PE_inst0_read_config_data;
	wire [0:0] PE_output_width_17_num_0_loopback_valid_out;
	wire [0:0] PE_output_width_17_num_1_loopback_valid_out;
	wire [0:0] PE_output_width_17_num_2_loopback_valid_out;
	wire [0:0] PE_output_width_1_num_0_loopback_valid_out;
	wire PondCore_inst0_PondTop_input_width_17_num_0_ready;
	wire PondCore_inst0_PondTop_input_width_17_num_1_ready;
	wire [16:0] PondCore_inst0_PondTop_output_width_17_num_0;
	wire PondCore_inst0_PondTop_output_width_17_num_0_valid;
	wire [16:0] PondCore_inst0_PondTop_output_width_17_num_1;
	wire PondCore_inst0_PondTop_output_width_17_num_1_valid;
	wire [0:0] PondCore_inst0_PondTop_output_width_1_num_0;
	wire PondCore_inst0_PondTop_output_width_1_num_0_valid;
	wire [0:0] PondCore_inst0_PondTop_output_width_1_num_1;
	wire PondCore_inst0_PondTop_output_width_1_num_1_valid;
	wire [31:0] PondCore_inst0_read_config_data;
	wire [31:0] PondCore_inst0_read_config_data_1;
	wire [0:0] PondTop_output_width_17_num_0_loopback_valid_out;
	wire [0:0] PondTop_output_width_17_num_1_loopback_valid_out;
	wire [0:0] PondTop_output_width_1_num_0_loopback_valid_out;
	wire [0:0] PondTop_output_width_1_num_1_loopback_valid_out;
	wire [0:0] PowerDomainConfigReg_inst0_ps_en_out;
	wire [31:0] PowerDomainConfigReg_inst0_read_config_data;
	wire [31:0] PowerDomainOR_O;
	wire SB_ID0_5TRACKS_B17_PE_PE_output_width_17_num_0_ready_out;
	wire SB_ID0_5TRACKS_B17_PE_PE_output_width_17_num_1_ready_out;
	wire SB_ID0_5TRACKS_B17_PE_PE_output_width_17_num_2_ready_out;
	wire SB_ID0_5TRACKS_B17_PE_PondTop_output_width_17_num_0_ready_out;
	wire SB_ID0_5TRACKS_B17_PE_PondTop_output_width_17_num_1_ready_out;
	wire SB_ID0_5TRACKS_B17_PE_SB_T0_EAST_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T0_EAST_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T0_EAST_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_PE_SB_T0_EAST_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T0_EAST_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_PE_SB_T0_NORTH_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T0_NORTH_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T0_NORTH_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_PE_SB_T0_NORTH_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T0_NORTH_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_PE_SB_T0_SOUTH_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T0_SOUTH_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T0_SOUTH_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_PE_SB_T0_SOUTH_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T0_SOUTH_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_PE_SB_T0_WEST_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T0_WEST_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T0_WEST_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_PE_SB_T0_WEST_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T0_WEST_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_PE_SB_T1_EAST_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T1_EAST_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T1_EAST_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_PE_SB_T1_EAST_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T1_EAST_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_PE_SB_T1_NORTH_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T1_NORTH_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T1_NORTH_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_PE_SB_T1_NORTH_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T1_NORTH_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_PE_SB_T1_SOUTH_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T1_SOUTH_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T1_SOUTH_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_PE_SB_T1_SOUTH_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T1_SOUTH_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_PE_SB_T1_WEST_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T1_WEST_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T1_WEST_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_PE_SB_T1_WEST_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T1_WEST_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_PE_SB_T2_EAST_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T2_EAST_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T2_EAST_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_PE_SB_T2_EAST_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T2_EAST_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_PE_SB_T2_NORTH_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T2_NORTH_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T2_NORTH_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_PE_SB_T2_NORTH_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T2_NORTH_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_PE_SB_T2_SOUTH_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T2_SOUTH_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T2_SOUTH_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_PE_SB_T2_SOUTH_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T2_SOUTH_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_PE_SB_T2_WEST_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T2_WEST_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T2_WEST_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_PE_SB_T2_WEST_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T2_WEST_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_PE_SB_T3_EAST_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T3_EAST_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T3_EAST_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_PE_SB_T3_EAST_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T3_EAST_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_PE_SB_T3_NORTH_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T3_NORTH_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T3_NORTH_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_PE_SB_T3_NORTH_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T3_NORTH_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_PE_SB_T3_SOUTH_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T3_SOUTH_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T3_SOUTH_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_PE_SB_T3_SOUTH_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T3_SOUTH_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_PE_SB_T3_WEST_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T3_WEST_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T3_WEST_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_PE_SB_T3_WEST_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T3_WEST_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_PE_SB_T4_EAST_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T4_EAST_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T4_EAST_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_PE_SB_T4_EAST_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T4_EAST_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_PE_SB_T4_NORTH_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T4_NORTH_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T4_NORTH_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_PE_SB_T4_NORTH_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T4_NORTH_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_PE_SB_T4_SOUTH_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T4_SOUTH_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T4_SOUTH_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_PE_SB_T4_SOUTH_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T4_SOUTH_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_PE_SB_T4_WEST_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T4_WEST_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T4_WEST_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_PE_SB_T4_WEST_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_PE_SB_T4_WEST_SB_OUT_B17_valid_out;
	wire [31:0] SB_ID0_5TRACKS_B17_PE_read_config_data;
	wire SB_ID0_5TRACKS_B1_PE_PE_output_width_1_num_0_ready_out;
	wire SB_ID0_5TRACKS_B1_PE_PondTop_output_width_1_num_0_ready_out;
	wire SB_ID0_5TRACKS_B1_PE_PondTop_output_width_1_num_1_ready_out;
	wire SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_OUT_B1_valid_out;
	wire [31:0] SB_ID0_5TRACKS_B1_PE_read_config_data;
	wire SB_T0_EAST_SB_OUT_B17_ready_and_Z;
	wire SB_T0_EAST_SB_OUT_B1_ready_and_Z;
	wire SB_T0_NORTH_SB_OUT_B17_ready_and_Z;
	wire SB_T0_NORTH_SB_OUT_B1_ready_and_Z;
	wire SB_T0_SOUTH_SB_OUT_B17_ready_and_Z;
	wire SB_T0_SOUTH_SB_OUT_B1_ready_and_Z;
	wire SB_T0_WEST_SB_OUT_B17_ready_and_Z;
	wire SB_T0_WEST_SB_OUT_B1_ready_and_Z;
	wire SB_T1_EAST_SB_OUT_B17_ready_and_Z;
	wire SB_T1_EAST_SB_OUT_B1_ready_and_Z;
	wire SB_T1_NORTH_SB_OUT_B17_ready_and_Z;
	wire SB_T1_NORTH_SB_OUT_B1_ready_and_Z;
	wire SB_T1_SOUTH_SB_OUT_B17_ready_and_Z;
	wire SB_T1_SOUTH_SB_OUT_B1_ready_and_Z;
	wire SB_T1_WEST_SB_OUT_B17_ready_and_Z;
	wire SB_T1_WEST_SB_OUT_B1_ready_and_Z;
	wire SB_T2_EAST_SB_OUT_B17_ready_and_Z;
	wire SB_T2_EAST_SB_OUT_B1_ready_and_Z;
	wire SB_T2_NORTH_SB_OUT_B17_ready_and_Z;
	wire SB_T2_NORTH_SB_OUT_B1_ready_and_Z;
	wire SB_T2_SOUTH_SB_OUT_B17_ready_and_Z;
	wire SB_T2_SOUTH_SB_OUT_B1_ready_and_Z;
	wire SB_T2_WEST_SB_OUT_B17_ready_and_Z;
	wire SB_T2_WEST_SB_OUT_B1_ready_and_Z;
	wire SB_T3_EAST_SB_OUT_B17_ready_and_Z;
	wire SB_T3_EAST_SB_OUT_B1_ready_and_Z;
	wire SB_T3_NORTH_SB_OUT_B17_ready_and_Z;
	wire SB_T3_NORTH_SB_OUT_B1_ready_and_Z;
	wire SB_T3_SOUTH_SB_OUT_B17_ready_and_Z;
	wire SB_T3_SOUTH_SB_OUT_B1_ready_and_Z;
	wire SB_T3_WEST_SB_OUT_B17_ready_and_Z;
	wire SB_T3_WEST_SB_OUT_B1_ready_and_Z;
	wire SB_T4_EAST_SB_OUT_B17_ready_and_Z;
	wire SB_T4_EAST_SB_OUT_B1_ready_and_Z;
	wire SB_T4_NORTH_SB_OUT_B17_ready_and_Z;
	wire SB_T4_NORTH_SB_OUT_B1_ready_and_Z;
	wire SB_T4_SOUTH_SB_OUT_B17_ready_and_Z;
	wire SB_T4_SOUTH_SB_OUT_B1_ready_and_Z;
	wire SB_T4_WEST_SB_OUT_B17_ready_and_Z;
	wire SB_T4_WEST_SB_OUT_B1_ready_and_Z;
	wire and_inst0_out;
	wire and_inst1_out;
	wire bit_const_1_None_out;
	wire [7:0] const_0_8_out;
	wire [8:0] const_511_9_out;
	wire coreir_eq_16_inst0_out;
	wire coreir_wrapOutClock_inst0_out;
	wire coreir_wrapOutClock_inst1_out;
	wire [31:0] read_data_mux_O;
	wire [31:0] self_config_config_addr_out;
	wire [356:0] CB_PE_input_width_17_num_0_I;
	assign CB_PE_input_width_17_num_0_I[340+:17] = PondCore_inst0_PondTop_output_width_17_num_0;
	assign CB_PE_input_width_17_num_0_I[323+:17] = SB_T4_WEST_SB_IN_B17;
	assign CB_PE_input_width_17_num_0_I[306+:17] = SB_T4_EAST_SB_IN_B17;
	assign CB_PE_input_width_17_num_0_I[289+:17] = SB_T4_SOUTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_0_I[272+:17] = SB_T4_NORTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_0_I[255+:17] = SB_T3_WEST_SB_IN_B17;
	assign CB_PE_input_width_17_num_0_I[238+:17] = SB_T3_EAST_SB_IN_B17;
	assign CB_PE_input_width_17_num_0_I[221+:17] = SB_T3_SOUTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_0_I[204+:17] = SB_T3_NORTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_0_I[187+:17] = SB_T2_WEST_SB_IN_B17;
	assign CB_PE_input_width_17_num_0_I[170+:17] = SB_T2_EAST_SB_IN_B17;
	assign CB_PE_input_width_17_num_0_I[153+:17] = SB_T2_SOUTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_0_I[136+:17] = SB_T2_NORTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_0_I[119+:17] = SB_T1_WEST_SB_IN_B17;
	assign CB_PE_input_width_17_num_0_I[102+:17] = SB_T1_EAST_SB_IN_B17;
	assign CB_PE_input_width_17_num_0_I[85+:17] = SB_T1_SOUTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_0_I[68+:17] = SB_T1_NORTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_0_I[51+:17] = SB_T0_WEST_SB_IN_B17;
	assign CB_PE_input_width_17_num_0_I[34+:17] = SB_T0_EAST_SB_IN_B17;
	assign CB_PE_input_width_17_num_0_I[17+:17] = SB_T0_SOUTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_0_I[0+:17] = SB_T0_NORTH_SB_IN_B17;
	wire [20:0] CB_PE_input_width_17_num_0_valid_in;
	assign CB_PE_input_width_17_num_0_valid_in = {PondCore_inst0_PondTop_output_width_17_num_0_valid, SB_T4_WEST_SB_IN_B17_valid, SB_T4_EAST_SB_IN_B17_valid, SB_T4_SOUTH_SB_IN_B17_valid, SB_T4_NORTH_SB_IN_B17_valid, SB_T3_WEST_SB_IN_B17_valid, SB_T3_EAST_SB_IN_B17_valid, SB_T3_SOUTH_SB_IN_B17_valid, SB_T3_NORTH_SB_IN_B17_valid, SB_T2_WEST_SB_IN_B17_valid, SB_T2_EAST_SB_IN_B17_valid, SB_T2_SOUTH_SB_IN_B17_valid, SB_T2_NORTH_SB_IN_B17_valid, SB_T1_WEST_SB_IN_B17_valid, SB_T1_EAST_SB_IN_B17_valid, SB_T1_SOUTH_SB_IN_B17_valid, SB_T1_NORTH_SB_IN_B17_valid, SB_T0_WEST_SB_IN_B17_valid, SB_T0_EAST_SB_IN_B17_valid, SB_T0_SOUTH_SB_IN_B17_valid, SB_T0_NORTH_SB_IN_B17_valid};
	CB_PE_input_width_17_num_0 CB_PE_input_width_17_num_0(
		.I(CB_PE_input_width_17_num_0_I),
		.O(CB_PE_input_width_17_num_0_O),
		.clk(clk),
		.config_config_addr(self_config_config_addr_out[31:24]),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_3_out),
		.enable(CB_PE_input_width_17_num_0_enable),
		.out_sel(CB_PE_input_width_17_num_0_out_sel),
		.read_config_data(CB_PE_input_width_17_num_0_read_config_data),
		.ready_in(PE_inst0_PE_input_width_17_num_0_ready[0]),
		.ready_out(CB_PE_input_width_17_num_0_ready_out),
		.reset(reset),
		.valid_in(CB_PE_input_width_17_num_0_valid_in),
		.valid_out(CB_PE_input_width_17_num_0_valid_out)
	);
	wire [356:0] CB_PE_input_width_17_num_1_I;
	assign CB_PE_input_width_17_num_1_I[340+:17] = PondCore_inst0_PondTop_output_width_17_num_0;
	assign CB_PE_input_width_17_num_1_I[323+:17] = SB_T4_WEST_SB_IN_B17;
	assign CB_PE_input_width_17_num_1_I[306+:17] = SB_T4_EAST_SB_IN_B17;
	assign CB_PE_input_width_17_num_1_I[289+:17] = SB_T4_SOUTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_1_I[272+:17] = SB_T4_NORTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_1_I[255+:17] = SB_T3_WEST_SB_IN_B17;
	assign CB_PE_input_width_17_num_1_I[238+:17] = SB_T3_EAST_SB_IN_B17;
	assign CB_PE_input_width_17_num_1_I[221+:17] = SB_T3_SOUTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_1_I[204+:17] = SB_T3_NORTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_1_I[187+:17] = SB_T2_WEST_SB_IN_B17;
	assign CB_PE_input_width_17_num_1_I[170+:17] = SB_T2_EAST_SB_IN_B17;
	assign CB_PE_input_width_17_num_1_I[153+:17] = SB_T2_SOUTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_1_I[136+:17] = SB_T2_NORTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_1_I[119+:17] = SB_T1_WEST_SB_IN_B17;
	assign CB_PE_input_width_17_num_1_I[102+:17] = SB_T1_EAST_SB_IN_B17;
	assign CB_PE_input_width_17_num_1_I[85+:17] = SB_T1_SOUTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_1_I[68+:17] = SB_T1_NORTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_1_I[51+:17] = SB_T0_WEST_SB_IN_B17;
	assign CB_PE_input_width_17_num_1_I[34+:17] = SB_T0_EAST_SB_IN_B17;
	assign CB_PE_input_width_17_num_1_I[17+:17] = SB_T0_SOUTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_1_I[0+:17] = SB_T0_NORTH_SB_IN_B17;
	wire [20:0] CB_PE_input_width_17_num_1_valid_in;
	assign CB_PE_input_width_17_num_1_valid_in = {PondCore_inst0_PondTop_output_width_17_num_0_valid, SB_T4_WEST_SB_IN_B17_valid, SB_T4_EAST_SB_IN_B17_valid, SB_T4_SOUTH_SB_IN_B17_valid, SB_T4_NORTH_SB_IN_B17_valid, SB_T3_WEST_SB_IN_B17_valid, SB_T3_EAST_SB_IN_B17_valid, SB_T3_SOUTH_SB_IN_B17_valid, SB_T3_NORTH_SB_IN_B17_valid, SB_T2_WEST_SB_IN_B17_valid, SB_T2_EAST_SB_IN_B17_valid, SB_T2_SOUTH_SB_IN_B17_valid, SB_T2_NORTH_SB_IN_B17_valid, SB_T1_WEST_SB_IN_B17_valid, SB_T1_EAST_SB_IN_B17_valid, SB_T1_SOUTH_SB_IN_B17_valid, SB_T1_NORTH_SB_IN_B17_valid, SB_T0_WEST_SB_IN_B17_valid, SB_T0_EAST_SB_IN_B17_valid, SB_T0_SOUTH_SB_IN_B17_valid, SB_T0_NORTH_SB_IN_B17_valid};
	CB_PE_input_width_17_num_1 CB_PE_input_width_17_num_1(
		.I(CB_PE_input_width_17_num_1_I),
		.O(CB_PE_input_width_17_num_1_O),
		.clk(clk),
		.config_config_addr(self_config_config_addr_out[31:24]),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_4_out),
		.enable(CB_PE_input_width_17_num_1_enable),
		.out_sel(CB_PE_input_width_17_num_1_out_sel),
		.read_config_data(CB_PE_input_width_17_num_1_read_config_data),
		.ready_in(PE_inst0_PE_input_width_17_num_1_ready[0]),
		.ready_out(CB_PE_input_width_17_num_1_ready_out),
		.reset(reset),
		.valid_in(CB_PE_input_width_17_num_1_valid_in),
		.valid_out(CB_PE_input_width_17_num_1_valid_out)
	);
	wire [356:0] CB_PE_input_width_17_num_2_I;
	assign CB_PE_input_width_17_num_2_I[340+:17] = PondCore_inst0_PondTop_output_width_17_num_0;
	assign CB_PE_input_width_17_num_2_I[323+:17] = SB_T4_WEST_SB_IN_B17;
	assign CB_PE_input_width_17_num_2_I[306+:17] = SB_T4_EAST_SB_IN_B17;
	assign CB_PE_input_width_17_num_2_I[289+:17] = SB_T4_SOUTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_2_I[272+:17] = SB_T4_NORTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_2_I[255+:17] = SB_T3_WEST_SB_IN_B17;
	assign CB_PE_input_width_17_num_2_I[238+:17] = SB_T3_EAST_SB_IN_B17;
	assign CB_PE_input_width_17_num_2_I[221+:17] = SB_T3_SOUTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_2_I[204+:17] = SB_T3_NORTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_2_I[187+:17] = SB_T2_WEST_SB_IN_B17;
	assign CB_PE_input_width_17_num_2_I[170+:17] = SB_T2_EAST_SB_IN_B17;
	assign CB_PE_input_width_17_num_2_I[153+:17] = SB_T2_SOUTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_2_I[136+:17] = SB_T2_NORTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_2_I[119+:17] = SB_T1_WEST_SB_IN_B17;
	assign CB_PE_input_width_17_num_2_I[102+:17] = SB_T1_EAST_SB_IN_B17;
	assign CB_PE_input_width_17_num_2_I[85+:17] = SB_T1_SOUTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_2_I[68+:17] = SB_T1_NORTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_2_I[51+:17] = SB_T0_WEST_SB_IN_B17;
	assign CB_PE_input_width_17_num_2_I[34+:17] = SB_T0_EAST_SB_IN_B17;
	assign CB_PE_input_width_17_num_2_I[17+:17] = SB_T0_SOUTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_2_I[0+:17] = SB_T0_NORTH_SB_IN_B17;
	wire [20:0] CB_PE_input_width_17_num_2_valid_in;
	assign CB_PE_input_width_17_num_2_valid_in = {PondCore_inst0_PondTop_output_width_17_num_0_valid, SB_T4_WEST_SB_IN_B17_valid, SB_T4_EAST_SB_IN_B17_valid, SB_T4_SOUTH_SB_IN_B17_valid, SB_T4_NORTH_SB_IN_B17_valid, SB_T3_WEST_SB_IN_B17_valid, SB_T3_EAST_SB_IN_B17_valid, SB_T3_SOUTH_SB_IN_B17_valid, SB_T3_NORTH_SB_IN_B17_valid, SB_T2_WEST_SB_IN_B17_valid, SB_T2_EAST_SB_IN_B17_valid, SB_T2_SOUTH_SB_IN_B17_valid, SB_T2_NORTH_SB_IN_B17_valid, SB_T1_WEST_SB_IN_B17_valid, SB_T1_EAST_SB_IN_B17_valid, SB_T1_SOUTH_SB_IN_B17_valid, SB_T1_NORTH_SB_IN_B17_valid, SB_T0_WEST_SB_IN_B17_valid, SB_T0_EAST_SB_IN_B17_valid, SB_T0_SOUTH_SB_IN_B17_valid, SB_T0_NORTH_SB_IN_B17_valid};
	CB_PE_input_width_17_num_2 CB_PE_input_width_17_num_2(
		.I(CB_PE_input_width_17_num_2_I),
		.O(CB_PE_input_width_17_num_2_O),
		.clk(clk),
		.config_config_addr(self_config_config_addr_out[31:24]),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_5_out),
		.enable(CB_PE_input_width_17_num_2_enable),
		.out_sel(CB_PE_input_width_17_num_2_out_sel),
		.read_config_data(CB_PE_input_width_17_num_2_read_config_data),
		.ready_in(PE_inst0_PE_input_width_17_num_2_ready[0]),
		.ready_out(CB_PE_input_width_17_num_2_ready_out),
		.reset(reset),
		.valid_in(CB_PE_input_width_17_num_2_valid_in),
		.valid_out(CB_PE_input_width_17_num_2_valid_out)
	);
	wire [339:0] CB_PE_input_width_17_num_3_I;
	assign CB_PE_input_width_17_num_3_I[323+:17] = SB_T4_WEST_SB_IN_B17;
	assign CB_PE_input_width_17_num_3_I[306+:17] = SB_T4_EAST_SB_IN_B17;
	assign CB_PE_input_width_17_num_3_I[289+:17] = SB_T4_SOUTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_3_I[272+:17] = SB_T4_NORTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_3_I[255+:17] = SB_T3_WEST_SB_IN_B17;
	assign CB_PE_input_width_17_num_3_I[238+:17] = SB_T3_EAST_SB_IN_B17;
	assign CB_PE_input_width_17_num_3_I[221+:17] = SB_T3_SOUTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_3_I[204+:17] = SB_T3_NORTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_3_I[187+:17] = SB_T2_WEST_SB_IN_B17;
	assign CB_PE_input_width_17_num_3_I[170+:17] = SB_T2_EAST_SB_IN_B17;
	assign CB_PE_input_width_17_num_3_I[153+:17] = SB_T2_SOUTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_3_I[136+:17] = SB_T2_NORTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_3_I[119+:17] = SB_T1_WEST_SB_IN_B17;
	assign CB_PE_input_width_17_num_3_I[102+:17] = SB_T1_EAST_SB_IN_B17;
	assign CB_PE_input_width_17_num_3_I[85+:17] = SB_T1_SOUTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_3_I[68+:17] = SB_T1_NORTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_3_I[51+:17] = SB_T0_WEST_SB_IN_B17;
	assign CB_PE_input_width_17_num_3_I[34+:17] = SB_T0_EAST_SB_IN_B17;
	assign CB_PE_input_width_17_num_3_I[17+:17] = SB_T0_SOUTH_SB_IN_B17;
	assign CB_PE_input_width_17_num_3_I[0+:17] = SB_T0_NORTH_SB_IN_B17;
	wire [19:0] CB_PE_input_width_17_num_3_valid_in;
	assign CB_PE_input_width_17_num_3_valid_in = {SB_T4_WEST_SB_IN_B17_valid, SB_T4_EAST_SB_IN_B17_valid, SB_T4_SOUTH_SB_IN_B17_valid, SB_T4_NORTH_SB_IN_B17_valid, SB_T3_WEST_SB_IN_B17_valid, SB_T3_EAST_SB_IN_B17_valid, SB_T3_SOUTH_SB_IN_B17_valid, SB_T3_NORTH_SB_IN_B17_valid, SB_T2_WEST_SB_IN_B17_valid, SB_T2_EAST_SB_IN_B17_valid, SB_T2_SOUTH_SB_IN_B17_valid, SB_T2_NORTH_SB_IN_B17_valid, SB_T1_WEST_SB_IN_B17_valid, SB_T1_EAST_SB_IN_B17_valid, SB_T1_SOUTH_SB_IN_B17_valid, SB_T1_NORTH_SB_IN_B17_valid, SB_T0_WEST_SB_IN_B17_valid, SB_T0_EAST_SB_IN_B17_valid, SB_T0_SOUTH_SB_IN_B17_valid, SB_T0_NORTH_SB_IN_B17_valid};
	CB_PE_input_width_17_num_3 CB_PE_input_width_17_num_3(
		.I(CB_PE_input_width_17_num_3_I),
		.O(CB_PE_input_width_17_num_3_O),
		.clk(clk),
		.config_config_addr(self_config_config_addr_out[31:24]),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_6_out),
		.enable(CB_PE_input_width_17_num_3_enable),
		.out_sel(CB_PE_input_width_17_num_3_out_sel),
		.read_config_data(CB_PE_input_width_17_num_3_read_config_data),
		.ready_in(PE_inst0_PE_input_width_17_num_3_ready[0]),
		.ready_out(CB_PE_input_width_17_num_3_ready_out),
		.reset(reset),
		.valid_in(CB_PE_input_width_17_num_3_valid_in),
		.valid_out(CB_PE_input_width_17_num_3_valid_out)
	);
	wire [20:0] CB_PE_input_width_1_num_0_I;
	assign CB_PE_input_width_1_num_0_I[20+:1] = PondCore_inst0_PondTop_output_width_1_num_0;
	assign CB_PE_input_width_1_num_0_I[19+:1] = SB_T4_WEST_SB_IN_B1;
	assign CB_PE_input_width_1_num_0_I[18+:1] = SB_T4_EAST_SB_IN_B1;
	assign CB_PE_input_width_1_num_0_I[17+:1] = SB_T4_SOUTH_SB_IN_B1;
	assign CB_PE_input_width_1_num_0_I[16+:1] = SB_T4_NORTH_SB_IN_B1;
	assign CB_PE_input_width_1_num_0_I[15+:1] = SB_T3_WEST_SB_IN_B1;
	assign CB_PE_input_width_1_num_0_I[14+:1] = SB_T3_EAST_SB_IN_B1;
	assign CB_PE_input_width_1_num_0_I[13+:1] = SB_T3_SOUTH_SB_IN_B1;
	assign CB_PE_input_width_1_num_0_I[12+:1] = SB_T3_NORTH_SB_IN_B1;
	assign CB_PE_input_width_1_num_0_I[11+:1] = SB_T2_WEST_SB_IN_B1;
	assign CB_PE_input_width_1_num_0_I[10+:1] = SB_T2_EAST_SB_IN_B1;
	assign CB_PE_input_width_1_num_0_I[9+:1] = SB_T2_SOUTH_SB_IN_B1;
	assign CB_PE_input_width_1_num_0_I[8+:1] = SB_T2_NORTH_SB_IN_B1;
	assign CB_PE_input_width_1_num_0_I[7+:1] = SB_T1_WEST_SB_IN_B1;
	assign CB_PE_input_width_1_num_0_I[6+:1] = SB_T1_EAST_SB_IN_B1;
	assign CB_PE_input_width_1_num_0_I[5+:1] = SB_T1_SOUTH_SB_IN_B1;
	assign CB_PE_input_width_1_num_0_I[4+:1] = SB_T1_NORTH_SB_IN_B1;
	assign CB_PE_input_width_1_num_0_I[3+:1] = SB_T0_WEST_SB_IN_B1;
	assign CB_PE_input_width_1_num_0_I[2+:1] = SB_T0_EAST_SB_IN_B1;
	assign CB_PE_input_width_1_num_0_I[1+:1] = SB_T0_SOUTH_SB_IN_B1;
	assign CB_PE_input_width_1_num_0_I[0+:1] = SB_T0_NORTH_SB_IN_B1;
	wire [20:0] CB_PE_input_width_1_num_0_valid_in;
	assign CB_PE_input_width_1_num_0_valid_in = {PondCore_inst0_PondTop_output_width_1_num_0_valid, SB_T4_WEST_SB_IN_B1_valid, SB_T4_EAST_SB_IN_B1_valid, SB_T4_SOUTH_SB_IN_B1_valid, SB_T4_NORTH_SB_IN_B1_valid, SB_T3_WEST_SB_IN_B1_valid, SB_T3_EAST_SB_IN_B1_valid, SB_T3_SOUTH_SB_IN_B1_valid, SB_T3_NORTH_SB_IN_B1_valid, SB_T2_WEST_SB_IN_B1_valid, SB_T2_EAST_SB_IN_B1_valid, SB_T2_SOUTH_SB_IN_B1_valid, SB_T2_NORTH_SB_IN_B1_valid, SB_T1_WEST_SB_IN_B1_valid, SB_T1_EAST_SB_IN_B1_valid, SB_T1_SOUTH_SB_IN_B1_valid, SB_T1_NORTH_SB_IN_B1_valid, SB_T0_WEST_SB_IN_B1_valid, SB_T0_EAST_SB_IN_B1_valid, SB_T0_SOUTH_SB_IN_B1_valid, SB_T0_NORTH_SB_IN_B1_valid};
	CB_PE_input_width_1_num_0 CB_PE_input_width_1_num_0(
		.I(CB_PE_input_width_1_num_0_I),
		.O(CB_PE_input_width_1_num_0_O),
		.clk(clk),
		.config_config_addr(self_config_config_addr_out[31:24]),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_7_out),
		.enable(CB_PE_input_width_1_num_0_enable),
		.out_sel(CB_PE_input_width_1_num_0_out_sel),
		.read_config_data(CB_PE_input_width_1_num_0_read_config_data),
		.ready_in(PE_inst0_PE_input_width_1_num_0_ready),
		.ready_out(CB_PE_input_width_1_num_0_ready_out),
		.reset(reset),
		.valid_in(CB_PE_input_width_1_num_0_valid_in),
		.valid_out(CB_PE_input_width_1_num_0_valid_out)
	);
	wire [19:0] CB_PE_input_width_1_num_1_I;
	assign CB_PE_input_width_1_num_1_I[19+:1] = SB_T4_WEST_SB_IN_B1;
	assign CB_PE_input_width_1_num_1_I[18+:1] = SB_T4_EAST_SB_IN_B1;
	assign CB_PE_input_width_1_num_1_I[17+:1] = SB_T4_SOUTH_SB_IN_B1;
	assign CB_PE_input_width_1_num_1_I[16+:1] = SB_T4_NORTH_SB_IN_B1;
	assign CB_PE_input_width_1_num_1_I[15+:1] = SB_T3_WEST_SB_IN_B1;
	assign CB_PE_input_width_1_num_1_I[14+:1] = SB_T3_EAST_SB_IN_B1;
	assign CB_PE_input_width_1_num_1_I[13+:1] = SB_T3_SOUTH_SB_IN_B1;
	assign CB_PE_input_width_1_num_1_I[12+:1] = SB_T3_NORTH_SB_IN_B1;
	assign CB_PE_input_width_1_num_1_I[11+:1] = SB_T2_WEST_SB_IN_B1;
	assign CB_PE_input_width_1_num_1_I[10+:1] = SB_T2_EAST_SB_IN_B1;
	assign CB_PE_input_width_1_num_1_I[9+:1] = SB_T2_SOUTH_SB_IN_B1;
	assign CB_PE_input_width_1_num_1_I[8+:1] = SB_T2_NORTH_SB_IN_B1;
	assign CB_PE_input_width_1_num_1_I[7+:1] = SB_T1_WEST_SB_IN_B1;
	assign CB_PE_input_width_1_num_1_I[6+:1] = SB_T1_EAST_SB_IN_B1;
	assign CB_PE_input_width_1_num_1_I[5+:1] = SB_T1_SOUTH_SB_IN_B1;
	assign CB_PE_input_width_1_num_1_I[4+:1] = SB_T1_NORTH_SB_IN_B1;
	assign CB_PE_input_width_1_num_1_I[3+:1] = SB_T0_WEST_SB_IN_B1;
	assign CB_PE_input_width_1_num_1_I[2+:1] = SB_T0_EAST_SB_IN_B1;
	assign CB_PE_input_width_1_num_1_I[1+:1] = SB_T0_SOUTH_SB_IN_B1;
	assign CB_PE_input_width_1_num_1_I[0+:1] = SB_T0_NORTH_SB_IN_B1;
	wire [19:0] CB_PE_input_width_1_num_1_valid_in;
	assign CB_PE_input_width_1_num_1_valid_in = {SB_T4_WEST_SB_IN_B1_valid, SB_T4_EAST_SB_IN_B1_valid, SB_T4_SOUTH_SB_IN_B1_valid, SB_T4_NORTH_SB_IN_B1_valid, SB_T3_WEST_SB_IN_B1_valid, SB_T3_EAST_SB_IN_B1_valid, SB_T3_SOUTH_SB_IN_B1_valid, SB_T3_NORTH_SB_IN_B1_valid, SB_T2_WEST_SB_IN_B1_valid, SB_T2_EAST_SB_IN_B1_valid, SB_T2_SOUTH_SB_IN_B1_valid, SB_T2_NORTH_SB_IN_B1_valid, SB_T1_WEST_SB_IN_B1_valid, SB_T1_EAST_SB_IN_B1_valid, SB_T1_SOUTH_SB_IN_B1_valid, SB_T1_NORTH_SB_IN_B1_valid, SB_T0_WEST_SB_IN_B1_valid, SB_T0_EAST_SB_IN_B1_valid, SB_T0_SOUTH_SB_IN_B1_valid, SB_T0_NORTH_SB_IN_B1_valid};
	CB_PE_input_width_1_num_1 CB_PE_input_width_1_num_1(
		.I(CB_PE_input_width_1_num_1_I),
		.O(CB_PE_input_width_1_num_1_O),
		.clk(clk),
		.config_config_addr(self_config_config_addr_out[31:24]),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_8_out),
		.enable(CB_PE_input_width_1_num_1_enable),
		.out_sel(CB_PE_input_width_1_num_1_out_sel),
		.read_config_data(CB_PE_input_width_1_num_1_read_config_data),
		.ready_in(PE_inst0_PE_input_width_1_num_1_ready),
		.ready_out(CB_PE_input_width_1_num_1_ready_out),
		.reset(reset),
		.valid_in(CB_PE_input_width_1_num_1_valid_in),
		.valid_out(CB_PE_input_width_1_num_1_valid_out)
	);
	wire [19:0] CB_PE_input_width_1_num_2_I;
	assign CB_PE_input_width_1_num_2_I[19+:1] = SB_T4_WEST_SB_IN_B1;
	assign CB_PE_input_width_1_num_2_I[18+:1] = SB_T4_EAST_SB_IN_B1;
	assign CB_PE_input_width_1_num_2_I[17+:1] = SB_T4_SOUTH_SB_IN_B1;
	assign CB_PE_input_width_1_num_2_I[16+:1] = SB_T4_NORTH_SB_IN_B1;
	assign CB_PE_input_width_1_num_2_I[15+:1] = SB_T3_WEST_SB_IN_B1;
	assign CB_PE_input_width_1_num_2_I[14+:1] = SB_T3_EAST_SB_IN_B1;
	assign CB_PE_input_width_1_num_2_I[13+:1] = SB_T3_SOUTH_SB_IN_B1;
	assign CB_PE_input_width_1_num_2_I[12+:1] = SB_T3_NORTH_SB_IN_B1;
	assign CB_PE_input_width_1_num_2_I[11+:1] = SB_T2_WEST_SB_IN_B1;
	assign CB_PE_input_width_1_num_2_I[10+:1] = SB_T2_EAST_SB_IN_B1;
	assign CB_PE_input_width_1_num_2_I[9+:1] = SB_T2_SOUTH_SB_IN_B1;
	assign CB_PE_input_width_1_num_2_I[8+:1] = SB_T2_NORTH_SB_IN_B1;
	assign CB_PE_input_width_1_num_2_I[7+:1] = SB_T1_WEST_SB_IN_B1;
	assign CB_PE_input_width_1_num_2_I[6+:1] = SB_T1_EAST_SB_IN_B1;
	assign CB_PE_input_width_1_num_2_I[5+:1] = SB_T1_SOUTH_SB_IN_B1;
	assign CB_PE_input_width_1_num_2_I[4+:1] = SB_T1_NORTH_SB_IN_B1;
	assign CB_PE_input_width_1_num_2_I[3+:1] = SB_T0_WEST_SB_IN_B1;
	assign CB_PE_input_width_1_num_2_I[2+:1] = SB_T0_EAST_SB_IN_B1;
	assign CB_PE_input_width_1_num_2_I[1+:1] = SB_T0_SOUTH_SB_IN_B1;
	assign CB_PE_input_width_1_num_2_I[0+:1] = SB_T0_NORTH_SB_IN_B1;
	wire [19:0] CB_PE_input_width_1_num_2_valid_in;
	assign CB_PE_input_width_1_num_2_valid_in = {SB_T4_WEST_SB_IN_B1_valid, SB_T4_EAST_SB_IN_B1_valid, SB_T4_SOUTH_SB_IN_B1_valid, SB_T4_NORTH_SB_IN_B1_valid, SB_T3_WEST_SB_IN_B1_valid, SB_T3_EAST_SB_IN_B1_valid, SB_T3_SOUTH_SB_IN_B1_valid, SB_T3_NORTH_SB_IN_B1_valid, SB_T2_WEST_SB_IN_B1_valid, SB_T2_EAST_SB_IN_B1_valid, SB_T2_SOUTH_SB_IN_B1_valid, SB_T2_NORTH_SB_IN_B1_valid, SB_T1_WEST_SB_IN_B1_valid, SB_T1_EAST_SB_IN_B1_valid, SB_T1_SOUTH_SB_IN_B1_valid, SB_T1_NORTH_SB_IN_B1_valid, SB_T0_WEST_SB_IN_B1_valid, SB_T0_EAST_SB_IN_B1_valid, SB_T0_SOUTH_SB_IN_B1_valid, SB_T0_NORTH_SB_IN_B1_valid};
	CB_PE_input_width_1_num_2 CB_PE_input_width_1_num_2(
		.I(CB_PE_input_width_1_num_2_I),
		.O(CB_PE_input_width_1_num_2_O),
		.clk(clk),
		.config_config_addr(self_config_config_addr_out[31:24]),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_9_out),
		.enable(CB_PE_input_width_1_num_2_enable),
		.out_sel(CB_PE_input_width_1_num_2_out_sel),
		.read_config_data(CB_PE_input_width_1_num_2_read_config_data),
		.ready_in(PE_inst0_PE_input_width_1_num_2_ready),
		.ready_out(CB_PE_input_width_1_num_2_ready_out),
		.reset(reset),
		.valid_in(CB_PE_input_width_1_num_2_valid_in),
		.valid_out(CB_PE_input_width_1_num_2_valid_out)
	);
	wire [356:0] CB_PondTop_input_width_17_num_0_I;
	assign CB_PondTop_input_width_17_num_0_I[340+:17] = PE_inst0_PE_output_width_17_num_0;
	assign CB_PondTop_input_width_17_num_0_I[323+:17] = SB_T4_WEST_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_0_I[306+:17] = SB_T4_EAST_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_0_I[289+:17] = SB_T4_SOUTH_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_0_I[272+:17] = SB_T4_NORTH_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_0_I[255+:17] = SB_T3_WEST_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_0_I[238+:17] = SB_T3_EAST_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_0_I[221+:17] = SB_T3_SOUTH_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_0_I[204+:17] = SB_T3_NORTH_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_0_I[187+:17] = SB_T2_WEST_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_0_I[170+:17] = SB_T2_EAST_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_0_I[153+:17] = SB_T2_SOUTH_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_0_I[136+:17] = SB_T2_NORTH_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_0_I[119+:17] = SB_T1_WEST_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_0_I[102+:17] = SB_T1_EAST_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_0_I[85+:17] = SB_T1_SOUTH_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_0_I[68+:17] = SB_T1_NORTH_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_0_I[51+:17] = SB_T0_WEST_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_0_I[34+:17] = SB_T0_EAST_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_0_I[17+:17] = SB_T0_SOUTH_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_0_I[0+:17] = SB_T0_NORTH_SB_IN_B17;
	wire [20:0] CB_PondTop_input_width_17_num_0_valid_in;
	assign CB_PondTop_input_width_17_num_0_valid_in = {PE_inst0_PE_output_width_17_num_0_valid[0], SB_T4_WEST_SB_IN_B17_valid, SB_T4_EAST_SB_IN_B17_valid, SB_T4_SOUTH_SB_IN_B17_valid, SB_T4_NORTH_SB_IN_B17_valid, SB_T3_WEST_SB_IN_B17_valid, SB_T3_EAST_SB_IN_B17_valid, SB_T3_SOUTH_SB_IN_B17_valid, SB_T3_NORTH_SB_IN_B17_valid, SB_T2_WEST_SB_IN_B17_valid, SB_T2_EAST_SB_IN_B17_valid, SB_T2_SOUTH_SB_IN_B17_valid, SB_T2_NORTH_SB_IN_B17_valid, SB_T1_WEST_SB_IN_B17_valid, SB_T1_EAST_SB_IN_B17_valid, SB_T1_SOUTH_SB_IN_B17_valid, SB_T1_NORTH_SB_IN_B17_valid, SB_T0_WEST_SB_IN_B17_valid, SB_T0_EAST_SB_IN_B17_valid, SB_T0_SOUTH_SB_IN_B17_valid, SB_T0_NORTH_SB_IN_B17_valid};
	CB_PondTop_input_width_17_num_0 CB_PondTop_input_width_17_num_0(
		.I(CB_PondTop_input_width_17_num_0_I),
		.O(CB_PondTop_input_width_17_num_0_O),
		.clk(clk),
		.config_config_addr(self_config_config_addr_out[31:24]),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_10_out),
		.enable(CB_PondTop_input_width_17_num_0_enable),
		.out_sel(CB_PondTop_input_width_17_num_0_out_sel),
		.read_config_data(CB_PondTop_input_width_17_num_0_read_config_data),
		.ready_in(PondCore_inst0_PondTop_input_width_17_num_0_ready),
		.ready_out(CB_PondTop_input_width_17_num_0_ready_out),
		.reset(reset),
		.valid_in(CB_PondTop_input_width_17_num_0_valid_in),
		.valid_out(CB_PondTop_input_width_17_num_0_valid_out)
	);
	wire [356:0] CB_PondTop_input_width_17_num_1_I;
	assign CB_PondTop_input_width_17_num_1_I[340+:17] = PE_inst0_PE_output_width_17_num_0;
	assign CB_PondTop_input_width_17_num_1_I[323+:17] = SB_T4_WEST_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_1_I[306+:17] = SB_T4_EAST_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_1_I[289+:17] = SB_T4_SOUTH_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_1_I[272+:17] = SB_T4_NORTH_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_1_I[255+:17] = SB_T3_WEST_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_1_I[238+:17] = SB_T3_EAST_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_1_I[221+:17] = SB_T3_SOUTH_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_1_I[204+:17] = SB_T3_NORTH_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_1_I[187+:17] = SB_T2_WEST_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_1_I[170+:17] = SB_T2_EAST_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_1_I[153+:17] = SB_T2_SOUTH_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_1_I[136+:17] = SB_T2_NORTH_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_1_I[119+:17] = SB_T1_WEST_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_1_I[102+:17] = SB_T1_EAST_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_1_I[85+:17] = SB_T1_SOUTH_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_1_I[68+:17] = SB_T1_NORTH_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_1_I[51+:17] = SB_T0_WEST_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_1_I[34+:17] = SB_T0_EAST_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_1_I[17+:17] = SB_T0_SOUTH_SB_IN_B17;
	assign CB_PondTop_input_width_17_num_1_I[0+:17] = SB_T0_NORTH_SB_IN_B17;
	wire [20:0] CB_PondTop_input_width_17_num_1_valid_in;
	assign CB_PondTop_input_width_17_num_1_valid_in = {PE_inst0_PE_output_width_17_num_0_valid[0], SB_T4_WEST_SB_IN_B17_valid, SB_T4_EAST_SB_IN_B17_valid, SB_T4_SOUTH_SB_IN_B17_valid, SB_T4_NORTH_SB_IN_B17_valid, SB_T3_WEST_SB_IN_B17_valid, SB_T3_EAST_SB_IN_B17_valid, SB_T3_SOUTH_SB_IN_B17_valid, SB_T3_NORTH_SB_IN_B17_valid, SB_T2_WEST_SB_IN_B17_valid, SB_T2_EAST_SB_IN_B17_valid, SB_T2_SOUTH_SB_IN_B17_valid, SB_T2_NORTH_SB_IN_B17_valid, SB_T1_WEST_SB_IN_B17_valid, SB_T1_EAST_SB_IN_B17_valid, SB_T1_SOUTH_SB_IN_B17_valid, SB_T1_NORTH_SB_IN_B17_valid, SB_T0_WEST_SB_IN_B17_valid, SB_T0_EAST_SB_IN_B17_valid, SB_T0_SOUTH_SB_IN_B17_valid, SB_T0_NORTH_SB_IN_B17_valid};
	CB_PondTop_input_width_17_num_1 CB_PondTop_input_width_17_num_1(
		.I(CB_PondTop_input_width_17_num_1_I),
		.O(CB_PondTop_input_width_17_num_1_O),
		.clk(clk),
		.config_config_addr(self_config_config_addr_out[31:24]),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_11_out),
		.enable(CB_PondTop_input_width_17_num_1_enable),
		.out_sel(CB_PondTop_input_width_17_num_1_out_sel),
		.read_config_data(CB_PondTop_input_width_17_num_1_read_config_data),
		.ready_in(PondCore_inst0_PondTop_input_width_17_num_1_ready),
		.ready_out(CB_PondTop_input_width_17_num_1_ready_out),
		.reset(reset),
		.valid_in(CB_PondTop_input_width_17_num_1_valid_in),
		.valid_out(CB_PondTop_input_width_17_num_1_valid_out)
	);
	wire [19:0] CB_flush_I;
	assign CB_flush_I[19+:1] = SB_T4_WEST_SB_IN_B1;
	assign CB_flush_I[18+:1] = SB_T4_EAST_SB_IN_B1;
	assign CB_flush_I[17+:1] = SB_T4_SOUTH_SB_IN_B1;
	assign CB_flush_I[16+:1] = SB_T4_NORTH_SB_IN_B1;
	assign CB_flush_I[15+:1] = SB_T3_WEST_SB_IN_B1;
	assign CB_flush_I[14+:1] = SB_T3_EAST_SB_IN_B1;
	assign CB_flush_I[13+:1] = SB_T3_SOUTH_SB_IN_B1;
	assign CB_flush_I[12+:1] = SB_T3_NORTH_SB_IN_B1;
	assign CB_flush_I[11+:1] = SB_T2_WEST_SB_IN_B1;
	assign CB_flush_I[10+:1] = SB_T2_EAST_SB_IN_B1;
	assign CB_flush_I[9+:1] = SB_T2_SOUTH_SB_IN_B1;
	assign CB_flush_I[8+:1] = SB_T2_NORTH_SB_IN_B1;
	assign CB_flush_I[7+:1] = SB_T1_WEST_SB_IN_B1;
	assign CB_flush_I[6+:1] = SB_T1_EAST_SB_IN_B1;
	assign CB_flush_I[5+:1] = SB_T1_SOUTH_SB_IN_B1;
	assign CB_flush_I[4+:1] = SB_T1_NORTH_SB_IN_B1;
	assign CB_flush_I[3+:1] = SB_T0_WEST_SB_IN_B1;
	assign CB_flush_I[2+:1] = SB_T0_EAST_SB_IN_B1;
	assign CB_flush_I[1+:1] = SB_T0_SOUTH_SB_IN_B1;
	assign CB_flush_I[0+:1] = SB_T0_NORTH_SB_IN_B1;
	wire [19:0] CB_flush_valid_in;
	assign CB_flush_valid_in = {SB_T4_WEST_SB_IN_B1_valid, SB_T4_EAST_SB_IN_B1_valid, SB_T4_SOUTH_SB_IN_B1_valid, SB_T4_NORTH_SB_IN_B1_valid, SB_T3_WEST_SB_IN_B1_valid, SB_T3_EAST_SB_IN_B1_valid, SB_T3_SOUTH_SB_IN_B1_valid, SB_T3_NORTH_SB_IN_B1_valid, SB_T2_WEST_SB_IN_B1_valid, SB_T2_EAST_SB_IN_B1_valid, SB_T2_SOUTH_SB_IN_B1_valid, SB_T2_NORTH_SB_IN_B1_valid, SB_T1_WEST_SB_IN_B1_valid, SB_T1_EAST_SB_IN_B1_valid, SB_T1_SOUTH_SB_IN_B1_valid, SB_T1_NORTH_SB_IN_B1_valid, SB_T0_WEST_SB_IN_B1_valid, SB_T0_EAST_SB_IN_B1_valid, SB_T0_SOUTH_SB_IN_B1_valid, SB_T0_NORTH_SB_IN_B1_valid};
	CB_flush CB_flush(
		.I(CB_flush_I),
		.O(CB_flush_O),
		.clk(clk),
		.config_config_addr(self_config_config_addr_out[31:24]),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_12_out),
		.enable(CB_flush_enable),
		.out_sel(CB_flush_out_sel),
		.read_config_data(CB_flush_read_config_data),
		.ready_in(bit_const_1_None_out),
		.ready_out(CB_flush_ready_out),
		.reset(reset),
		.valid_in(CB_flush_valid_in),
		.valid_out(CB_flush_valid_out)
	);
	Decode08 DECODE_FEATURE_0(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_0_O)
	);
	Decode18 DECODE_FEATURE_1(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_1_O)
	);
	Decode108 DECODE_FEATURE_10(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_10_O)
	);
	Decode118 DECODE_FEATURE_11(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_11_O)
	);
	Decode128 DECODE_FEATURE_12(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_12_O)
	);
	Decode138 DECODE_FEATURE_13(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_13_O)
	);
	Decode148 DECODE_FEATURE_14(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_14_O)
	);
	Decode158 DECODE_FEATURE_15(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_15_O)
	);
	Decode28 DECODE_FEATURE_2(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_2_O)
	);
	Decode38 DECODE_FEATURE_3(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_3_O)
	);
	Decode48 DECODE_FEATURE_4(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_4_O)
	);
	Decode58 DECODE_FEATURE_5(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_5_O)
	);
	Decode68 DECODE_FEATURE_6(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_6_O)
	);
	Decode78 DECODE_FEATURE_7(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_7_O)
	);
	Decode88 DECODE_FEATURE_8(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_8_O)
	);
	Decode98 DECODE_FEATURE_9(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_9_O)
	);
	corebit_and FEATURE_AND_0(
		.in0(DECODE_FEATURE_0_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_0_out)
	);
	corebit_and FEATURE_AND_1(
		.in0(DECODE_FEATURE_1_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_1_out)
	);
	corebit_and FEATURE_AND_10(
		.in0(DECODE_FEATURE_10_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_10_out)
	);
	corebit_and FEATURE_AND_11(
		.in0(DECODE_FEATURE_11_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_11_out)
	);
	corebit_and FEATURE_AND_12(
		.in0(DECODE_FEATURE_12_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_12_out)
	);
	corebit_and FEATURE_AND_13(
		.in0(DECODE_FEATURE_13_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_13_out)
	);
	corebit_and FEATURE_AND_14(
		.in0(DECODE_FEATURE_14_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_14_out)
	);
	corebit_and FEATURE_AND_15(
		.in0(DECODE_FEATURE_15_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_15_out)
	);
	corebit_and FEATURE_AND_2(
		.in0(DECODE_FEATURE_2_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_2_out)
	);
	corebit_and FEATURE_AND_3(
		.in0(DECODE_FEATURE_3_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_3_out)
	);
	corebit_and FEATURE_AND_4(
		.in0(DECODE_FEATURE_4_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_4_out)
	);
	corebit_and FEATURE_AND_5(
		.in0(DECODE_FEATURE_5_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_5_out)
	);
	corebit_and FEATURE_AND_6(
		.in0(DECODE_FEATURE_6_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_6_out)
	);
	corebit_and FEATURE_AND_7(
		.in0(DECODE_FEATURE_7_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_7_out)
	);
	corebit_and FEATURE_AND_8(
		.in0(DECODE_FEATURE_8_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_8_out)
	);
	corebit_and FEATURE_AND_9(
		.in0(DECODE_FEATURE_9_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_9_out)
	);
	PE PE_inst0(
		.PE_input_width_17_num_0(CB_PE_input_width_17_num_0_O),
		.PE_input_width_17_num_0_ready(PE_inst0_PE_input_width_17_num_0_ready),
		.PE_input_width_17_num_0_valid(CB_PE_input_width_17_num_0_valid_out),
		.PE_input_width_17_num_1(CB_PE_input_width_17_num_1_O),
		.PE_input_width_17_num_1_ready(PE_inst0_PE_input_width_17_num_1_ready),
		.PE_input_width_17_num_1_valid(CB_PE_input_width_17_num_1_valid_out),
		.PE_input_width_17_num_2(CB_PE_input_width_17_num_2_O),
		.PE_input_width_17_num_2_ready(PE_inst0_PE_input_width_17_num_2_ready),
		.PE_input_width_17_num_2_valid(CB_PE_input_width_17_num_2_valid_out),
		.PE_input_width_17_num_3(CB_PE_input_width_17_num_3_O),
		.PE_input_width_17_num_3_ready(PE_inst0_PE_input_width_17_num_3_ready),
		.PE_input_width_17_num_3_valid(CB_PE_input_width_17_num_3_valid_out),
		.PE_input_width_1_num_0(CB_PE_input_width_1_num_0_O),
		.PE_input_width_1_num_0_ready(PE_inst0_PE_input_width_1_num_0_ready),
		.PE_input_width_1_num_0_valid(CB_PE_input_width_1_num_0_valid_out),
		.PE_input_width_1_num_1(CB_PE_input_width_1_num_1_O),
		.PE_input_width_1_num_1_ready(PE_inst0_PE_input_width_1_num_1_ready),
		.PE_input_width_1_num_1_valid(CB_PE_input_width_1_num_1_valid_out),
		.PE_input_width_1_num_2(CB_PE_input_width_1_num_2_O),
		.PE_input_width_1_num_2_ready(PE_inst0_PE_input_width_1_num_2_ready),
		.PE_input_width_1_num_2_valid(CB_PE_input_width_1_num_2_valid_out),
		.PE_output_width_17_num_0(PE_inst0_PE_output_width_17_num_0),
		.PE_output_width_17_num_0_ready(SB_ID0_5TRACKS_B17_PE_PE_output_width_17_num_0_ready_out),
		.PE_output_width_17_num_0_valid(PE_inst0_PE_output_width_17_num_0_valid),
		.PE_output_width_17_num_1(PE_inst0_PE_output_width_17_num_1),
		.PE_output_width_17_num_1_ready(SB_ID0_5TRACKS_B17_PE_PE_output_width_17_num_1_ready_out),
		.PE_output_width_17_num_1_valid(PE_inst0_PE_output_width_17_num_1_valid),
		.PE_output_width_17_num_2(PE_inst0_PE_output_width_17_num_2),
		.PE_output_width_17_num_2_ready(SB_ID0_5TRACKS_B17_PE_PE_output_width_17_num_2_ready_out),
		.PE_output_width_17_num_2_valid(PE_inst0_PE_output_width_17_num_2_valid),
		.PE_output_width_1_num_0(PE_inst0_PE_output_width_1_num_0),
		.PE_output_width_1_num_0_ready(SB_ID0_5TRACKS_B1_PE_PE_output_width_1_num_0_ready_out),
		.PE_output_width_1_num_0_valid(PE_inst0_PE_output_width_1_num_0_valid),
		.clk(clk),
		.config_config_addr(self_config_config_addr_out[31:24]),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_0_out),
		.flush(CB_flush_O),
		.flush_core(flush),
		.read_config_data(PE_inst0_read_config_data),
		.reset(reset),
		.stall(stall)
	);
	ReadyValidLoopBack PE_output_width_17_num_0_loopback(
		.valid_out(PE_output_width_17_num_0_loopback_valid_out),
		.ready_in(SB_ID0_5TRACKS_B17_PE_PE_output_width_17_num_0_ready_out),
		.valid_in(PE_inst0_PE_output_width_17_num_0_valid)
	);
	ReadyValidLoopBack PE_output_width_17_num_1_loopback(
		.valid_out(PE_output_width_17_num_1_loopback_valid_out),
		.ready_in(SB_ID0_5TRACKS_B17_PE_PE_output_width_17_num_1_ready_out),
		.valid_in(PE_inst0_PE_output_width_17_num_1_valid)
	);
	ReadyValidLoopBack PE_output_width_17_num_2_loopback(
		.valid_out(PE_output_width_17_num_2_loopback_valid_out),
		.ready_in(SB_ID0_5TRACKS_B17_PE_PE_output_width_17_num_2_ready_out),
		.valid_in(PE_inst0_PE_output_width_17_num_2_valid)
	);
	ReadyValidLoopBack PE_output_width_1_num_0_loopback(
		.valid_out(PE_output_width_1_num_0_loopback_valid_out),
		.ready_in(SB_ID0_5TRACKS_B1_PE_PE_output_width_1_num_0_ready_out),
		.valid_in(PE_inst0_PE_output_width_1_num_0_valid)
	);
	PondCore PondCore_inst0(
		.PondTop_input_width_17_num_0(CB_PondTop_input_width_17_num_0_O),
		.PondTop_input_width_17_num_0_ready(PondCore_inst0_PondTop_input_width_17_num_0_ready),
		.PondTop_input_width_17_num_0_valid(CB_PondTop_input_width_17_num_0_valid_out),
		.PondTop_input_width_17_num_1(CB_PondTop_input_width_17_num_1_O),
		.PondTop_input_width_17_num_1_ready(PondCore_inst0_PondTop_input_width_17_num_1_ready),
		.PondTop_input_width_17_num_1_valid(CB_PondTop_input_width_17_num_1_valid_out),
		.PondTop_output_width_17_num_0(PondCore_inst0_PondTop_output_width_17_num_0),
		.PondTop_output_width_17_num_0_ready(SB_ID0_5TRACKS_B17_PE_PondTop_output_width_17_num_0_ready_out),
		.PondTop_output_width_17_num_0_valid(PondCore_inst0_PondTop_output_width_17_num_0_valid),
		.PondTop_output_width_17_num_1(PondCore_inst0_PondTop_output_width_17_num_1),
		.PondTop_output_width_17_num_1_ready(SB_ID0_5TRACKS_B17_PE_PondTop_output_width_17_num_1_ready_out),
		.PondTop_output_width_17_num_1_valid(PondCore_inst0_PondTop_output_width_17_num_1_valid),
		.PondTop_output_width_1_num_0(PondCore_inst0_PondTop_output_width_1_num_0),
		.PondTop_output_width_1_num_0_ready(SB_ID0_5TRACKS_B1_PE_PondTop_output_width_1_num_0_ready_out),
		.PondTop_output_width_1_num_0_valid(PondCore_inst0_PondTop_output_width_1_num_0_valid),
		.PondTop_output_width_1_num_1(PondCore_inst0_PondTop_output_width_1_num_1),
		.PondTop_output_width_1_num_1_ready(SB_ID0_5TRACKS_B1_PE_PondTop_output_width_1_num_1_ready_out),
		.PondTop_output_width_1_num_1_valid(PondCore_inst0_PondTop_output_width_1_num_1_valid),
		.clk(clk),
		.config_1_config_addr(self_config_config_addr_out[31:24]),
		.config_1_config_data(config_config_data),
		.config_1_read(config_read),
		.config_1_write(FEATURE_AND_2_out),
		.config_config_addr(self_config_config_addr_out[31:24]),
		.config_config_data(config_config_data),
		.config_en_0(DECODE_FEATURE_2_O),
		.config_read(config_read),
		.config_write(FEATURE_AND_1_out),
		.flush(CB_flush_O),
		.flush_core(flush),
		.read_config_data(PondCore_inst0_read_config_data),
		.read_config_data_1(PondCore_inst0_read_config_data_1),
		.reset(reset),
		.stall(stall)
	);
	ReadyValidLoopBack PondTop_output_width_17_num_0_loopback(
		.valid_out(PondTop_output_width_17_num_0_loopback_valid_out),
		.ready_in(SB_ID0_5TRACKS_B17_PE_PondTop_output_width_17_num_0_ready_out),
		.valid_in(PondCore_inst0_PondTop_output_width_17_num_0_valid)
	);
	ReadyValidLoopBack PondTop_output_width_17_num_1_loopback(
		.valid_out(PondTop_output_width_17_num_1_loopback_valid_out),
		.ready_in(SB_ID0_5TRACKS_B17_PE_PondTop_output_width_17_num_1_ready_out),
		.valid_in(PondCore_inst0_PondTop_output_width_17_num_1_valid)
	);
	ReadyValidLoopBack PondTop_output_width_1_num_0_loopback(
		.valid_out(PondTop_output_width_1_num_0_loopback_valid_out),
		.ready_in(SB_ID0_5TRACKS_B1_PE_PondTop_output_width_1_num_0_ready_out),
		.valid_in(PondCore_inst0_PondTop_output_width_1_num_0_valid)
	);
	ReadyValidLoopBack PondTop_output_width_1_num_1_loopback(
		.valid_out(PondTop_output_width_1_num_1_loopback_valid_out),
		.ready_in(SB_ID0_5TRACKS_B1_PE_PondTop_output_width_1_num_1_ready_out),
		.valid_in(PondCore_inst0_PondTop_output_width_1_num_1_valid)
	);
	PowerDomainConfigReg PowerDomainConfigReg_inst0(
		.clk(clk),
		.config_config_addr(self_config_config_addr_out[31:24]),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_15_out),
		.ps_en_out(PowerDomainConfigReg_inst0_ps_en_out),
		.read_config_data(PowerDomainConfigReg_inst0_read_config_data),
		.reset(reset)
	);
	PowerDomainOR PowerDomainOR(
		.I0(read_data_mux_O),
		.I1(read_config_data_in),
		.O(PowerDomainOR_O),
		.I_not(PowerDomainConfigReg_inst0_ps_en_out)
	);
	SB_ID0_5TRACKS_B17_PE SB_ID0_5TRACKS_B17_PE(
		.PE_input_width_17_num_0_enable(CB_PE_input_width_17_num_0_enable),
		.PE_input_width_17_num_0_out_sel(CB_PE_input_width_17_num_0_out_sel),
		.PE_input_width_17_num_0_ready(CB_PE_input_width_17_num_0_ready_out),
		.PE_input_width_17_num_1_enable(CB_PE_input_width_17_num_1_enable),
		.PE_input_width_17_num_1_out_sel(CB_PE_input_width_17_num_1_out_sel),
		.PE_input_width_17_num_1_ready(CB_PE_input_width_17_num_1_ready_out),
		.PE_input_width_17_num_2_enable(CB_PE_input_width_17_num_2_enable),
		.PE_input_width_17_num_2_out_sel(CB_PE_input_width_17_num_2_out_sel),
		.PE_input_width_17_num_2_ready(CB_PE_input_width_17_num_2_ready_out),
		.PE_input_width_17_num_3_enable(CB_PE_input_width_17_num_3_enable),
		.PE_input_width_17_num_3_out_sel(CB_PE_input_width_17_num_3_out_sel),
		.PE_input_width_17_num_3_ready(CB_PE_input_width_17_num_3_ready_out),
		.PE_output_width_17_num_0(PE_inst0_PE_output_width_17_num_0),
		.PE_output_width_17_num_0_ready_out(SB_ID0_5TRACKS_B17_PE_PE_output_width_17_num_0_ready_out),
		.PE_output_width_17_num_0_valid(PE_output_width_17_num_0_loopback_valid_out[0]),
		.PE_output_width_17_num_1(PE_inst0_PE_output_width_17_num_1),
		.PE_output_width_17_num_1_ready_out(SB_ID0_5TRACKS_B17_PE_PE_output_width_17_num_1_ready_out),
		.PE_output_width_17_num_1_valid(PE_output_width_17_num_1_loopback_valid_out[0]),
		.PE_output_width_17_num_2(PE_inst0_PE_output_width_17_num_2),
		.PE_output_width_17_num_2_ready_out(SB_ID0_5TRACKS_B17_PE_PE_output_width_17_num_2_ready_out),
		.PE_output_width_17_num_2_valid(PE_output_width_17_num_2_loopback_valid_out[0]),
		.PondTop_input_width_17_num_0_enable(CB_PondTop_input_width_17_num_0_enable),
		.PondTop_input_width_17_num_0_out_sel(CB_PondTop_input_width_17_num_0_out_sel),
		.PondTop_input_width_17_num_0_ready(CB_PondTop_input_width_17_num_0_ready_out),
		.PondTop_input_width_17_num_1_enable(CB_PondTop_input_width_17_num_1_enable),
		.PondTop_input_width_17_num_1_out_sel(CB_PondTop_input_width_17_num_1_out_sel),
		.PondTop_input_width_17_num_1_ready(CB_PondTop_input_width_17_num_1_ready_out),
		.PondTop_output_width_17_num_0_ready_out(SB_ID0_5TRACKS_B17_PE_PondTop_output_width_17_num_0_ready_out),
		.PondTop_output_width_17_num_0_valid(PondTop_output_width_17_num_0_loopback_valid_out[0]),
		.PondTop_output_width_17_num_1(PondCore_inst0_PondTop_output_width_17_num_1),
		.PondTop_output_width_17_num_1_ready_out(SB_ID0_5TRACKS_B17_PE_PondTop_output_width_17_num_1_ready_out),
		.PondTop_output_width_17_num_1_valid(PondTop_output_width_17_num_1_loopback_valid_out[0]),
		.SB_T0_EAST_SB_IN_B17(SB_T0_EAST_SB_IN_B17),
		.SB_T0_EAST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T0_EAST_SB_IN_B17_enable),
		.SB_T0_EAST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T0_EAST_SB_IN_B17_ready_out),
		.SB_T0_EAST_SB_IN_B17_valid_in(SB_T0_EAST_SB_IN_B17_valid),
		.SB_T0_EAST_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_EAST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T0_EAST_SB_OUT_B17_enable),
		.SB_T0_EAST_SB_OUT_B17_ready_in(SB_T0_EAST_SB_OUT_B17_ready_and_Z),
		.SB_T0_EAST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T0_EAST_SB_OUT_B17_valid_out),
		.SB_T0_NORTH_SB_IN_B17(SB_T0_NORTH_SB_IN_B17),
		.SB_T0_NORTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T0_NORTH_SB_IN_B17_enable),
		.SB_T0_NORTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T0_NORTH_SB_IN_B17_ready_out),
		.SB_T0_NORTH_SB_IN_B17_valid_in(SB_T0_NORTH_SB_IN_B17_valid),
		.SB_T0_NORTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T0_NORTH_SB_OUT_B17_enable),
		.SB_T0_NORTH_SB_OUT_B17_ready_in(SB_T0_NORTH_SB_OUT_B17_ready_and_Z),
		.SB_T0_NORTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T0_NORTH_SB_OUT_B17_valid_out),
		.SB_T0_SOUTH_SB_IN_B17(SB_T0_SOUTH_SB_IN_B17),
		.SB_T0_SOUTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T0_SOUTH_SB_IN_B17_enable),
		.SB_T0_SOUTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T0_SOUTH_SB_IN_B17_ready_out),
		.SB_T0_SOUTH_SB_IN_B17_valid_in(SB_T0_SOUTH_SB_IN_B17_valid),
		.SB_T0_SOUTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T0_SOUTH_SB_OUT_B17_enable),
		.SB_T0_SOUTH_SB_OUT_B17_ready_in(SB_T0_SOUTH_SB_OUT_B17_ready_and_Z),
		.SB_T0_SOUTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T0_SOUTH_SB_OUT_B17_valid_out),
		.SB_T0_WEST_SB_IN_B17(SB_T0_WEST_SB_IN_B17),
		.SB_T0_WEST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T0_WEST_SB_IN_B17_enable),
		.SB_T0_WEST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T0_WEST_SB_IN_B17_ready_out),
		.SB_T0_WEST_SB_IN_B17_valid_in(SB_T0_WEST_SB_IN_B17_valid),
		.SB_T0_WEST_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_WEST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T0_WEST_SB_OUT_B17_enable),
		.SB_T0_WEST_SB_OUT_B17_ready_in(SB_T0_WEST_SB_OUT_B17_ready_and_Z),
		.SB_T0_WEST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T0_WEST_SB_OUT_B17_valid_out),
		.SB_T1_EAST_SB_IN_B17(SB_T1_EAST_SB_IN_B17),
		.SB_T1_EAST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T1_EAST_SB_IN_B17_enable),
		.SB_T1_EAST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T1_EAST_SB_IN_B17_ready_out),
		.SB_T1_EAST_SB_IN_B17_valid_in(SB_T1_EAST_SB_IN_B17_valid),
		.SB_T1_EAST_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_EAST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T1_EAST_SB_OUT_B17_enable),
		.SB_T1_EAST_SB_OUT_B17_ready_in(SB_T1_EAST_SB_OUT_B17_ready_and_Z),
		.SB_T1_EAST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T1_EAST_SB_OUT_B17_valid_out),
		.SB_T1_NORTH_SB_IN_B17(SB_T1_NORTH_SB_IN_B17),
		.SB_T1_NORTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T1_NORTH_SB_IN_B17_enable),
		.SB_T1_NORTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T1_NORTH_SB_IN_B17_ready_out),
		.SB_T1_NORTH_SB_IN_B17_valid_in(SB_T1_NORTH_SB_IN_B17_valid),
		.SB_T1_NORTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T1_NORTH_SB_OUT_B17_enable),
		.SB_T1_NORTH_SB_OUT_B17_ready_in(SB_T1_NORTH_SB_OUT_B17_ready_and_Z),
		.SB_T1_NORTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T1_NORTH_SB_OUT_B17_valid_out),
		.SB_T1_SOUTH_SB_IN_B17(SB_T1_SOUTH_SB_IN_B17),
		.SB_T1_SOUTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T1_SOUTH_SB_IN_B17_enable),
		.SB_T1_SOUTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T1_SOUTH_SB_IN_B17_ready_out),
		.SB_T1_SOUTH_SB_IN_B17_valid_in(SB_T1_SOUTH_SB_IN_B17_valid),
		.SB_T1_SOUTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T1_SOUTH_SB_OUT_B17_enable),
		.SB_T1_SOUTH_SB_OUT_B17_ready_in(SB_T1_SOUTH_SB_OUT_B17_ready_and_Z),
		.SB_T1_SOUTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T1_SOUTH_SB_OUT_B17_valid_out),
		.SB_T1_WEST_SB_IN_B17(SB_T1_WEST_SB_IN_B17),
		.SB_T1_WEST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T1_WEST_SB_IN_B17_enable),
		.SB_T1_WEST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T1_WEST_SB_IN_B17_ready_out),
		.SB_T1_WEST_SB_IN_B17_valid_in(SB_T1_WEST_SB_IN_B17_valid),
		.SB_T1_WEST_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_WEST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T1_WEST_SB_OUT_B17_enable),
		.SB_T1_WEST_SB_OUT_B17_ready_in(SB_T1_WEST_SB_OUT_B17_ready_and_Z),
		.SB_T1_WEST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T1_WEST_SB_OUT_B17_valid_out),
		.SB_T2_EAST_SB_IN_B17(SB_T2_EAST_SB_IN_B17),
		.SB_T2_EAST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T2_EAST_SB_IN_B17_enable),
		.SB_T2_EAST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T2_EAST_SB_IN_B17_ready_out),
		.SB_T2_EAST_SB_IN_B17_valid_in(SB_T2_EAST_SB_IN_B17_valid),
		.SB_T2_EAST_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_EAST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T2_EAST_SB_OUT_B17_enable),
		.SB_T2_EAST_SB_OUT_B17_ready_in(SB_T2_EAST_SB_OUT_B17_ready_and_Z),
		.SB_T2_EAST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T2_EAST_SB_OUT_B17_valid_out),
		.SB_T2_NORTH_SB_IN_B17(SB_T2_NORTH_SB_IN_B17),
		.SB_T2_NORTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T2_NORTH_SB_IN_B17_enable),
		.SB_T2_NORTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T2_NORTH_SB_IN_B17_ready_out),
		.SB_T2_NORTH_SB_IN_B17_valid_in(SB_T2_NORTH_SB_IN_B17_valid),
		.SB_T2_NORTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T2_NORTH_SB_OUT_B17_enable),
		.SB_T2_NORTH_SB_OUT_B17_ready_in(SB_T2_NORTH_SB_OUT_B17_ready_and_Z),
		.SB_T2_NORTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T2_NORTH_SB_OUT_B17_valid_out),
		.SB_T2_SOUTH_SB_IN_B17(SB_T2_SOUTH_SB_IN_B17),
		.SB_T2_SOUTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T2_SOUTH_SB_IN_B17_enable),
		.SB_T2_SOUTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T2_SOUTH_SB_IN_B17_ready_out),
		.SB_T2_SOUTH_SB_IN_B17_valid_in(SB_T2_SOUTH_SB_IN_B17_valid),
		.SB_T2_SOUTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T2_SOUTH_SB_OUT_B17_enable),
		.SB_T2_SOUTH_SB_OUT_B17_ready_in(SB_T2_SOUTH_SB_OUT_B17_ready_and_Z),
		.SB_T2_SOUTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T2_SOUTH_SB_OUT_B17_valid_out),
		.SB_T2_WEST_SB_IN_B17(SB_T2_WEST_SB_IN_B17),
		.SB_T2_WEST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T2_WEST_SB_IN_B17_enable),
		.SB_T2_WEST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T2_WEST_SB_IN_B17_ready_out),
		.SB_T2_WEST_SB_IN_B17_valid_in(SB_T2_WEST_SB_IN_B17_valid),
		.SB_T2_WEST_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_WEST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T2_WEST_SB_OUT_B17_enable),
		.SB_T2_WEST_SB_OUT_B17_ready_in(SB_T2_WEST_SB_OUT_B17_ready_and_Z),
		.SB_T2_WEST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T2_WEST_SB_OUT_B17_valid_out),
		.SB_T3_EAST_SB_IN_B17(SB_T3_EAST_SB_IN_B17),
		.SB_T3_EAST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T3_EAST_SB_IN_B17_enable),
		.SB_T3_EAST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T3_EAST_SB_IN_B17_ready_out),
		.SB_T3_EAST_SB_IN_B17_valid_in(SB_T3_EAST_SB_IN_B17_valid),
		.SB_T3_EAST_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_EAST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T3_EAST_SB_OUT_B17_enable),
		.SB_T3_EAST_SB_OUT_B17_ready_in(SB_T3_EAST_SB_OUT_B17_ready_and_Z),
		.SB_T3_EAST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T3_EAST_SB_OUT_B17_valid_out),
		.SB_T3_NORTH_SB_IN_B17(SB_T3_NORTH_SB_IN_B17),
		.SB_T3_NORTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T3_NORTH_SB_IN_B17_enable),
		.SB_T3_NORTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T3_NORTH_SB_IN_B17_ready_out),
		.SB_T3_NORTH_SB_IN_B17_valid_in(SB_T3_NORTH_SB_IN_B17_valid),
		.SB_T3_NORTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T3_NORTH_SB_OUT_B17_enable),
		.SB_T3_NORTH_SB_OUT_B17_ready_in(SB_T3_NORTH_SB_OUT_B17_ready_and_Z),
		.SB_T3_NORTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T3_NORTH_SB_OUT_B17_valid_out),
		.SB_T3_SOUTH_SB_IN_B17(SB_T3_SOUTH_SB_IN_B17),
		.SB_T3_SOUTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T3_SOUTH_SB_IN_B17_enable),
		.SB_T3_SOUTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T3_SOUTH_SB_IN_B17_ready_out),
		.SB_T3_SOUTH_SB_IN_B17_valid_in(SB_T3_SOUTH_SB_IN_B17_valid),
		.SB_T3_SOUTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T3_SOUTH_SB_OUT_B17_enable),
		.SB_T3_SOUTH_SB_OUT_B17_ready_in(SB_T3_SOUTH_SB_OUT_B17_ready_and_Z),
		.SB_T3_SOUTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T3_SOUTH_SB_OUT_B17_valid_out),
		.SB_T3_WEST_SB_IN_B17(SB_T3_WEST_SB_IN_B17),
		.SB_T3_WEST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T3_WEST_SB_IN_B17_enable),
		.SB_T3_WEST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T3_WEST_SB_IN_B17_ready_out),
		.SB_T3_WEST_SB_IN_B17_valid_in(SB_T3_WEST_SB_IN_B17_valid),
		.SB_T3_WEST_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_WEST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T3_WEST_SB_OUT_B17_enable),
		.SB_T3_WEST_SB_OUT_B17_ready_in(SB_T3_WEST_SB_OUT_B17_ready_and_Z),
		.SB_T3_WEST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T3_WEST_SB_OUT_B17_valid_out),
		.SB_T4_EAST_SB_IN_B17(SB_T4_EAST_SB_IN_B17),
		.SB_T4_EAST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T4_EAST_SB_IN_B17_enable),
		.SB_T4_EAST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T4_EAST_SB_IN_B17_ready_out),
		.SB_T4_EAST_SB_IN_B17_valid_in(SB_T4_EAST_SB_IN_B17_valid),
		.SB_T4_EAST_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_EAST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T4_EAST_SB_OUT_B17_enable),
		.SB_T4_EAST_SB_OUT_B17_ready_in(SB_T4_EAST_SB_OUT_B17_ready_and_Z),
		.SB_T4_EAST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T4_EAST_SB_OUT_B17_valid_out),
		.SB_T4_NORTH_SB_IN_B17(SB_T4_NORTH_SB_IN_B17),
		.SB_T4_NORTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T4_NORTH_SB_IN_B17_enable),
		.SB_T4_NORTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T4_NORTH_SB_IN_B17_ready_out),
		.SB_T4_NORTH_SB_IN_B17_valid_in(SB_T4_NORTH_SB_IN_B17_valid),
		.SB_T4_NORTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T4_NORTH_SB_OUT_B17_enable),
		.SB_T4_NORTH_SB_OUT_B17_ready_in(SB_T4_NORTH_SB_OUT_B17_ready_and_Z),
		.SB_T4_NORTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T4_NORTH_SB_OUT_B17_valid_out),
		.SB_T4_SOUTH_SB_IN_B17(SB_T4_SOUTH_SB_IN_B17),
		.SB_T4_SOUTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T4_SOUTH_SB_IN_B17_enable),
		.SB_T4_SOUTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T4_SOUTH_SB_IN_B17_ready_out),
		.SB_T4_SOUTH_SB_IN_B17_valid_in(SB_T4_SOUTH_SB_IN_B17_valid),
		.SB_T4_SOUTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T4_SOUTH_SB_OUT_B17_enable),
		.SB_T4_SOUTH_SB_OUT_B17_ready_in(SB_T4_SOUTH_SB_OUT_B17_ready_and_Z),
		.SB_T4_SOUTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T4_SOUTH_SB_OUT_B17_valid_out),
		.SB_T4_WEST_SB_IN_B17(SB_T4_WEST_SB_IN_B17),
		.SB_T4_WEST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T4_WEST_SB_IN_B17_enable),
		.SB_T4_WEST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T4_WEST_SB_IN_B17_ready_out),
		.SB_T4_WEST_SB_IN_B17_valid_in(SB_T4_WEST_SB_IN_B17_valid),
		.SB_T4_WEST_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_WEST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T4_WEST_SB_OUT_B17_enable),
		.SB_T4_WEST_SB_OUT_B17_ready_in(SB_T4_WEST_SB_OUT_B17_ready_and_Z),
		.SB_T4_WEST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T4_WEST_SB_OUT_B17_valid_out),
		.clk(clk),
		.config_config_addr(self_config_config_addr_out[31:24]),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_14_out),
		.read_config_data(SB_ID0_5TRACKS_B17_PE_read_config_data),
		.reset(reset),
		.stall(stall)
	);
	SB_ID0_5TRACKS_B1_PE SB_ID0_5TRACKS_B1_PE(
		.PE_input_width_1_num_0_enable(CB_PE_input_width_1_num_0_enable),
		.PE_input_width_1_num_0_out_sel(CB_PE_input_width_1_num_0_out_sel),
		.PE_input_width_1_num_0_ready(CB_PE_input_width_1_num_0_ready_out),
		.PE_input_width_1_num_1_enable(CB_PE_input_width_1_num_1_enable),
		.PE_input_width_1_num_1_out_sel(CB_PE_input_width_1_num_1_out_sel),
		.PE_input_width_1_num_1_ready(CB_PE_input_width_1_num_1_ready_out),
		.PE_input_width_1_num_2_enable(CB_PE_input_width_1_num_2_enable),
		.PE_input_width_1_num_2_out_sel(CB_PE_input_width_1_num_2_out_sel),
		.PE_input_width_1_num_2_ready(CB_PE_input_width_1_num_2_ready_out),
		.PE_output_width_1_num_0(PE_inst0_PE_output_width_1_num_0),
		.PE_output_width_1_num_0_ready_out(SB_ID0_5TRACKS_B1_PE_PE_output_width_1_num_0_ready_out),
		.PE_output_width_1_num_0_valid(PE_output_width_1_num_0_loopback_valid_out[0]),
		.PondTop_output_width_1_num_0(PondCore_inst0_PondTop_output_width_1_num_0),
		.PondTop_output_width_1_num_0_ready_out(SB_ID0_5TRACKS_B1_PE_PondTop_output_width_1_num_0_ready_out),
		.PondTop_output_width_1_num_0_valid(PondTop_output_width_1_num_0_loopback_valid_out[0]),
		.PondTop_output_width_1_num_1(PondCore_inst0_PondTop_output_width_1_num_1),
		.PondTop_output_width_1_num_1_ready_out(SB_ID0_5TRACKS_B1_PE_PondTop_output_width_1_num_1_ready_out),
		.PondTop_output_width_1_num_1_valid(PondTop_output_width_1_num_1_loopback_valid_out[0]),
		.SB_T0_EAST_SB_IN_B1(SB_T0_EAST_SB_IN_B1),
		.SB_T0_EAST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_IN_B1_enable),
		.SB_T0_EAST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_IN_B1_ready_out),
		.SB_T0_EAST_SB_IN_B1_valid_in(SB_T0_EAST_SB_IN_B1_valid),
		.SB_T0_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_EAST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_OUT_B1_enable),
		.SB_T0_EAST_SB_OUT_B1_ready_in(SB_T0_EAST_SB_OUT_B1_ready_and_Z),
		.SB_T0_EAST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_OUT_B1_valid_out),
		.SB_T0_NORTH_SB_IN_B1(SB_T0_NORTH_SB_IN_B1),
		.SB_T0_NORTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_IN_B1_enable),
		.SB_T0_NORTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_IN_B1_ready_out),
		.SB_T0_NORTH_SB_IN_B1_valid_in(SB_T0_NORTH_SB_IN_B1_valid),
		.SB_T0_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_OUT_B1_enable),
		.SB_T0_NORTH_SB_OUT_B1_ready_in(SB_T0_NORTH_SB_OUT_B1_ready_and_Z),
		.SB_T0_NORTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_OUT_B1_valid_out),
		.SB_T0_SOUTH_SB_IN_B1(SB_T0_SOUTH_SB_IN_B1),
		.SB_T0_SOUTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_IN_B1_enable),
		.SB_T0_SOUTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_IN_B1_ready_out),
		.SB_T0_SOUTH_SB_IN_B1_valid_in(SB_T0_SOUTH_SB_IN_B1_valid),
		.SB_T0_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_OUT_B1_enable),
		.SB_T0_SOUTH_SB_OUT_B1_ready_in(SB_T0_SOUTH_SB_OUT_B1_ready_and_Z),
		.SB_T0_SOUTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_OUT_B1_valid_out),
		.SB_T0_WEST_SB_IN_B1(SB_T0_WEST_SB_IN_B1),
		.SB_T0_WEST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_IN_B1_enable),
		.SB_T0_WEST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_IN_B1_ready_out),
		.SB_T0_WEST_SB_IN_B1_valid_in(SB_T0_WEST_SB_IN_B1_valid),
		.SB_T0_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_WEST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_OUT_B1_enable),
		.SB_T0_WEST_SB_OUT_B1_ready_in(SB_T0_WEST_SB_OUT_B1_ready_and_Z),
		.SB_T0_WEST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_OUT_B1_valid_out),
		.SB_T1_EAST_SB_IN_B1(SB_T1_EAST_SB_IN_B1),
		.SB_T1_EAST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_IN_B1_enable),
		.SB_T1_EAST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_IN_B1_ready_out),
		.SB_T1_EAST_SB_IN_B1_valid_in(SB_T1_EAST_SB_IN_B1_valid),
		.SB_T1_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_EAST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_OUT_B1_enable),
		.SB_T1_EAST_SB_OUT_B1_ready_in(SB_T1_EAST_SB_OUT_B1_ready_and_Z),
		.SB_T1_EAST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_OUT_B1_valid_out),
		.SB_T1_NORTH_SB_IN_B1(SB_T1_NORTH_SB_IN_B1),
		.SB_T1_NORTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_IN_B1_enable),
		.SB_T1_NORTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_IN_B1_ready_out),
		.SB_T1_NORTH_SB_IN_B1_valid_in(SB_T1_NORTH_SB_IN_B1_valid),
		.SB_T1_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_OUT_B1_enable),
		.SB_T1_NORTH_SB_OUT_B1_ready_in(SB_T1_NORTH_SB_OUT_B1_ready_and_Z),
		.SB_T1_NORTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_OUT_B1_valid_out),
		.SB_T1_SOUTH_SB_IN_B1(SB_T1_SOUTH_SB_IN_B1),
		.SB_T1_SOUTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_IN_B1_enable),
		.SB_T1_SOUTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_IN_B1_ready_out),
		.SB_T1_SOUTH_SB_IN_B1_valid_in(SB_T1_SOUTH_SB_IN_B1_valid),
		.SB_T1_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_OUT_B1_enable),
		.SB_T1_SOUTH_SB_OUT_B1_ready_in(SB_T1_SOUTH_SB_OUT_B1_ready_and_Z),
		.SB_T1_SOUTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_OUT_B1_valid_out),
		.SB_T1_WEST_SB_IN_B1(SB_T1_WEST_SB_IN_B1),
		.SB_T1_WEST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_IN_B1_enable),
		.SB_T1_WEST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_IN_B1_ready_out),
		.SB_T1_WEST_SB_IN_B1_valid_in(SB_T1_WEST_SB_IN_B1_valid),
		.SB_T1_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_WEST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_OUT_B1_enable),
		.SB_T1_WEST_SB_OUT_B1_ready_in(SB_T1_WEST_SB_OUT_B1_ready_and_Z),
		.SB_T1_WEST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_OUT_B1_valid_out),
		.SB_T2_EAST_SB_IN_B1(SB_T2_EAST_SB_IN_B1),
		.SB_T2_EAST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_IN_B1_enable),
		.SB_T2_EAST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_IN_B1_ready_out),
		.SB_T2_EAST_SB_IN_B1_valid_in(SB_T2_EAST_SB_IN_B1_valid),
		.SB_T2_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_EAST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_OUT_B1_enable),
		.SB_T2_EAST_SB_OUT_B1_ready_in(SB_T2_EAST_SB_OUT_B1_ready_and_Z),
		.SB_T2_EAST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_OUT_B1_valid_out),
		.SB_T2_NORTH_SB_IN_B1(SB_T2_NORTH_SB_IN_B1),
		.SB_T2_NORTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_IN_B1_enable),
		.SB_T2_NORTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_IN_B1_ready_out),
		.SB_T2_NORTH_SB_IN_B1_valid_in(SB_T2_NORTH_SB_IN_B1_valid),
		.SB_T2_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_OUT_B1_enable),
		.SB_T2_NORTH_SB_OUT_B1_ready_in(SB_T2_NORTH_SB_OUT_B1_ready_and_Z),
		.SB_T2_NORTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_OUT_B1_valid_out),
		.SB_T2_SOUTH_SB_IN_B1(SB_T2_SOUTH_SB_IN_B1),
		.SB_T2_SOUTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_IN_B1_enable),
		.SB_T2_SOUTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_IN_B1_ready_out),
		.SB_T2_SOUTH_SB_IN_B1_valid_in(SB_T2_SOUTH_SB_IN_B1_valid),
		.SB_T2_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_OUT_B1_enable),
		.SB_T2_SOUTH_SB_OUT_B1_ready_in(SB_T2_SOUTH_SB_OUT_B1_ready_and_Z),
		.SB_T2_SOUTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_OUT_B1_valid_out),
		.SB_T2_WEST_SB_IN_B1(SB_T2_WEST_SB_IN_B1),
		.SB_T2_WEST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_IN_B1_enable),
		.SB_T2_WEST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_IN_B1_ready_out),
		.SB_T2_WEST_SB_IN_B1_valid_in(SB_T2_WEST_SB_IN_B1_valid),
		.SB_T2_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_WEST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_OUT_B1_enable),
		.SB_T2_WEST_SB_OUT_B1_ready_in(SB_T2_WEST_SB_OUT_B1_ready_and_Z),
		.SB_T2_WEST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_OUT_B1_valid_out),
		.SB_T3_EAST_SB_IN_B1(SB_T3_EAST_SB_IN_B1),
		.SB_T3_EAST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_IN_B1_enable),
		.SB_T3_EAST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_IN_B1_ready_out),
		.SB_T3_EAST_SB_IN_B1_valid_in(SB_T3_EAST_SB_IN_B1_valid),
		.SB_T3_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_EAST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_OUT_B1_enable),
		.SB_T3_EAST_SB_OUT_B1_ready_in(SB_T3_EAST_SB_OUT_B1_ready_and_Z),
		.SB_T3_EAST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_OUT_B1_valid_out),
		.SB_T3_NORTH_SB_IN_B1(SB_T3_NORTH_SB_IN_B1),
		.SB_T3_NORTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_IN_B1_enable),
		.SB_T3_NORTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_IN_B1_ready_out),
		.SB_T3_NORTH_SB_IN_B1_valid_in(SB_T3_NORTH_SB_IN_B1_valid),
		.SB_T3_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_OUT_B1_enable),
		.SB_T3_NORTH_SB_OUT_B1_ready_in(SB_T3_NORTH_SB_OUT_B1_ready_and_Z),
		.SB_T3_NORTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_OUT_B1_valid_out),
		.SB_T3_SOUTH_SB_IN_B1(SB_T3_SOUTH_SB_IN_B1),
		.SB_T3_SOUTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_IN_B1_enable),
		.SB_T3_SOUTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_IN_B1_ready_out),
		.SB_T3_SOUTH_SB_IN_B1_valid_in(SB_T3_SOUTH_SB_IN_B1_valid),
		.SB_T3_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_OUT_B1_enable),
		.SB_T3_SOUTH_SB_OUT_B1_ready_in(SB_T3_SOUTH_SB_OUT_B1_ready_and_Z),
		.SB_T3_SOUTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_OUT_B1_valid_out),
		.SB_T3_WEST_SB_IN_B1(SB_T3_WEST_SB_IN_B1),
		.SB_T3_WEST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_IN_B1_enable),
		.SB_T3_WEST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_IN_B1_ready_out),
		.SB_T3_WEST_SB_IN_B1_valid_in(SB_T3_WEST_SB_IN_B1_valid),
		.SB_T3_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_WEST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_OUT_B1_enable),
		.SB_T3_WEST_SB_OUT_B1_ready_in(SB_T3_WEST_SB_OUT_B1_ready_and_Z),
		.SB_T3_WEST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_OUT_B1_valid_out),
		.SB_T4_EAST_SB_IN_B1(SB_T4_EAST_SB_IN_B1),
		.SB_T4_EAST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_IN_B1_enable),
		.SB_T4_EAST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_IN_B1_ready_out),
		.SB_T4_EAST_SB_IN_B1_valid_in(SB_T4_EAST_SB_IN_B1_valid),
		.SB_T4_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_EAST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_OUT_B1_enable),
		.SB_T4_EAST_SB_OUT_B1_ready_in(SB_T4_EAST_SB_OUT_B1_ready_and_Z),
		.SB_T4_EAST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_OUT_B1_valid_out),
		.SB_T4_NORTH_SB_IN_B1(SB_T4_NORTH_SB_IN_B1),
		.SB_T4_NORTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_IN_B1_enable),
		.SB_T4_NORTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_IN_B1_ready_out),
		.SB_T4_NORTH_SB_IN_B1_valid_in(SB_T4_NORTH_SB_IN_B1_valid),
		.SB_T4_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_OUT_B1_enable),
		.SB_T4_NORTH_SB_OUT_B1_ready_in(SB_T4_NORTH_SB_OUT_B1_ready_and_Z),
		.SB_T4_NORTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_OUT_B1_valid_out),
		.SB_T4_SOUTH_SB_IN_B1(SB_T4_SOUTH_SB_IN_B1),
		.SB_T4_SOUTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_IN_B1_enable),
		.SB_T4_SOUTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_IN_B1_ready_out),
		.SB_T4_SOUTH_SB_IN_B1_valid_in(SB_T4_SOUTH_SB_IN_B1_valid),
		.SB_T4_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_OUT_B1_enable),
		.SB_T4_SOUTH_SB_OUT_B1_ready_in(SB_T4_SOUTH_SB_OUT_B1_ready_and_Z),
		.SB_T4_SOUTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_OUT_B1_valid_out),
		.SB_T4_WEST_SB_IN_B1(SB_T4_WEST_SB_IN_B1),
		.SB_T4_WEST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_IN_B1_enable),
		.SB_T4_WEST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_IN_B1_ready_out),
		.SB_T4_WEST_SB_IN_B1_valid_in(SB_T4_WEST_SB_IN_B1_valid),
		.SB_T4_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_WEST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_OUT_B1_enable),
		.SB_T4_WEST_SB_OUT_B1_ready_in(SB_T4_WEST_SB_OUT_B1_ready_and_Z),
		.SB_T4_WEST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_OUT_B1_valid_out),
		.clk(clk),
		.config_config_addr(self_config_config_addr_out[31:24]),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_13_out),
		.read_config_data(SB_ID0_5TRACKS_B1_PE_read_config_data),
		.reset(reset),
		.stall(stall)
	);
	and_cell SB_T0_EAST_SB_OUT_B17_ready_and(
		.A(SB_T0_EAST_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_PE_SB_T0_EAST_SB_OUT_B17_enable),
		.Z(SB_T0_EAST_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T0_EAST_SB_OUT_B1_ready_and(
		.A(SB_T0_EAST_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_OUT_B1_enable),
		.Z(SB_T0_EAST_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T0_NORTH_SB_OUT_B17_ready_and(
		.A(SB_T0_NORTH_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_PE_SB_T0_NORTH_SB_OUT_B17_enable),
		.Z(SB_T0_NORTH_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T0_NORTH_SB_OUT_B1_ready_and(
		.A(SB_T0_NORTH_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_OUT_B1_enable),
		.Z(SB_T0_NORTH_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T0_SOUTH_SB_OUT_B17_ready_and(
		.A(SB_T0_SOUTH_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_PE_SB_T0_SOUTH_SB_OUT_B17_enable),
		.Z(SB_T0_SOUTH_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T0_SOUTH_SB_OUT_B1_ready_and(
		.A(SB_T0_SOUTH_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_OUT_B1_enable),
		.Z(SB_T0_SOUTH_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T0_WEST_SB_OUT_B17_ready_and(
		.A(SB_T0_WEST_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_PE_SB_T0_WEST_SB_OUT_B17_enable),
		.Z(SB_T0_WEST_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T0_WEST_SB_OUT_B1_ready_and(
		.A(SB_T0_WEST_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_OUT_B1_enable),
		.Z(SB_T0_WEST_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T1_EAST_SB_OUT_B17_ready_and(
		.A(SB_T1_EAST_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_PE_SB_T1_EAST_SB_OUT_B17_enable),
		.Z(SB_T1_EAST_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T1_EAST_SB_OUT_B1_ready_and(
		.A(SB_T1_EAST_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_OUT_B1_enable),
		.Z(SB_T1_EAST_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T1_NORTH_SB_OUT_B17_ready_and(
		.A(SB_T1_NORTH_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_PE_SB_T1_NORTH_SB_OUT_B17_enable),
		.Z(SB_T1_NORTH_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T1_NORTH_SB_OUT_B1_ready_and(
		.A(SB_T1_NORTH_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_OUT_B1_enable),
		.Z(SB_T1_NORTH_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T1_SOUTH_SB_OUT_B17_ready_and(
		.A(SB_T1_SOUTH_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_PE_SB_T1_SOUTH_SB_OUT_B17_enable),
		.Z(SB_T1_SOUTH_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T1_SOUTH_SB_OUT_B1_ready_and(
		.A(SB_T1_SOUTH_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_OUT_B1_enable),
		.Z(SB_T1_SOUTH_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T1_WEST_SB_OUT_B17_ready_and(
		.A(SB_T1_WEST_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_PE_SB_T1_WEST_SB_OUT_B17_enable),
		.Z(SB_T1_WEST_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T1_WEST_SB_OUT_B1_ready_and(
		.A(SB_T1_WEST_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_OUT_B1_enable),
		.Z(SB_T1_WEST_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T2_EAST_SB_OUT_B17_ready_and(
		.A(SB_T2_EAST_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_PE_SB_T2_EAST_SB_OUT_B17_enable),
		.Z(SB_T2_EAST_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T2_EAST_SB_OUT_B1_ready_and(
		.A(SB_T2_EAST_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_OUT_B1_enable),
		.Z(SB_T2_EAST_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T2_NORTH_SB_OUT_B17_ready_and(
		.A(SB_T2_NORTH_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_PE_SB_T2_NORTH_SB_OUT_B17_enable),
		.Z(SB_T2_NORTH_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T2_NORTH_SB_OUT_B1_ready_and(
		.A(SB_T2_NORTH_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_OUT_B1_enable),
		.Z(SB_T2_NORTH_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T2_SOUTH_SB_OUT_B17_ready_and(
		.A(SB_T2_SOUTH_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_PE_SB_T2_SOUTH_SB_OUT_B17_enable),
		.Z(SB_T2_SOUTH_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T2_SOUTH_SB_OUT_B1_ready_and(
		.A(SB_T2_SOUTH_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_OUT_B1_enable),
		.Z(SB_T2_SOUTH_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T2_WEST_SB_OUT_B17_ready_and(
		.A(SB_T2_WEST_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_PE_SB_T2_WEST_SB_OUT_B17_enable),
		.Z(SB_T2_WEST_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T2_WEST_SB_OUT_B1_ready_and(
		.A(SB_T2_WEST_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_OUT_B1_enable),
		.Z(SB_T2_WEST_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T3_EAST_SB_OUT_B17_ready_and(
		.A(SB_T3_EAST_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_PE_SB_T3_EAST_SB_OUT_B17_enable),
		.Z(SB_T3_EAST_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T3_EAST_SB_OUT_B1_ready_and(
		.A(SB_T3_EAST_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_OUT_B1_enable),
		.Z(SB_T3_EAST_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T3_NORTH_SB_OUT_B17_ready_and(
		.A(SB_T3_NORTH_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_PE_SB_T3_NORTH_SB_OUT_B17_enable),
		.Z(SB_T3_NORTH_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T3_NORTH_SB_OUT_B1_ready_and(
		.A(SB_T3_NORTH_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_OUT_B1_enable),
		.Z(SB_T3_NORTH_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T3_SOUTH_SB_OUT_B17_ready_and(
		.A(SB_T3_SOUTH_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_PE_SB_T3_SOUTH_SB_OUT_B17_enable),
		.Z(SB_T3_SOUTH_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T3_SOUTH_SB_OUT_B1_ready_and(
		.A(SB_T3_SOUTH_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_OUT_B1_enable),
		.Z(SB_T3_SOUTH_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T3_WEST_SB_OUT_B17_ready_and(
		.A(SB_T3_WEST_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_PE_SB_T3_WEST_SB_OUT_B17_enable),
		.Z(SB_T3_WEST_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T3_WEST_SB_OUT_B1_ready_and(
		.A(SB_T3_WEST_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_OUT_B1_enable),
		.Z(SB_T3_WEST_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T4_EAST_SB_OUT_B17_ready_and(
		.A(SB_T4_EAST_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_PE_SB_T4_EAST_SB_OUT_B17_enable),
		.Z(SB_T4_EAST_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T4_EAST_SB_OUT_B1_ready_and(
		.A(SB_T4_EAST_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_OUT_B1_enable),
		.Z(SB_T4_EAST_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T4_NORTH_SB_OUT_B17_ready_and(
		.A(SB_T4_NORTH_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_PE_SB_T4_NORTH_SB_OUT_B17_enable),
		.Z(SB_T4_NORTH_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T4_NORTH_SB_OUT_B1_ready_and(
		.A(SB_T4_NORTH_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_OUT_B1_enable),
		.Z(SB_T4_NORTH_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T4_SOUTH_SB_OUT_B17_ready_and(
		.A(SB_T4_SOUTH_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_PE_SB_T4_SOUTH_SB_OUT_B17_enable),
		.Z(SB_T4_SOUTH_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T4_SOUTH_SB_OUT_B1_ready_and(
		.A(SB_T4_SOUTH_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_OUT_B1_enable),
		.Z(SB_T4_SOUTH_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T4_WEST_SB_OUT_B17_ready_and(
		.A(SB_T4_WEST_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_PE_SB_T4_WEST_SB_OUT_B17_enable),
		.Z(SB_T4_WEST_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T4_WEST_SB_OUT_B1_ready_and(
		.A(SB_T4_WEST_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_OUT_B1_enable),
		.Z(SB_T4_WEST_SB_OUT_B1_ready_and_Z)
	);
	corebit_and and_inst0(
		.in0(coreir_eq_16_inst0_out),
		.in1(config_read[0]),
		.out(and_inst0_out)
	);
	corebit_and and_inst1(
		.in0(coreir_eq_16_inst0_out),
		.in1(config_write[0]),
		.out(and_inst1_out)
	);
	corebit_const #(.value(1'b1)) bit_const_1_None(.out(bit_const_1_None_out));
	coreir_const #(
		.value(8'h00),
		.width(8)
	) const_0_8(.out(const_0_8_out));
	coreir_const #(
		.value(9'h1ff),
		.width(9)
	) const_511_9(.out(const_511_9_out));
	coreir_eq #(.width(16)) coreir_eq_16_inst0(
		.in0(tile_id),
		.in1(self_config_config_addr_out[15:0]),
		.out(coreir_eq_16_inst0_out)
	);
	coreir_wrap coreir_wrapOutClock_inst0(
		.in(clk_pass_through),
		.out(coreir_wrapOutClock_inst0_out)
	);
	coreir_wrap coreir_wrapOutClock_inst1(
		.in(clk_pass_through),
		.out(coreir_wrapOutClock_inst1_out)
	);
	wire [511:0] read_data_mux_I;
	assign read_data_mux_I[480+:32] = PowerDomainConfigReg_inst0_read_config_data;
	assign read_data_mux_I[448+:32] = SB_ID0_5TRACKS_B17_PE_read_config_data;
	assign read_data_mux_I[416+:32] = SB_ID0_5TRACKS_B1_PE_read_config_data;
	assign read_data_mux_I[384+:32] = CB_flush_read_config_data;
	assign read_data_mux_I[352+:32] = CB_PondTop_input_width_17_num_1_read_config_data;
	assign read_data_mux_I[320+:32] = CB_PondTop_input_width_17_num_0_read_config_data;
	assign read_data_mux_I[288+:32] = CB_PE_input_width_1_num_2_read_config_data;
	assign read_data_mux_I[256+:32] = CB_PE_input_width_1_num_1_read_config_data;
	assign read_data_mux_I[224+:32] = CB_PE_input_width_1_num_0_read_config_data;
	assign read_data_mux_I[192+:32] = CB_PE_input_width_17_num_3_read_config_data;
	assign read_data_mux_I[160+:32] = CB_PE_input_width_17_num_2_read_config_data;
	assign read_data_mux_I[128+:32] = CB_PE_input_width_17_num_1_read_config_data;
	assign read_data_mux_I[96+:32] = CB_PE_input_width_17_num_0_read_config_data;
	assign read_data_mux_I[64+:32] = PondCore_inst0_read_config_data_1;
	assign read_data_mux_I[32+:32] = PondCore_inst0_read_config_data;
	assign read_data_mux_I[0+:32] = PE_inst0_read_config_data;
	MuxWithDefaultWrapper_16_32_8_0 read_data_mux(
		.I(read_data_mux_I),
		.S(self_config_config_addr_out[23:16]),
		.EN(and_inst0_out),
		.O(read_data_mux_O)
	);
	mantle_wire__typeBit32 self_config_config_addr(
		.in(config_config_addr),
		.out(self_config_config_addr_out)
	);
	assign SB_T0_EAST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T0_EAST_SB_IN_B17_ready_out;
	assign SB_T0_EAST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_IN_B1_ready_out;
	assign SB_T0_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_OUT_B1;
	assign SB_T0_EAST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T0_EAST_SB_OUT_B17;
	assign SB_T0_EAST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T0_EAST_SB_OUT_B17_valid_out;
	assign SB_T0_EAST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_OUT_B1_valid_out;
	assign SB_T0_NORTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T0_NORTH_SB_IN_B17_ready_out;
	assign SB_T0_NORTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_IN_B1_ready_out;
	assign SB_T0_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_OUT_B1;
	assign SB_T0_NORTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T0_NORTH_SB_OUT_B17;
	assign SB_T0_NORTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T0_NORTH_SB_OUT_B17_valid_out;
	assign SB_T0_NORTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_OUT_B1_valid_out;
	assign SB_T0_SOUTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T0_SOUTH_SB_IN_B17_ready_out;
	assign SB_T0_SOUTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_IN_B1_ready_out;
	assign SB_T0_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_OUT_B1;
	assign SB_T0_SOUTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T0_SOUTH_SB_OUT_B17;
	assign SB_T0_SOUTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T0_SOUTH_SB_OUT_B17_valid_out;
	assign SB_T0_SOUTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_OUT_B1_valid_out;
	assign SB_T0_WEST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T0_WEST_SB_IN_B17_ready_out;
	assign SB_T0_WEST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_IN_B1_ready_out;
	assign SB_T0_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_OUT_B1;
	assign SB_T0_WEST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T0_WEST_SB_OUT_B17;
	assign SB_T0_WEST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T0_WEST_SB_OUT_B17_valid_out;
	assign SB_T0_WEST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_OUT_B1_valid_out;
	assign SB_T1_EAST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T1_EAST_SB_IN_B17_ready_out;
	assign SB_T1_EAST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_IN_B1_ready_out;
	assign SB_T1_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_OUT_B1;
	assign SB_T1_EAST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T1_EAST_SB_OUT_B17;
	assign SB_T1_EAST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T1_EAST_SB_OUT_B17_valid_out;
	assign SB_T1_EAST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_OUT_B1_valid_out;
	assign SB_T1_NORTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T1_NORTH_SB_IN_B17_ready_out;
	assign SB_T1_NORTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_IN_B1_ready_out;
	assign SB_T1_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_OUT_B1;
	assign SB_T1_NORTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T1_NORTH_SB_OUT_B17;
	assign SB_T1_NORTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T1_NORTH_SB_OUT_B17_valid_out;
	assign SB_T1_NORTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_OUT_B1_valid_out;
	assign SB_T1_SOUTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T1_SOUTH_SB_IN_B17_ready_out;
	assign SB_T1_SOUTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_IN_B1_ready_out;
	assign SB_T1_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_OUT_B1;
	assign SB_T1_SOUTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T1_SOUTH_SB_OUT_B17;
	assign SB_T1_SOUTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T1_SOUTH_SB_OUT_B17_valid_out;
	assign SB_T1_SOUTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_OUT_B1_valid_out;
	assign SB_T1_WEST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T1_WEST_SB_IN_B17_ready_out;
	assign SB_T1_WEST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_IN_B1_ready_out;
	assign SB_T1_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_OUT_B1;
	assign SB_T1_WEST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T1_WEST_SB_OUT_B17;
	assign SB_T1_WEST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T1_WEST_SB_OUT_B17_valid_out;
	assign SB_T1_WEST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_OUT_B1_valid_out;
	assign SB_T2_EAST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T2_EAST_SB_IN_B17_ready_out;
	assign SB_T2_EAST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_IN_B1_ready_out;
	assign SB_T2_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_OUT_B1;
	assign SB_T2_EAST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T2_EAST_SB_OUT_B17;
	assign SB_T2_EAST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T2_EAST_SB_OUT_B17_valid_out;
	assign SB_T2_EAST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_OUT_B1_valid_out;
	assign SB_T2_NORTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T2_NORTH_SB_IN_B17_ready_out;
	assign SB_T2_NORTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_IN_B1_ready_out;
	assign SB_T2_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_OUT_B1;
	assign SB_T2_NORTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T2_NORTH_SB_OUT_B17;
	assign SB_T2_NORTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T2_NORTH_SB_OUT_B17_valid_out;
	assign SB_T2_NORTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_OUT_B1_valid_out;
	assign SB_T2_SOUTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T2_SOUTH_SB_IN_B17_ready_out;
	assign SB_T2_SOUTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_IN_B1_ready_out;
	assign SB_T2_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_OUT_B1;
	assign SB_T2_SOUTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T2_SOUTH_SB_OUT_B17;
	assign SB_T2_SOUTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T2_SOUTH_SB_OUT_B17_valid_out;
	assign SB_T2_SOUTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_OUT_B1_valid_out;
	assign SB_T2_WEST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T2_WEST_SB_IN_B17_ready_out;
	assign SB_T2_WEST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_IN_B1_ready_out;
	assign SB_T2_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_OUT_B1;
	assign SB_T2_WEST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T2_WEST_SB_OUT_B17;
	assign SB_T2_WEST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T2_WEST_SB_OUT_B17_valid_out;
	assign SB_T2_WEST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_OUT_B1_valid_out;
	assign SB_T3_EAST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T3_EAST_SB_IN_B17_ready_out;
	assign SB_T3_EAST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_IN_B1_ready_out;
	assign SB_T3_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_OUT_B1;
	assign SB_T3_EAST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T3_EAST_SB_OUT_B17;
	assign SB_T3_EAST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T3_EAST_SB_OUT_B17_valid_out;
	assign SB_T3_EAST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_OUT_B1_valid_out;
	assign SB_T3_NORTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T3_NORTH_SB_IN_B17_ready_out;
	assign SB_T3_NORTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_IN_B1_ready_out;
	assign SB_T3_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_OUT_B1;
	assign SB_T3_NORTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T3_NORTH_SB_OUT_B17;
	assign SB_T3_NORTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T3_NORTH_SB_OUT_B17_valid_out;
	assign SB_T3_NORTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_OUT_B1_valid_out;
	assign SB_T3_SOUTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T3_SOUTH_SB_IN_B17_ready_out;
	assign SB_T3_SOUTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_IN_B1_ready_out;
	assign SB_T3_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_OUT_B1;
	assign SB_T3_SOUTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T3_SOUTH_SB_OUT_B17;
	assign SB_T3_SOUTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T3_SOUTH_SB_OUT_B17_valid_out;
	assign SB_T3_SOUTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_OUT_B1_valid_out;
	assign SB_T3_WEST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T3_WEST_SB_IN_B17_ready_out;
	assign SB_T3_WEST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_IN_B1_ready_out;
	assign SB_T3_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_OUT_B1;
	assign SB_T3_WEST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T3_WEST_SB_OUT_B17;
	assign SB_T3_WEST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T3_WEST_SB_OUT_B17_valid_out;
	assign SB_T3_WEST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_OUT_B1_valid_out;
	assign SB_T4_EAST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T4_EAST_SB_IN_B17_ready_out;
	assign SB_T4_EAST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_IN_B1_ready_out;
	assign SB_T4_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_OUT_B1;
	assign SB_T4_EAST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T4_EAST_SB_OUT_B17;
	assign SB_T4_EAST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T4_EAST_SB_OUT_B17_valid_out;
	assign SB_T4_EAST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_OUT_B1_valid_out;
	assign SB_T4_NORTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T4_NORTH_SB_IN_B17_ready_out;
	assign SB_T4_NORTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_IN_B1_ready_out;
	assign SB_T4_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_OUT_B1;
	assign SB_T4_NORTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T4_NORTH_SB_OUT_B17;
	assign SB_T4_NORTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T4_NORTH_SB_OUT_B17_valid_out;
	assign SB_T4_NORTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_OUT_B1_valid_out;
	assign SB_T4_SOUTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T4_SOUTH_SB_IN_B17_ready_out;
	assign SB_T4_SOUTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_IN_B1_ready_out;
	assign SB_T4_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_OUT_B1;
	assign SB_T4_SOUTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T4_SOUTH_SB_OUT_B17;
	assign SB_T4_SOUTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T4_SOUTH_SB_OUT_B17_valid_out;
	assign SB_T4_SOUTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_OUT_B1_valid_out;
	assign SB_T4_WEST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T4_WEST_SB_IN_B17_ready_out;
	assign SB_T4_WEST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_IN_B1_ready_out;
	assign SB_T4_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_OUT_B1;
	assign SB_T4_WEST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T4_WEST_SB_OUT_B17;
	assign SB_T4_WEST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T4_WEST_SB_OUT_B17_valid_out;
	assign SB_T4_WEST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_OUT_B1_valid_out;
	assign clk_out = coreir_wrapOutClock_inst0_out;
	assign clk_pass_through_out_bot = clk_pass_through;
	assign clk_pass_through_out_right = coreir_wrapOutClock_inst1_out;
	assign config_out_config_addr = config_config_addr;
	assign config_out_config_data = config_config_data;
	assign config_out_read = config_read;
	assign config_out_write = config_write;
	assign flush_out = flush;
	assign hi = const_511_9_out;
	assign lo = const_0_8_out;
	assign read_config_data = PowerDomainOR_O;
	assign reset_out = reset;
	assign stall_out = stall;
endmodule
module CB_MEM_input_width_1_num_1 (
	I,
	O,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	enable,
	out_sel,
	read_config_data,
	ready_in,
	ready_out,
	reset,
	valid_in,
	valid_out
);
	input [19:0] I;
	output wire [0:0] O;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output wire enable;
	output wire [31:0] out_sel;
	output wire [31:0] read_config_data;
	input ready_in;
	output wire ready_out;
	input reset;
	input [19:0] valid_in;
	output wire valid_out;
	wire [0:0] CB_MEM_input_width_1_num_1_O;
	wire CB_MEM_input_width_1_num_1_ready_out;
	wire CB_MEM_input_width_1_num_1_valid_out;
	wire [31:0] CB_MEM_input_width_1_num_1_out_sel;
	wire [0:0] CB_MEM_input_width_1_num_1_enable_value_O;
	wire [4:0] CB_MEM_input_width_1_num_1_sel_value_O;
	wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
	wire [5:0] config_reg_0_O;
	wire [19:0] CB_MEM_input_width_1_num_1_I;
	assign CB_MEM_input_width_1_num_1_I[19+:1] = I[19+:1];
	assign CB_MEM_input_width_1_num_1_I[18+:1] = I[18+:1];
	assign CB_MEM_input_width_1_num_1_I[17+:1] = I[17+:1];
	assign CB_MEM_input_width_1_num_1_I[16+:1] = I[16+:1];
	assign CB_MEM_input_width_1_num_1_I[15+:1] = I[15+:1];
	assign CB_MEM_input_width_1_num_1_I[14+:1] = I[14+:1];
	assign CB_MEM_input_width_1_num_1_I[13+:1] = I[13+:1];
	assign CB_MEM_input_width_1_num_1_I[12+:1] = I[12+:1];
	assign CB_MEM_input_width_1_num_1_I[11+:1] = I[11+:1];
	assign CB_MEM_input_width_1_num_1_I[10+:1] = I[10+:1];
	assign CB_MEM_input_width_1_num_1_I[9+:1] = I[9+:1];
	assign CB_MEM_input_width_1_num_1_I[8+:1] = I[8+:1];
	assign CB_MEM_input_width_1_num_1_I[7+:1] = I[7+:1];
	assign CB_MEM_input_width_1_num_1_I[6+:1] = I[6+:1];
	assign CB_MEM_input_width_1_num_1_I[5+:1] = I[5+:1];
	assign CB_MEM_input_width_1_num_1_I[4+:1] = I[4+:1];
	assign CB_MEM_input_width_1_num_1_I[3+:1] = I[3+:1];
	assign CB_MEM_input_width_1_num_1_I[2+:1] = I[2+:1];
	assign CB_MEM_input_width_1_num_1_I[1+:1] = I[1+:1];
	assign CB_MEM_input_width_1_num_1_I[0+:1] = I[0+:1];
	mux_aoi_ready_valid_const_20_1 CB_MEM_input_width_1_num_1(
		.I(CB_MEM_input_width_1_num_1_I),
		.O(CB_MEM_input_width_1_num_1_O),
		.ready_in(ready_in),
		.ready_out(CB_MEM_input_width_1_num_1_ready_out),
		.valid_in(valid_in),
		.valid_out(CB_MEM_input_width_1_num_1_valid_out),
		.S(CB_MEM_input_width_1_num_1_sel_value_O),
		.out_sel(CB_MEM_input_width_1_num_1_out_sel)
	);
	SliceWrapper_6_0_1 CB_MEM_input_width_1_num_1_enable_value(
		.I(config_reg_0_O),
		.O(CB_MEM_input_width_1_num_1_enable_value_O)
	);
	SliceWrapper_6_1_6 CB_MEM_input_width_1_num_1_sel_value(
		.I(config_reg_0_O),
		.O(CB_MEM_input_width_1_num_1_sel_value_O)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_6_32_inst0$bit_const_0_None(.out(ZextWrapper_6_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
	assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, config_reg_0_O};
	mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O(
		.in(ZextWrapper_6_32_inst0$self_O_in),
		.out(ZextWrapper_6_32_inst0$self_O_out)
	);
	ConfigRegister_6_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	assign O = CB_MEM_input_width_1_num_1_O;
	assign enable = CB_MEM_input_width_1_num_1_enable_value_O[0];
	assign out_sel = CB_MEM_input_width_1_num_1_out_sel;
	assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
	assign ready_out = CB_MEM_input_width_1_num_1_ready_out;
	assign valid_out = CB_MEM_input_width_1_num_1_valid_out;
endmodule
module CB_MEM_input_width_1_num_0 (
	I,
	O,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	enable,
	out_sel,
	read_config_data,
	ready_in,
	ready_out,
	reset,
	valid_in,
	valid_out
);
	input [19:0] I;
	output wire [0:0] O;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output wire enable;
	output wire [31:0] out_sel;
	output wire [31:0] read_config_data;
	input ready_in;
	output wire ready_out;
	input reset;
	input [19:0] valid_in;
	output wire valid_out;
	wire [0:0] CB_MEM_input_width_1_num_0_O;
	wire CB_MEM_input_width_1_num_0_ready_out;
	wire CB_MEM_input_width_1_num_0_valid_out;
	wire [31:0] CB_MEM_input_width_1_num_0_out_sel;
	wire [0:0] CB_MEM_input_width_1_num_0_enable_value_O;
	wire [4:0] CB_MEM_input_width_1_num_0_sel_value_O;
	wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
	wire [5:0] config_reg_0_O;
	wire [19:0] CB_MEM_input_width_1_num_0_I;
	assign CB_MEM_input_width_1_num_0_I[19+:1] = I[19+:1];
	assign CB_MEM_input_width_1_num_0_I[18+:1] = I[18+:1];
	assign CB_MEM_input_width_1_num_0_I[17+:1] = I[17+:1];
	assign CB_MEM_input_width_1_num_0_I[16+:1] = I[16+:1];
	assign CB_MEM_input_width_1_num_0_I[15+:1] = I[15+:1];
	assign CB_MEM_input_width_1_num_0_I[14+:1] = I[14+:1];
	assign CB_MEM_input_width_1_num_0_I[13+:1] = I[13+:1];
	assign CB_MEM_input_width_1_num_0_I[12+:1] = I[12+:1];
	assign CB_MEM_input_width_1_num_0_I[11+:1] = I[11+:1];
	assign CB_MEM_input_width_1_num_0_I[10+:1] = I[10+:1];
	assign CB_MEM_input_width_1_num_0_I[9+:1] = I[9+:1];
	assign CB_MEM_input_width_1_num_0_I[8+:1] = I[8+:1];
	assign CB_MEM_input_width_1_num_0_I[7+:1] = I[7+:1];
	assign CB_MEM_input_width_1_num_0_I[6+:1] = I[6+:1];
	assign CB_MEM_input_width_1_num_0_I[5+:1] = I[5+:1];
	assign CB_MEM_input_width_1_num_0_I[4+:1] = I[4+:1];
	assign CB_MEM_input_width_1_num_0_I[3+:1] = I[3+:1];
	assign CB_MEM_input_width_1_num_0_I[2+:1] = I[2+:1];
	assign CB_MEM_input_width_1_num_0_I[1+:1] = I[1+:1];
	assign CB_MEM_input_width_1_num_0_I[0+:1] = I[0+:1];
	mux_aoi_ready_valid_const_20_1 CB_MEM_input_width_1_num_0(
		.I(CB_MEM_input_width_1_num_0_I),
		.O(CB_MEM_input_width_1_num_0_O),
		.ready_in(ready_in),
		.ready_out(CB_MEM_input_width_1_num_0_ready_out),
		.valid_in(valid_in),
		.valid_out(CB_MEM_input_width_1_num_0_valid_out),
		.S(CB_MEM_input_width_1_num_0_sel_value_O),
		.out_sel(CB_MEM_input_width_1_num_0_out_sel)
	);
	SliceWrapper_6_0_1 CB_MEM_input_width_1_num_0_enable_value(
		.I(config_reg_0_O),
		.O(CB_MEM_input_width_1_num_0_enable_value_O)
	);
	SliceWrapper_6_1_6 CB_MEM_input_width_1_num_0_sel_value(
		.I(config_reg_0_O),
		.O(CB_MEM_input_width_1_num_0_sel_value_O)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_6_32_inst0$bit_const_0_None(.out(ZextWrapper_6_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
	assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, config_reg_0_O};
	mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O(
		.in(ZextWrapper_6_32_inst0$self_O_in),
		.out(ZextWrapper_6_32_inst0$self_O_out)
	);
	ConfigRegister_6_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	assign O = CB_MEM_input_width_1_num_0_O;
	assign enable = CB_MEM_input_width_1_num_0_enable_value_O[0];
	assign out_sel = CB_MEM_input_width_1_num_0_out_sel;
	assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
	assign ready_out = CB_MEM_input_width_1_num_0_ready_out;
	assign valid_out = CB_MEM_input_width_1_num_0_valid_out;
endmodule
module CB_MEM_input_width_17_num_3 (
	I,
	O,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	enable,
	out_sel,
	read_config_data,
	ready_in,
	ready_out,
	reset,
	valid_in,
	valid_out
);
	input [339:0] I;
	output wire [16:0] O;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output wire enable;
	output wire [31:0] out_sel;
	output wire [31:0] read_config_data;
	input ready_in;
	output wire ready_out;
	input reset;
	input [19:0] valid_in;
	output wire valid_out;
	wire [16:0] CB_MEM_input_width_17_num_3_O;
	wire CB_MEM_input_width_17_num_3_ready_out;
	wire CB_MEM_input_width_17_num_3_valid_out;
	wire [31:0] CB_MEM_input_width_17_num_3_out_sel;
	wire [0:0] CB_MEM_input_width_17_num_3_enable_value_O;
	wire [4:0] CB_MEM_input_width_17_num_3_sel_value_O;
	wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
	wire [5:0] config_reg_0_O;
	wire [339:0] CB_MEM_input_width_17_num_3_I;
	assign CB_MEM_input_width_17_num_3_I[323+:17] = I[323+:17];
	assign CB_MEM_input_width_17_num_3_I[306+:17] = I[306+:17];
	assign CB_MEM_input_width_17_num_3_I[289+:17] = I[289+:17];
	assign CB_MEM_input_width_17_num_3_I[272+:17] = I[272+:17];
	assign CB_MEM_input_width_17_num_3_I[255+:17] = I[255+:17];
	assign CB_MEM_input_width_17_num_3_I[238+:17] = I[238+:17];
	assign CB_MEM_input_width_17_num_3_I[221+:17] = I[221+:17];
	assign CB_MEM_input_width_17_num_3_I[204+:17] = I[204+:17];
	assign CB_MEM_input_width_17_num_3_I[187+:17] = I[187+:17];
	assign CB_MEM_input_width_17_num_3_I[170+:17] = I[170+:17];
	assign CB_MEM_input_width_17_num_3_I[153+:17] = I[153+:17];
	assign CB_MEM_input_width_17_num_3_I[136+:17] = I[136+:17];
	assign CB_MEM_input_width_17_num_3_I[119+:17] = I[119+:17];
	assign CB_MEM_input_width_17_num_3_I[102+:17] = I[102+:17];
	assign CB_MEM_input_width_17_num_3_I[85+:17] = I[85+:17];
	assign CB_MEM_input_width_17_num_3_I[68+:17] = I[68+:17];
	assign CB_MEM_input_width_17_num_3_I[51+:17] = I[51+:17];
	assign CB_MEM_input_width_17_num_3_I[34+:17] = I[34+:17];
	assign CB_MEM_input_width_17_num_3_I[17+:17] = I[17+:17];
	assign CB_MEM_input_width_17_num_3_I[0+:17] = I[0+:17];
	mux_aoi_ready_valid_const_20_17 CB_MEM_input_width_17_num_3(
		.I(CB_MEM_input_width_17_num_3_I),
		.O(CB_MEM_input_width_17_num_3_O),
		.ready_in(ready_in),
		.ready_out(CB_MEM_input_width_17_num_3_ready_out),
		.valid_in(valid_in),
		.valid_out(CB_MEM_input_width_17_num_3_valid_out),
		.S(CB_MEM_input_width_17_num_3_sel_value_O),
		.out_sel(CB_MEM_input_width_17_num_3_out_sel)
	);
	SliceWrapper_6_0_1 CB_MEM_input_width_17_num_3_enable_value(
		.I(config_reg_0_O),
		.O(CB_MEM_input_width_17_num_3_enable_value_O)
	);
	SliceWrapper_6_1_6 CB_MEM_input_width_17_num_3_sel_value(
		.I(config_reg_0_O),
		.O(CB_MEM_input_width_17_num_3_sel_value_O)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_6_32_inst0$bit_const_0_None(.out(ZextWrapper_6_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
	assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, config_reg_0_O};
	mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O(
		.in(ZextWrapper_6_32_inst0$self_O_in),
		.out(ZextWrapper_6_32_inst0$self_O_out)
	);
	ConfigRegister_6_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	assign O = CB_MEM_input_width_17_num_3_O;
	assign enable = CB_MEM_input_width_17_num_3_enable_value_O[0];
	assign out_sel = CB_MEM_input_width_17_num_3_out_sel;
	assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
	assign ready_out = CB_MEM_input_width_17_num_3_ready_out;
	assign valid_out = CB_MEM_input_width_17_num_3_valid_out;
endmodule
module CB_MEM_input_width_17_num_2 (
	I,
	O,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	enable,
	out_sel,
	read_config_data,
	ready_in,
	ready_out,
	reset,
	valid_in,
	valid_out
);
	input [339:0] I;
	output wire [16:0] O;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output wire enable;
	output wire [31:0] out_sel;
	output wire [31:0] read_config_data;
	input ready_in;
	output wire ready_out;
	input reset;
	input [19:0] valid_in;
	output wire valid_out;
	wire [16:0] CB_MEM_input_width_17_num_2_O;
	wire CB_MEM_input_width_17_num_2_ready_out;
	wire CB_MEM_input_width_17_num_2_valid_out;
	wire [31:0] CB_MEM_input_width_17_num_2_out_sel;
	wire [0:0] CB_MEM_input_width_17_num_2_enable_value_O;
	wire [4:0] CB_MEM_input_width_17_num_2_sel_value_O;
	wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
	wire [5:0] config_reg_0_O;
	wire [339:0] CB_MEM_input_width_17_num_2_I;
	assign CB_MEM_input_width_17_num_2_I[323+:17] = I[323+:17];
	assign CB_MEM_input_width_17_num_2_I[306+:17] = I[306+:17];
	assign CB_MEM_input_width_17_num_2_I[289+:17] = I[289+:17];
	assign CB_MEM_input_width_17_num_2_I[272+:17] = I[272+:17];
	assign CB_MEM_input_width_17_num_2_I[255+:17] = I[255+:17];
	assign CB_MEM_input_width_17_num_2_I[238+:17] = I[238+:17];
	assign CB_MEM_input_width_17_num_2_I[221+:17] = I[221+:17];
	assign CB_MEM_input_width_17_num_2_I[204+:17] = I[204+:17];
	assign CB_MEM_input_width_17_num_2_I[187+:17] = I[187+:17];
	assign CB_MEM_input_width_17_num_2_I[170+:17] = I[170+:17];
	assign CB_MEM_input_width_17_num_2_I[153+:17] = I[153+:17];
	assign CB_MEM_input_width_17_num_2_I[136+:17] = I[136+:17];
	assign CB_MEM_input_width_17_num_2_I[119+:17] = I[119+:17];
	assign CB_MEM_input_width_17_num_2_I[102+:17] = I[102+:17];
	assign CB_MEM_input_width_17_num_2_I[85+:17] = I[85+:17];
	assign CB_MEM_input_width_17_num_2_I[68+:17] = I[68+:17];
	assign CB_MEM_input_width_17_num_2_I[51+:17] = I[51+:17];
	assign CB_MEM_input_width_17_num_2_I[34+:17] = I[34+:17];
	assign CB_MEM_input_width_17_num_2_I[17+:17] = I[17+:17];
	assign CB_MEM_input_width_17_num_2_I[0+:17] = I[0+:17];
	mux_aoi_ready_valid_const_20_17 CB_MEM_input_width_17_num_2(
		.I(CB_MEM_input_width_17_num_2_I),
		.O(CB_MEM_input_width_17_num_2_O),
		.ready_in(ready_in),
		.ready_out(CB_MEM_input_width_17_num_2_ready_out),
		.valid_in(valid_in),
		.valid_out(CB_MEM_input_width_17_num_2_valid_out),
		.S(CB_MEM_input_width_17_num_2_sel_value_O),
		.out_sel(CB_MEM_input_width_17_num_2_out_sel)
	);
	SliceWrapper_6_0_1 CB_MEM_input_width_17_num_2_enable_value(
		.I(config_reg_0_O),
		.O(CB_MEM_input_width_17_num_2_enable_value_O)
	);
	SliceWrapper_6_1_6 CB_MEM_input_width_17_num_2_sel_value(
		.I(config_reg_0_O),
		.O(CB_MEM_input_width_17_num_2_sel_value_O)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_6_32_inst0$bit_const_0_None(.out(ZextWrapper_6_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
	assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, config_reg_0_O};
	mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O(
		.in(ZextWrapper_6_32_inst0$self_O_in),
		.out(ZextWrapper_6_32_inst0$self_O_out)
	);
	ConfigRegister_6_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	assign O = CB_MEM_input_width_17_num_2_O;
	assign enable = CB_MEM_input_width_17_num_2_enable_value_O[0];
	assign out_sel = CB_MEM_input_width_17_num_2_out_sel;
	assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
	assign ready_out = CB_MEM_input_width_17_num_2_ready_out;
	assign valid_out = CB_MEM_input_width_17_num_2_valid_out;
endmodule
module CB_MEM_input_width_17_num_1 (
	I,
	O,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	enable,
	out_sel,
	read_config_data,
	ready_in,
	ready_out,
	reset,
	valid_in,
	valid_out
);
	input [339:0] I;
	output wire [16:0] O;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output wire enable;
	output wire [31:0] out_sel;
	output wire [31:0] read_config_data;
	input ready_in;
	output wire ready_out;
	input reset;
	input [19:0] valid_in;
	output wire valid_out;
	wire [16:0] CB_MEM_input_width_17_num_1_O;
	wire CB_MEM_input_width_17_num_1_ready_out;
	wire CB_MEM_input_width_17_num_1_valid_out;
	wire [31:0] CB_MEM_input_width_17_num_1_out_sel;
	wire [0:0] CB_MEM_input_width_17_num_1_enable_value_O;
	wire [4:0] CB_MEM_input_width_17_num_1_sel_value_O;
	wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
	wire [5:0] config_reg_0_O;
	wire [339:0] CB_MEM_input_width_17_num_1_I;
	assign CB_MEM_input_width_17_num_1_I[323+:17] = I[323+:17];
	assign CB_MEM_input_width_17_num_1_I[306+:17] = I[306+:17];
	assign CB_MEM_input_width_17_num_1_I[289+:17] = I[289+:17];
	assign CB_MEM_input_width_17_num_1_I[272+:17] = I[272+:17];
	assign CB_MEM_input_width_17_num_1_I[255+:17] = I[255+:17];
	assign CB_MEM_input_width_17_num_1_I[238+:17] = I[238+:17];
	assign CB_MEM_input_width_17_num_1_I[221+:17] = I[221+:17];
	assign CB_MEM_input_width_17_num_1_I[204+:17] = I[204+:17];
	assign CB_MEM_input_width_17_num_1_I[187+:17] = I[187+:17];
	assign CB_MEM_input_width_17_num_1_I[170+:17] = I[170+:17];
	assign CB_MEM_input_width_17_num_1_I[153+:17] = I[153+:17];
	assign CB_MEM_input_width_17_num_1_I[136+:17] = I[136+:17];
	assign CB_MEM_input_width_17_num_1_I[119+:17] = I[119+:17];
	assign CB_MEM_input_width_17_num_1_I[102+:17] = I[102+:17];
	assign CB_MEM_input_width_17_num_1_I[85+:17] = I[85+:17];
	assign CB_MEM_input_width_17_num_1_I[68+:17] = I[68+:17];
	assign CB_MEM_input_width_17_num_1_I[51+:17] = I[51+:17];
	assign CB_MEM_input_width_17_num_1_I[34+:17] = I[34+:17];
	assign CB_MEM_input_width_17_num_1_I[17+:17] = I[17+:17];
	assign CB_MEM_input_width_17_num_1_I[0+:17] = I[0+:17];
	mux_aoi_ready_valid_const_20_17 CB_MEM_input_width_17_num_1(
		.I(CB_MEM_input_width_17_num_1_I),
		.O(CB_MEM_input_width_17_num_1_O),
		.ready_in(ready_in),
		.ready_out(CB_MEM_input_width_17_num_1_ready_out),
		.valid_in(valid_in),
		.valid_out(CB_MEM_input_width_17_num_1_valid_out),
		.S(CB_MEM_input_width_17_num_1_sel_value_O),
		.out_sel(CB_MEM_input_width_17_num_1_out_sel)
	);
	SliceWrapper_6_0_1 CB_MEM_input_width_17_num_1_enable_value(
		.I(config_reg_0_O),
		.O(CB_MEM_input_width_17_num_1_enable_value_O)
	);
	SliceWrapper_6_1_6 CB_MEM_input_width_17_num_1_sel_value(
		.I(config_reg_0_O),
		.O(CB_MEM_input_width_17_num_1_sel_value_O)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_6_32_inst0$bit_const_0_None(.out(ZextWrapper_6_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
	assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, config_reg_0_O};
	mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O(
		.in(ZextWrapper_6_32_inst0$self_O_in),
		.out(ZextWrapper_6_32_inst0$self_O_out)
	);
	ConfigRegister_6_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	assign O = CB_MEM_input_width_17_num_1_O;
	assign enable = CB_MEM_input_width_17_num_1_enable_value_O[0];
	assign out_sel = CB_MEM_input_width_17_num_1_out_sel;
	assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
	assign ready_out = CB_MEM_input_width_17_num_1_ready_out;
	assign valid_out = CB_MEM_input_width_17_num_1_valid_out;
endmodule
module CB_MEM_input_width_17_num_0 (
	I,
	O,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	enable,
	out_sel,
	read_config_data,
	ready_in,
	ready_out,
	reset,
	valid_in,
	valid_out
);
	input [339:0] I;
	output wire [16:0] O;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output wire enable;
	output wire [31:0] out_sel;
	output wire [31:0] read_config_data;
	input ready_in;
	output wire ready_out;
	input reset;
	input [19:0] valid_in;
	output wire valid_out;
	wire [16:0] CB_MEM_input_width_17_num_0_O;
	wire CB_MEM_input_width_17_num_0_ready_out;
	wire CB_MEM_input_width_17_num_0_valid_out;
	wire [31:0] CB_MEM_input_width_17_num_0_out_sel;
	wire [0:0] CB_MEM_input_width_17_num_0_enable_value_O;
	wire [4:0] CB_MEM_input_width_17_num_0_sel_value_O;
	wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
	wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
	wire [5:0] config_reg_0_O;
	wire [339:0] CB_MEM_input_width_17_num_0_I;
	assign CB_MEM_input_width_17_num_0_I[323+:17] = I[323+:17];
	assign CB_MEM_input_width_17_num_0_I[306+:17] = I[306+:17];
	assign CB_MEM_input_width_17_num_0_I[289+:17] = I[289+:17];
	assign CB_MEM_input_width_17_num_0_I[272+:17] = I[272+:17];
	assign CB_MEM_input_width_17_num_0_I[255+:17] = I[255+:17];
	assign CB_MEM_input_width_17_num_0_I[238+:17] = I[238+:17];
	assign CB_MEM_input_width_17_num_0_I[221+:17] = I[221+:17];
	assign CB_MEM_input_width_17_num_0_I[204+:17] = I[204+:17];
	assign CB_MEM_input_width_17_num_0_I[187+:17] = I[187+:17];
	assign CB_MEM_input_width_17_num_0_I[170+:17] = I[170+:17];
	assign CB_MEM_input_width_17_num_0_I[153+:17] = I[153+:17];
	assign CB_MEM_input_width_17_num_0_I[136+:17] = I[136+:17];
	assign CB_MEM_input_width_17_num_0_I[119+:17] = I[119+:17];
	assign CB_MEM_input_width_17_num_0_I[102+:17] = I[102+:17];
	assign CB_MEM_input_width_17_num_0_I[85+:17] = I[85+:17];
	assign CB_MEM_input_width_17_num_0_I[68+:17] = I[68+:17];
	assign CB_MEM_input_width_17_num_0_I[51+:17] = I[51+:17];
	assign CB_MEM_input_width_17_num_0_I[34+:17] = I[34+:17];
	assign CB_MEM_input_width_17_num_0_I[17+:17] = I[17+:17];
	assign CB_MEM_input_width_17_num_0_I[0+:17] = I[0+:17];
	mux_aoi_ready_valid_const_20_17 CB_MEM_input_width_17_num_0(
		.I(CB_MEM_input_width_17_num_0_I),
		.O(CB_MEM_input_width_17_num_0_O),
		.ready_in(ready_in),
		.ready_out(CB_MEM_input_width_17_num_0_ready_out),
		.valid_in(valid_in),
		.valid_out(CB_MEM_input_width_17_num_0_valid_out),
		.S(CB_MEM_input_width_17_num_0_sel_value_O),
		.out_sel(CB_MEM_input_width_17_num_0_out_sel)
	);
	SliceWrapper_6_0_1 CB_MEM_input_width_17_num_0_enable_value(
		.I(config_reg_0_O),
		.O(CB_MEM_input_width_17_num_0_enable_value_O)
	);
	SliceWrapper_6_1_6 CB_MEM_input_width_17_num_0_sel_value(
		.I(config_reg_0_O),
		.O(CB_MEM_input_width_17_num_0_sel_value_O)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_6_32_inst0$bit_const_0_None(.out(ZextWrapper_6_32_inst0$bit_const_0_None_out));
	wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
	assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, ZextWrapper_6_32_inst0$bit_const_0_None_out, config_reg_0_O};
	mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O(
		.in(ZextWrapper_6_32_inst0$self_O_in),
		.out(ZextWrapper_6_32_inst0$self_O_out)
	);
	ConfigRegister_6_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	assign O = CB_MEM_input_width_17_num_0_O;
	assign enable = CB_MEM_input_width_17_num_0_enable_value_O[0];
	assign out_sel = CB_MEM_input_width_17_num_0_out_sel;
	assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
	assign ready_out = CB_MEM_input_width_17_num_0_ready_out;
	assign valid_out = CB_MEM_input_width_17_num_0_valid_out;
endmodule
module Tile_MemCore (
	SB_T0_EAST_SB_IN_B1,
	SB_T0_EAST_SB_IN_B17,
	SB_T0_EAST_SB_IN_B17_ready,
	SB_T0_EAST_SB_IN_B17_valid,
	SB_T0_EAST_SB_IN_B1_ready,
	SB_T0_EAST_SB_IN_B1_valid,
	SB_T0_EAST_SB_OUT_B1,
	SB_T0_EAST_SB_OUT_B17,
	SB_T0_EAST_SB_OUT_B17_ready,
	SB_T0_EAST_SB_OUT_B17_valid,
	SB_T0_EAST_SB_OUT_B1_ready,
	SB_T0_EAST_SB_OUT_B1_valid,
	SB_T0_NORTH_SB_IN_B1,
	SB_T0_NORTH_SB_IN_B17,
	SB_T0_NORTH_SB_IN_B17_ready,
	SB_T0_NORTH_SB_IN_B17_valid,
	SB_T0_NORTH_SB_IN_B1_ready,
	SB_T0_NORTH_SB_IN_B1_valid,
	SB_T0_NORTH_SB_OUT_B1,
	SB_T0_NORTH_SB_OUT_B17,
	SB_T0_NORTH_SB_OUT_B17_ready,
	SB_T0_NORTH_SB_OUT_B17_valid,
	SB_T0_NORTH_SB_OUT_B1_ready,
	SB_T0_NORTH_SB_OUT_B1_valid,
	SB_T0_SOUTH_SB_IN_B1,
	SB_T0_SOUTH_SB_IN_B17,
	SB_T0_SOUTH_SB_IN_B17_ready,
	SB_T0_SOUTH_SB_IN_B17_valid,
	SB_T0_SOUTH_SB_IN_B1_ready,
	SB_T0_SOUTH_SB_IN_B1_valid,
	SB_T0_SOUTH_SB_OUT_B1,
	SB_T0_SOUTH_SB_OUT_B17,
	SB_T0_SOUTH_SB_OUT_B17_ready,
	SB_T0_SOUTH_SB_OUT_B17_valid,
	SB_T0_SOUTH_SB_OUT_B1_ready,
	SB_T0_SOUTH_SB_OUT_B1_valid,
	SB_T0_WEST_SB_IN_B1,
	SB_T0_WEST_SB_IN_B17,
	SB_T0_WEST_SB_IN_B17_ready,
	SB_T0_WEST_SB_IN_B17_valid,
	SB_T0_WEST_SB_IN_B1_ready,
	SB_T0_WEST_SB_IN_B1_valid,
	SB_T0_WEST_SB_OUT_B1,
	SB_T0_WEST_SB_OUT_B17,
	SB_T0_WEST_SB_OUT_B17_ready,
	SB_T0_WEST_SB_OUT_B17_valid,
	SB_T0_WEST_SB_OUT_B1_ready,
	SB_T0_WEST_SB_OUT_B1_valid,
	SB_T1_EAST_SB_IN_B1,
	SB_T1_EAST_SB_IN_B17,
	SB_T1_EAST_SB_IN_B17_ready,
	SB_T1_EAST_SB_IN_B17_valid,
	SB_T1_EAST_SB_IN_B1_ready,
	SB_T1_EAST_SB_IN_B1_valid,
	SB_T1_EAST_SB_OUT_B1,
	SB_T1_EAST_SB_OUT_B17,
	SB_T1_EAST_SB_OUT_B17_ready,
	SB_T1_EAST_SB_OUT_B17_valid,
	SB_T1_EAST_SB_OUT_B1_ready,
	SB_T1_EAST_SB_OUT_B1_valid,
	SB_T1_NORTH_SB_IN_B1,
	SB_T1_NORTH_SB_IN_B17,
	SB_T1_NORTH_SB_IN_B17_ready,
	SB_T1_NORTH_SB_IN_B17_valid,
	SB_T1_NORTH_SB_IN_B1_ready,
	SB_T1_NORTH_SB_IN_B1_valid,
	SB_T1_NORTH_SB_OUT_B1,
	SB_T1_NORTH_SB_OUT_B17,
	SB_T1_NORTH_SB_OUT_B17_ready,
	SB_T1_NORTH_SB_OUT_B17_valid,
	SB_T1_NORTH_SB_OUT_B1_ready,
	SB_T1_NORTH_SB_OUT_B1_valid,
	SB_T1_SOUTH_SB_IN_B1,
	SB_T1_SOUTH_SB_IN_B17,
	SB_T1_SOUTH_SB_IN_B17_ready,
	SB_T1_SOUTH_SB_IN_B17_valid,
	SB_T1_SOUTH_SB_IN_B1_ready,
	SB_T1_SOUTH_SB_IN_B1_valid,
	SB_T1_SOUTH_SB_OUT_B1,
	SB_T1_SOUTH_SB_OUT_B17,
	SB_T1_SOUTH_SB_OUT_B17_ready,
	SB_T1_SOUTH_SB_OUT_B17_valid,
	SB_T1_SOUTH_SB_OUT_B1_ready,
	SB_T1_SOUTH_SB_OUT_B1_valid,
	SB_T1_WEST_SB_IN_B1,
	SB_T1_WEST_SB_IN_B17,
	SB_T1_WEST_SB_IN_B17_ready,
	SB_T1_WEST_SB_IN_B17_valid,
	SB_T1_WEST_SB_IN_B1_ready,
	SB_T1_WEST_SB_IN_B1_valid,
	SB_T1_WEST_SB_OUT_B1,
	SB_T1_WEST_SB_OUT_B17,
	SB_T1_WEST_SB_OUT_B17_ready,
	SB_T1_WEST_SB_OUT_B17_valid,
	SB_T1_WEST_SB_OUT_B1_ready,
	SB_T1_WEST_SB_OUT_B1_valid,
	SB_T2_EAST_SB_IN_B1,
	SB_T2_EAST_SB_IN_B17,
	SB_T2_EAST_SB_IN_B17_ready,
	SB_T2_EAST_SB_IN_B17_valid,
	SB_T2_EAST_SB_IN_B1_ready,
	SB_T2_EAST_SB_IN_B1_valid,
	SB_T2_EAST_SB_OUT_B1,
	SB_T2_EAST_SB_OUT_B17,
	SB_T2_EAST_SB_OUT_B17_ready,
	SB_T2_EAST_SB_OUT_B17_valid,
	SB_T2_EAST_SB_OUT_B1_ready,
	SB_T2_EAST_SB_OUT_B1_valid,
	SB_T2_NORTH_SB_IN_B1,
	SB_T2_NORTH_SB_IN_B17,
	SB_T2_NORTH_SB_IN_B17_ready,
	SB_T2_NORTH_SB_IN_B17_valid,
	SB_T2_NORTH_SB_IN_B1_ready,
	SB_T2_NORTH_SB_IN_B1_valid,
	SB_T2_NORTH_SB_OUT_B1,
	SB_T2_NORTH_SB_OUT_B17,
	SB_T2_NORTH_SB_OUT_B17_ready,
	SB_T2_NORTH_SB_OUT_B17_valid,
	SB_T2_NORTH_SB_OUT_B1_ready,
	SB_T2_NORTH_SB_OUT_B1_valid,
	SB_T2_SOUTH_SB_IN_B1,
	SB_T2_SOUTH_SB_IN_B17,
	SB_T2_SOUTH_SB_IN_B17_ready,
	SB_T2_SOUTH_SB_IN_B17_valid,
	SB_T2_SOUTH_SB_IN_B1_ready,
	SB_T2_SOUTH_SB_IN_B1_valid,
	SB_T2_SOUTH_SB_OUT_B1,
	SB_T2_SOUTH_SB_OUT_B17,
	SB_T2_SOUTH_SB_OUT_B17_ready,
	SB_T2_SOUTH_SB_OUT_B17_valid,
	SB_T2_SOUTH_SB_OUT_B1_ready,
	SB_T2_SOUTH_SB_OUT_B1_valid,
	SB_T2_WEST_SB_IN_B1,
	SB_T2_WEST_SB_IN_B17,
	SB_T2_WEST_SB_IN_B17_ready,
	SB_T2_WEST_SB_IN_B17_valid,
	SB_T2_WEST_SB_IN_B1_ready,
	SB_T2_WEST_SB_IN_B1_valid,
	SB_T2_WEST_SB_OUT_B1,
	SB_T2_WEST_SB_OUT_B17,
	SB_T2_WEST_SB_OUT_B17_ready,
	SB_T2_WEST_SB_OUT_B17_valid,
	SB_T2_WEST_SB_OUT_B1_ready,
	SB_T2_WEST_SB_OUT_B1_valid,
	SB_T3_EAST_SB_IN_B1,
	SB_T3_EAST_SB_IN_B17,
	SB_T3_EAST_SB_IN_B17_ready,
	SB_T3_EAST_SB_IN_B17_valid,
	SB_T3_EAST_SB_IN_B1_ready,
	SB_T3_EAST_SB_IN_B1_valid,
	SB_T3_EAST_SB_OUT_B1,
	SB_T3_EAST_SB_OUT_B17,
	SB_T3_EAST_SB_OUT_B17_ready,
	SB_T3_EAST_SB_OUT_B17_valid,
	SB_T3_EAST_SB_OUT_B1_ready,
	SB_T3_EAST_SB_OUT_B1_valid,
	SB_T3_NORTH_SB_IN_B1,
	SB_T3_NORTH_SB_IN_B17,
	SB_T3_NORTH_SB_IN_B17_ready,
	SB_T3_NORTH_SB_IN_B17_valid,
	SB_T3_NORTH_SB_IN_B1_ready,
	SB_T3_NORTH_SB_IN_B1_valid,
	SB_T3_NORTH_SB_OUT_B1,
	SB_T3_NORTH_SB_OUT_B17,
	SB_T3_NORTH_SB_OUT_B17_ready,
	SB_T3_NORTH_SB_OUT_B17_valid,
	SB_T3_NORTH_SB_OUT_B1_ready,
	SB_T3_NORTH_SB_OUT_B1_valid,
	SB_T3_SOUTH_SB_IN_B1,
	SB_T3_SOUTH_SB_IN_B17,
	SB_T3_SOUTH_SB_IN_B17_ready,
	SB_T3_SOUTH_SB_IN_B17_valid,
	SB_T3_SOUTH_SB_IN_B1_ready,
	SB_T3_SOUTH_SB_IN_B1_valid,
	SB_T3_SOUTH_SB_OUT_B1,
	SB_T3_SOUTH_SB_OUT_B17,
	SB_T3_SOUTH_SB_OUT_B17_ready,
	SB_T3_SOUTH_SB_OUT_B17_valid,
	SB_T3_SOUTH_SB_OUT_B1_ready,
	SB_T3_SOUTH_SB_OUT_B1_valid,
	SB_T3_WEST_SB_IN_B1,
	SB_T3_WEST_SB_IN_B17,
	SB_T3_WEST_SB_IN_B17_ready,
	SB_T3_WEST_SB_IN_B17_valid,
	SB_T3_WEST_SB_IN_B1_ready,
	SB_T3_WEST_SB_IN_B1_valid,
	SB_T3_WEST_SB_OUT_B1,
	SB_T3_WEST_SB_OUT_B17,
	SB_T3_WEST_SB_OUT_B17_ready,
	SB_T3_WEST_SB_OUT_B17_valid,
	SB_T3_WEST_SB_OUT_B1_ready,
	SB_T3_WEST_SB_OUT_B1_valid,
	SB_T4_EAST_SB_IN_B1,
	SB_T4_EAST_SB_IN_B17,
	SB_T4_EAST_SB_IN_B17_ready,
	SB_T4_EAST_SB_IN_B17_valid,
	SB_T4_EAST_SB_IN_B1_ready,
	SB_T4_EAST_SB_IN_B1_valid,
	SB_T4_EAST_SB_OUT_B1,
	SB_T4_EAST_SB_OUT_B17,
	SB_T4_EAST_SB_OUT_B17_ready,
	SB_T4_EAST_SB_OUT_B17_valid,
	SB_T4_EAST_SB_OUT_B1_ready,
	SB_T4_EAST_SB_OUT_B1_valid,
	SB_T4_NORTH_SB_IN_B1,
	SB_T4_NORTH_SB_IN_B17,
	SB_T4_NORTH_SB_IN_B17_ready,
	SB_T4_NORTH_SB_IN_B17_valid,
	SB_T4_NORTH_SB_IN_B1_ready,
	SB_T4_NORTH_SB_IN_B1_valid,
	SB_T4_NORTH_SB_OUT_B1,
	SB_T4_NORTH_SB_OUT_B17,
	SB_T4_NORTH_SB_OUT_B17_ready,
	SB_T4_NORTH_SB_OUT_B17_valid,
	SB_T4_NORTH_SB_OUT_B1_ready,
	SB_T4_NORTH_SB_OUT_B1_valid,
	SB_T4_SOUTH_SB_IN_B1,
	SB_T4_SOUTH_SB_IN_B17,
	SB_T4_SOUTH_SB_IN_B17_ready,
	SB_T4_SOUTH_SB_IN_B17_valid,
	SB_T4_SOUTH_SB_IN_B1_ready,
	SB_T4_SOUTH_SB_IN_B1_valid,
	SB_T4_SOUTH_SB_OUT_B1,
	SB_T4_SOUTH_SB_OUT_B17,
	SB_T4_SOUTH_SB_OUT_B17_ready,
	SB_T4_SOUTH_SB_OUT_B17_valid,
	SB_T4_SOUTH_SB_OUT_B1_ready,
	SB_T4_SOUTH_SB_OUT_B1_valid,
	SB_T4_WEST_SB_IN_B1,
	SB_T4_WEST_SB_IN_B17,
	SB_T4_WEST_SB_IN_B17_ready,
	SB_T4_WEST_SB_IN_B17_valid,
	SB_T4_WEST_SB_IN_B1_ready,
	SB_T4_WEST_SB_IN_B1_valid,
	SB_T4_WEST_SB_OUT_B1,
	SB_T4_WEST_SB_OUT_B17,
	SB_T4_WEST_SB_OUT_B17_ready,
	SB_T4_WEST_SB_OUT_B17_valid,
	SB_T4_WEST_SB_OUT_B1_ready,
	SB_T4_WEST_SB_OUT_B1_valid,
	clk,
	clk_out,
	config_config_addr,
	config_config_data,
	config_out_config_addr,
	config_out_config_data,
	config_out_read,
	config_out_write,
	config_read,
	config_write,
	flush,
	flush_out,
	hi,
	lo,
	read_config_data,
	read_config_data_in,
	reset,
	reset_out,
	stall,
	stall_out,
	tile_id
);
	input [0:0] SB_T0_EAST_SB_IN_B1;
	input [16:0] SB_T0_EAST_SB_IN_B17;
	output wire SB_T0_EAST_SB_IN_B17_ready;
	input SB_T0_EAST_SB_IN_B17_valid;
	output wire SB_T0_EAST_SB_IN_B1_ready;
	input SB_T0_EAST_SB_IN_B1_valid;
	output wire [0:0] SB_T0_EAST_SB_OUT_B1;
	output wire [16:0] SB_T0_EAST_SB_OUT_B17;
	input SB_T0_EAST_SB_OUT_B17_ready;
	output wire SB_T0_EAST_SB_OUT_B17_valid;
	input SB_T0_EAST_SB_OUT_B1_ready;
	output wire SB_T0_EAST_SB_OUT_B1_valid;
	input [0:0] SB_T0_NORTH_SB_IN_B1;
	input [16:0] SB_T0_NORTH_SB_IN_B17;
	output wire SB_T0_NORTH_SB_IN_B17_ready;
	input SB_T0_NORTH_SB_IN_B17_valid;
	output wire SB_T0_NORTH_SB_IN_B1_ready;
	input SB_T0_NORTH_SB_IN_B1_valid;
	output wire [0:0] SB_T0_NORTH_SB_OUT_B1;
	output wire [16:0] SB_T0_NORTH_SB_OUT_B17;
	input SB_T0_NORTH_SB_OUT_B17_ready;
	output wire SB_T0_NORTH_SB_OUT_B17_valid;
	input SB_T0_NORTH_SB_OUT_B1_ready;
	output wire SB_T0_NORTH_SB_OUT_B1_valid;
	input [0:0] SB_T0_SOUTH_SB_IN_B1;
	input [16:0] SB_T0_SOUTH_SB_IN_B17;
	output wire SB_T0_SOUTH_SB_IN_B17_ready;
	input SB_T0_SOUTH_SB_IN_B17_valid;
	output wire SB_T0_SOUTH_SB_IN_B1_ready;
	input SB_T0_SOUTH_SB_IN_B1_valid;
	output wire [0:0] SB_T0_SOUTH_SB_OUT_B1;
	output wire [16:0] SB_T0_SOUTH_SB_OUT_B17;
	input SB_T0_SOUTH_SB_OUT_B17_ready;
	output wire SB_T0_SOUTH_SB_OUT_B17_valid;
	input SB_T0_SOUTH_SB_OUT_B1_ready;
	output wire SB_T0_SOUTH_SB_OUT_B1_valid;
	input [0:0] SB_T0_WEST_SB_IN_B1;
	input [16:0] SB_T0_WEST_SB_IN_B17;
	output wire SB_T0_WEST_SB_IN_B17_ready;
	input SB_T0_WEST_SB_IN_B17_valid;
	output wire SB_T0_WEST_SB_IN_B1_ready;
	input SB_T0_WEST_SB_IN_B1_valid;
	output wire [0:0] SB_T0_WEST_SB_OUT_B1;
	output wire [16:0] SB_T0_WEST_SB_OUT_B17;
	input SB_T0_WEST_SB_OUT_B17_ready;
	output wire SB_T0_WEST_SB_OUT_B17_valid;
	input SB_T0_WEST_SB_OUT_B1_ready;
	output wire SB_T0_WEST_SB_OUT_B1_valid;
	input [0:0] SB_T1_EAST_SB_IN_B1;
	input [16:0] SB_T1_EAST_SB_IN_B17;
	output wire SB_T1_EAST_SB_IN_B17_ready;
	input SB_T1_EAST_SB_IN_B17_valid;
	output wire SB_T1_EAST_SB_IN_B1_ready;
	input SB_T1_EAST_SB_IN_B1_valid;
	output wire [0:0] SB_T1_EAST_SB_OUT_B1;
	output wire [16:0] SB_T1_EAST_SB_OUT_B17;
	input SB_T1_EAST_SB_OUT_B17_ready;
	output wire SB_T1_EAST_SB_OUT_B17_valid;
	input SB_T1_EAST_SB_OUT_B1_ready;
	output wire SB_T1_EAST_SB_OUT_B1_valid;
	input [0:0] SB_T1_NORTH_SB_IN_B1;
	input [16:0] SB_T1_NORTH_SB_IN_B17;
	output wire SB_T1_NORTH_SB_IN_B17_ready;
	input SB_T1_NORTH_SB_IN_B17_valid;
	output wire SB_T1_NORTH_SB_IN_B1_ready;
	input SB_T1_NORTH_SB_IN_B1_valid;
	output wire [0:0] SB_T1_NORTH_SB_OUT_B1;
	output wire [16:0] SB_T1_NORTH_SB_OUT_B17;
	input SB_T1_NORTH_SB_OUT_B17_ready;
	output wire SB_T1_NORTH_SB_OUT_B17_valid;
	input SB_T1_NORTH_SB_OUT_B1_ready;
	output wire SB_T1_NORTH_SB_OUT_B1_valid;
	input [0:0] SB_T1_SOUTH_SB_IN_B1;
	input [16:0] SB_T1_SOUTH_SB_IN_B17;
	output wire SB_T1_SOUTH_SB_IN_B17_ready;
	input SB_T1_SOUTH_SB_IN_B17_valid;
	output wire SB_T1_SOUTH_SB_IN_B1_ready;
	input SB_T1_SOUTH_SB_IN_B1_valid;
	output wire [0:0] SB_T1_SOUTH_SB_OUT_B1;
	output wire [16:0] SB_T1_SOUTH_SB_OUT_B17;
	input SB_T1_SOUTH_SB_OUT_B17_ready;
	output wire SB_T1_SOUTH_SB_OUT_B17_valid;
	input SB_T1_SOUTH_SB_OUT_B1_ready;
	output wire SB_T1_SOUTH_SB_OUT_B1_valid;
	input [0:0] SB_T1_WEST_SB_IN_B1;
	input [16:0] SB_T1_WEST_SB_IN_B17;
	output wire SB_T1_WEST_SB_IN_B17_ready;
	input SB_T1_WEST_SB_IN_B17_valid;
	output wire SB_T1_WEST_SB_IN_B1_ready;
	input SB_T1_WEST_SB_IN_B1_valid;
	output wire [0:0] SB_T1_WEST_SB_OUT_B1;
	output wire [16:0] SB_T1_WEST_SB_OUT_B17;
	input SB_T1_WEST_SB_OUT_B17_ready;
	output wire SB_T1_WEST_SB_OUT_B17_valid;
	input SB_T1_WEST_SB_OUT_B1_ready;
	output wire SB_T1_WEST_SB_OUT_B1_valid;
	input [0:0] SB_T2_EAST_SB_IN_B1;
	input [16:0] SB_T2_EAST_SB_IN_B17;
	output wire SB_T2_EAST_SB_IN_B17_ready;
	input SB_T2_EAST_SB_IN_B17_valid;
	output wire SB_T2_EAST_SB_IN_B1_ready;
	input SB_T2_EAST_SB_IN_B1_valid;
	output wire [0:0] SB_T2_EAST_SB_OUT_B1;
	output wire [16:0] SB_T2_EAST_SB_OUT_B17;
	input SB_T2_EAST_SB_OUT_B17_ready;
	output wire SB_T2_EAST_SB_OUT_B17_valid;
	input SB_T2_EAST_SB_OUT_B1_ready;
	output wire SB_T2_EAST_SB_OUT_B1_valid;
	input [0:0] SB_T2_NORTH_SB_IN_B1;
	input [16:0] SB_T2_NORTH_SB_IN_B17;
	output wire SB_T2_NORTH_SB_IN_B17_ready;
	input SB_T2_NORTH_SB_IN_B17_valid;
	output wire SB_T2_NORTH_SB_IN_B1_ready;
	input SB_T2_NORTH_SB_IN_B1_valid;
	output wire [0:0] SB_T2_NORTH_SB_OUT_B1;
	output wire [16:0] SB_T2_NORTH_SB_OUT_B17;
	input SB_T2_NORTH_SB_OUT_B17_ready;
	output wire SB_T2_NORTH_SB_OUT_B17_valid;
	input SB_T2_NORTH_SB_OUT_B1_ready;
	output wire SB_T2_NORTH_SB_OUT_B1_valid;
	input [0:0] SB_T2_SOUTH_SB_IN_B1;
	input [16:0] SB_T2_SOUTH_SB_IN_B17;
	output wire SB_T2_SOUTH_SB_IN_B17_ready;
	input SB_T2_SOUTH_SB_IN_B17_valid;
	output wire SB_T2_SOUTH_SB_IN_B1_ready;
	input SB_T2_SOUTH_SB_IN_B1_valid;
	output wire [0:0] SB_T2_SOUTH_SB_OUT_B1;
	output wire [16:0] SB_T2_SOUTH_SB_OUT_B17;
	input SB_T2_SOUTH_SB_OUT_B17_ready;
	output wire SB_T2_SOUTH_SB_OUT_B17_valid;
	input SB_T2_SOUTH_SB_OUT_B1_ready;
	output wire SB_T2_SOUTH_SB_OUT_B1_valid;
	input [0:0] SB_T2_WEST_SB_IN_B1;
	input [16:0] SB_T2_WEST_SB_IN_B17;
	output wire SB_T2_WEST_SB_IN_B17_ready;
	input SB_T2_WEST_SB_IN_B17_valid;
	output wire SB_T2_WEST_SB_IN_B1_ready;
	input SB_T2_WEST_SB_IN_B1_valid;
	output wire [0:0] SB_T2_WEST_SB_OUT_B1;
	output wire [16:0] SB_T2_WEST_SB_OUT_B17;
	input SB_T2_WEST_SB_OUT_B17_ready;
	output wire SB_T2_WEST_SB_OUT_B17_valid;
	input SB_T2_WEST_SB_OUT_B1_ready;
	output wire SB_T2_WEST_SB_OUT_B1_valid;
	input [0:0] SB_T3_EAST_SB_IN_B1;
	input [16:0] SB_T3_EAST_SB_IN_B17;
	output wire SB_T3_EAST_SB_IN_B17_ready;
	input SB_T3_EAST_SB_IN_B17_valid;
	output wire SB_T3_EAST_SB_IN_B1_ready;
	input SB_T3_EAST_SB_IN_B1_valid;
	output wire [0:0] SB_T3_EAST_SB_OUT_B1;
	output wire [16:0] SB_T3_EAST_SB_OUT_B17;
	input SB_T3_EAST_SB_OUT_B17_ready;
	output wire SB_T3_EAST_SB_OUT_B17_valid;
	input SB_T3_EAST_SB_OUT_B1_ready;
	output wire SB_T3_EAST_SB_OUT_B1_valid;
	input [0:0] SB_T3_NORTH_SB_IN_B1;
	input [16:0] SB_T3_NORTH_SB_IN_B17;
	output wire SB_T3_NORTH_SB_IN_B17_ready;
	input SB_T3_NORTH_SB_IN_B17_valid;
	output wire SB_T3_NORTH_SB_IN_B1_ready;
	input SB_T3_NORTH_SB_IN_B1_valid;
	output wire [0:0] SB_T3_NORTH_SB_OUT_B1;
	output wire [16:0] SB_T3_NORTH_SB_OUT_B17;
	input SB_T3_NORTH_SB_OUT_B17_ready;
	output wire SB_T3_NORTH_SB_OUT_B17_valid;
	input SB_T3_NORTH_SB_OUT_B1_ready;
	output wire SB_T3_NORTH_SB_OUT_B1_valid;
	input [0:0] SB_T3_SOUTH_SB_IN_B1;
	input [16:0] SB_T3_SOUTH_SB_IN_B17;
	output wire SB_T3_SOUTH_SB_IN_B17_ready;
	input SB_T3_SOUTH_SB_IN_B17_valid;
	output wire SB_T3_SOUTH_SB_IN_B1_ready;
	input SB_T3_SOUTH_SB_IN_B1_valid;
	output wire [0:0] SB_T3_SOUTH_SB_OUT_B1;
	output wire [16:0] SB_T3_SOUTH_SB_OUT_B17;
	input SB_T3_SOUTH_SB_OUT_B17_ready;
	output wire SB_T3_SOUTH_SB_OUT_B17_valid;
	input SB_T3_SOUTH_SB_OUT_B1_ready;
	output wire SB_T3_SOUTH_SB_OUT_B1_valid;
	input [0:0] SB_T3_WEST_SB_IN_B1;
	input [16:0] SB_T3_WEST_SB_IN_B17;
	output wire SB_T3_WEST_SB_IN_B17_ready;
	input SB_T3_WEST_SB_IN_B17_valid;
	output wire SB_T3_WEST_SB_IN_B1_ready;
	input SB_T3_WEST_SB_IN_B1_valid;
	output wire [0:0] SB_T3_WEST_SB_OUT_B1;
	output wire [16:0] SB_T3_WEST_SB_OUT_B17;
	input SB_T3_WEST_SB_OUT_B17_ready;
	output wire SB_T3_WEST_SB_OUT_B17_valid;
	input SB_T3_WEST_SB_OUT_B1_ready;
	output wire SB_T3_WEST_SB_OUT_B1_valid;
	input [0:0] SB_T4_EAST_SB_IN_B1;
	input [16:0] SB_T4_EAST_SB_IN_B17;
	output wire SB_T4_EAST_SB_IN_B17_ready;
	input SB_T4_EAST_SB_IN_B17_valid;
	output wire SB_T4_EAST_SB_IN_B1_ready;
	input SB_T4_EAST_SB_IN_B1_valid;
	output wire [0:0] SB_T4_EAST_SB_OUT_B1;
	output wire [16:0] SB_T4_EAST_SB_OUT_B17;
	input SB_T4_EAST_SB_OUT_B17_ready;
	output wire SB_T4_EAST_SB_OUT_B17_valid;
	input SB_T4_EAST_SB_OUT_B1_ready;
	output wire SB_T4_EAST_SB_OUT_B1_valid;
	input [0:0] SB_T4_NORTH_SB_IN_B1;
	input [16:0] SB_T4_NORTH_SB_IN_B17;
	output wire SB_T4_NORTH_SB_IN_B17_ready;
	input SB_T4_NORTH_SB_IN_B17_valid;
	output wire SB_T4_NORTH_SB_IN_B1_ready;
	input SB_T4_NORTH_SB_IN_B1_valid;
	output wire [0:0] SB_T4_NORTH_SB_OUT_B1;
	output wire [16:0] SB_T4_NORTH_SB_OUT_B17;
	input SB_T4_NORTH_SB_OUT_B17_ready;
	output wire SB_T4_NORTH_SB_OUT_B17_valid;
	input SB_T4_NORTH_SB_OUT_B1_ready;
	output wire SB_T4_NORTH_SB_OUT_B1_valid;
	input [0:0] SB_T4_SOUTH_SB_IN_B1;
	input [16:0] SB_T4_SOUTH_SB_IN_B17;
	output wire SB_T4_SOUTH_SB_IN_B17_ready;
	input SB_T4_SOUTH_SB_IN_B17_valid;
	output wire SB_T4_SOUTH_SB_IN_B1_ready;
	input SB_T4_SOUTH_SB_IN_B1_valid;
	output wire [0:0] SB_T4_SOUTH_SB_OUT_B1;
	output wire [16:0] SB_T4_SOUTH_SB_OUT_B17;
	input SB_T4_SOUTH_SB_OUT_B17_ready;
	output wire SB_T4_SOUTH_SB_OUT_B17_valid;
	input SB_T4_SOUTH_SB_OUT_B1_ready;
	output wire SB_T4_SOUTH_SB_OUT_B1_valid;
	input [0:0] SB_T4_WEST_SB_IN_B1;
	input [16:0] SB_T4_WEST_SB_IN_B17;
	output wire SB_T4_WEST_SB_IN_B17_ready;
	input SB_T4_WEST_SB_IN_B17_valid;
	output wire SB_T4_WEST_SB_IN_B1_ready;
	input SB_T4_WEST_SB_IN_B1_valid;
	output wire [0:0] SB_T4_WEST_SB_OUT_B1;
	output wire [16:0] SB_T4_WEST_SB_OUT_B17;
	input SB_T4_WEST_SB_OUT_B17_ready;
	output wire SB_T4_WEST_SB_OUT_B17_valid;
	input SB_T4_WEST_SB_OUT_B1_ready;
	output wire SB_T4_WEST_SB_OUT_B1_valid;
	input clk;
	output wire clk_out;
	input [31:0] config_config_addr;
	input [31:0] config_config_data;
	output wire [31:0] config_out_config_addr;
	output wire [31:0] config_out_config_data;
	output wire [0:0] config_out_read;
	output wire [0:0] config_out_write;
	input [0:0] config_read;
	input [0:0] config_write;
	input [0:0] flush;
	output wire [0:0] flush_out;
	output wire [8:0] hi;
	output wire [7:0] lo;
	output wire [31:0] read_config_data;
	input [31:0] read_config_data_in;
	input reset;
	output wire reset_out;
	input [0:0] stall;
	output wire [0:0] stall_out;
	input [15:0] tile_id;
	wire [16:0] CB_MEM_input_width_17_num_0_O;
	wire CB_MEM_input_width_17_num_0_enable;
	wire [31:0] CB_MEM_input_width_17_num_0_out_sel;
	wire [31:0] CB_MEM_input_width_17_num_0_read_config_data;
	wire CB_MEM_input_width_17_num_0_ready_out;
	wire CB_MEM_input_width_17_num_0_valid_out;
	wire [16:0] CB_MEM_input_width_17_num_1_O;
	wire CB_MEM_input_width_17_num_1_enable;
	wire [31:0] CB_MEM_input_width_17_num_1_out_sel;
	wire [31:0] CB_MEM_input_width_17_num_1_read_config_data;
	wire CB_MEM_input_width_17_num_1_ready_out;
	wire CB_MEM_input_width_17_num_1_valid_out;
	wire [16:0] CB_MEM_input_width_17_num_2_O;
	wire CB_MEM_input_width_17_num_2_enable;
	wire [31:0] CB_MEM_input_width_17_num_2_out_sel;
	wire [31:0] CB_MEM_input_width_17_num_2_read_config_data;
	wire CB_MEM_input_width_17_num_2_ready_out;
	wire CB_MEM_input_width_17_num_2_valid_out;
	wire [16:0] CB_MEM_input_width_17_num_3_O;
	wire CB_MEM_input_width_17_num_3_enable;
	wire [31:0] CB_MEM_input_width_17_num_3_out_sel;
	wire [31:0] CB_MEM_input_width_17_num_3_read_config_data;
	wire CB_MEM_input_width_17_num_3_ready_out;
	wire CB_MEM_input_width_17_num_3_valid_out;
	wire [0:0] CB_MEM_input_width_1_num_0_O;
	wire CB_MEM_input_width_1_num_0_enable;
	wire [31:0] CB_MEM_input_width_1_num_0_out_sel;
	wire [31:0] CB_MEM_input_width_1_num_0_read_config_data;
	wire CB_MEM_input_width_1_num_0_ready_out;
	wire CB_MEM_input_width_1_num_0_valid_out;
	wire [0:0] CB_MEM_input_width_1_num_1_O;
	wire CB_MEM_input_width_1_num_1_enable;
	wire [31:0] CB_MEM_input_width_1_num_1_out_sel;
	wire [31:0] CB_MEM_input_width_1_num_1_read_config_data;
	wire CB_MEM_input_width_1_num_1_ready_out;
	wire CB_MEM_input_width_1_num_1_valid_out;
	wire [0:0] CB_flush_O;
	wire CB_flush_enable;
	wire [31:0] CB_flush_out_sel;
	wire [31:0] CB_flush_read_config_data;
	wire CB_flush_ready_out;
	wire CB_flush_valid_out;
	wire DECODE_FEATURE_0_O;
	wire DECODE_FEATURE_1_O;
	wire DECODE_FEATURE_10_O;
	wire DECODE_FEATURE_11_O;
	wire DECODE_FEATURE_12_O;
	wire DECODE_FEATURE_2_O;
	wire DECODE_FEATURE_3_O;
	wire DECODE_FEATURE_4_O;
	wire DECODE_FEATURE_5_O;
	wire DECODE_FEATURE_6_O;
	wire DECODE_FEATURE_7_O;
	wire DECODE_FEATURE_8_O;
	wire DECODE_FEATURE_9_O;
	wire FEATURE_AND_0_out;
	wire FEATURE_AND_1_out;
	wire FEATURE_AND_10_out;
	wire FEATURE_AND_11_out;
	wire FEATURE_AND_12_out;
	wire FEATURE_AND_2_out;
	wire FEATURE_AND_3_out;
	wire FEATURE_AND_4_out;
	wire FEATURE_AND_5_out;
	wire FEATURE_AND_6_out;
	wire FEATURE_AND_7_out;
	wire FEATURE_AND_8_out;
	wire FEATURE_AND_9_out;
	wire [0:0] MEM_output_width_17_num_0_loopback_valid_out;
	wire [0:0] MEM_output_width_17_num_1_loopback_valid_out;
	wire [0:0] MEM_output_width_17_num_2_loopback_valid_out;
	wire [0:0] MEM_output_width_1_num_0_loopback_valid_out;
	wire [0:0] MEM_output_width_1_num_1_loopback_valid_out;
	wire [0:0] MEM_output_width_1_num_2_loopback_valid_out;
	wire [0:0] MemCore_inst0_MEM_input_width_17_num_0_ready;
	wire [0:0] MemCore_inst0_MEM_input_width_17_num_1_ready;
	wire [0:0] MemCore_inst0_MEM_input_width_17_num_2_ready;
	wire [0:0] MemCore_inst0_MEM_input_width_17_num_3_ready;
	wire MemCore_inst0_MEM_input_width_1_num_0_ready;
	wire MemCore_inst0_MEM_input_width_1_num_1_ready;
	wire [16:0] MemCore_inst0_MEM_output_width_17_num_0;
	wire [0:0] MemCore_inst0_MEM_output_width_17_num_0_valid;
	wire [16:0] MemCore_inst0_MEM_output_width_17_num_1;
	wire [0:0] MemCore_inst0_MEM_output_width_17_num_1_valid;
	wire [16:0] MemCore_inst0_MEM_output_width_17_num_2;
	wire [0:0] MemCore_inst0_MEM_output_width_17_num_2_valid;
	wire [0:0] MemCore_inst0_MEM_output_width_1_num_0;
	wire MemCore_inst0_MEM_output_width_1_num_0_valid;
	wire [0:0] MemCore_inst0_MEM_output_width_1_num_1;
	wire MemCore_inst0_MEM_output_width_1_num_1_valid;
	wire [0:0] MemCore_inst0_MEM_output_width_1_num_2;
	wire MemCore_inst0_MEM_output_width_1_num_2_valid;
	wire [31:0] MemCore_inst0_read_config_data;
	wire [31:0] MemCore_inst0_read_config_data_1;
	wire [31:0] MemCore_inst0_read_config_data_2;
	wire [0:0] PowerDomainConfigReg_inst0_ps_en_out;
	wire [31:0] PowerDomainConfigReg_inst0_read_config_data;
	wire [31:0] PowerDomainOR_O;
	wire SB_ID0_5TRACKS_B17_MemCore_MEM_output_width_17_num_0_ready_out;
	wire SB_ID0_5TRACKS_B17_MemCore_MEM_output_width_17_num_1_ready_out;
	wire SB_ID0_5TRACKS_B17_MemCore_MEM_output_width_17_num_2_ready_out;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_EAST_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_EAST_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T0_EAST_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_EAST_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_EAST_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_NORTH_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_NORTH_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T0_NORTH_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_NORTH_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_NORTH_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_SOUTH_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_SOUTH_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T0_SOUTH_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_SOUTH_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_SOUTH_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_WEST_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_WEST_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T0_WEST_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_WEST_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_WEST_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_EAST_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_EAST_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T1_EAST_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_EAST_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_EAST_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_NORTH_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_NORTH_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T1_NORTH_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_NORTH_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_NORTH_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_SOUTH_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_SOUTH_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T1_SOUTH_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_SOUTH_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_SOUTH_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_WEST_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_WEST_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T1_WEST_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_WEST_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_WEST_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_EAST_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_EAST_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T2_EAST_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_EAST_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_EAST_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_NORTH_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_NORTH_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T2_NORTH_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_NORTH_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_NORTH_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_SOUTH_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_SOUTH_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T2_SOUTH_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_SOUTH_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_SOUTH_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_WEST_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_WEST_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T2_WEST_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_WEST_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_WEST_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_EAST_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_EAST_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T3_EAST_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_EAST_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_EAST_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_NORTH_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_NORTH_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T3_NORTH_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_NORTH_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_NORTH_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_SOUTH_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_SOUTH_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T3_SOUTH_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_SOUTH_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_SOUTH_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_WEST_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_WEST_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T3_WEST_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_WEST_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_WEST_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_EAST_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_EAST_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T4_EAST_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_EAST_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_EAST_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_NORTH_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_NORTH_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T4_NORTH_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_NORTH_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_NORTH_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_SOUTH_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_SOUTH_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T4_SOUTH_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_SOUTH_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_SOUTH_SB_OUT_B17_valid_out;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_WEST_SB_IN_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_WEST_SB_IN_B17_ready_out;
	wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T4_WEST_SB_OUT_B17;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_WEST_SB_OUT_B17_enable;
	wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_WEST_SB_OUT_B17_valid_out;
	wire [31:0] SB_ID0_5TRACKS_B17_MemCore_read_config_data;
	wire SB_ID0_5TRACKS_B1_MemCore_MEM_output_width_1_num_0_ready_out;
	wire SB_ID0_5TRACKS_B1_MemCore_MEM_output_width_1_num_1_ready_out;
	wire SB_ID0_5TRACKS_B1_MemCore_MEM_output_width_1_num_2_ready_out;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_OUT_B1_valid_out;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_IN_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_IN_B1_ready_out;
	wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_OUT_B1;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_OUT_B1_enable;
	wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_OUT_B1_valid_out;
	wire [31:0] SB_ID0_5TRACKS_B1_MemCore_read_config_data;
	wire SB_T0_EAST_SB_OUT_B17_ready_and_Z;
	wire SB_T0_EAST_SB_OUT_B1_ready_and_Z;
	wire SB_T0_NORTH_SB_OUT_B17_ready_and_Z;
	wire SB_T0_NORTH_SB_OUT_B1_ready_and_Z;
	wire SB_T0_SOUTH_SB_OUT_B17_ready_and_Z;
	wire SB_T0_SOUTH_SB_OUT_B1_ready_and_Z;
	wire SB_T0_WEST_SB_OUT_B17_ready_and_Z;
	wire SB_T0_WEST_SB_OUT_B1_ready_and_Z;
	wire SB_T1_EAST_SB_OUT_B17_ready_and_Z;
	wire SB_T1_EAST_SB_OUT_B1_ready_and_Z;
	wire SB_T1_NORTH_SB_OUT_B17_ready_and_Z;
	wire SB_T1_NORTH_SB_OUT_B1_ready_and_Z;
	wire SB_T1_SOUTH_SB_OUT_B17_ready_and_Z;
	wire SB_T1_SOUTH_SB_OUT_B1_ready_and_Z;
	wire SB_T1_WEST_SB_OUT_B17_ready_and_Z;
	wire SB_T1_WEST_SB_OUT_B1_ready_and_Z;
	wire SB_T2_EAST_SB_OUT_B17_ready_and_Z;
	wire SB_T2_EAST_SB_OUT_B1_ready_and_Z;
	wire SB_T2_NORTH_SB_OUT_B17_ready_and_Z;
	wire SB_T2_NORTH_SB_OUT_B1_ready_and_Z;
	wire SB_T2_SOUTH_SB_OUT_B17_ready_and_Z;
	wire SB_T2_SOUTH_SB_OUT_B1_ready_and_Z;
	wire SB_T2_WEST_SB_OUT_B17_ready_and_Z;
	wire SB_T2_WEST_SB_OUT_B1_ready_and_Z;
	wire SB_T3_EAST_SB_OUT_B17_ready_and_Z;
	wire SB_T3_EAST_SB_OUT_B1_ready_and_Z;
	wire SB_T3_NORTH_SB_OUT_B17_ready_and_Z;
	wire SB_T3_NORTH_SB_OUT_B1_ready_and_Z;
	wire SB_T3_SOUTH_SB_OUT_B17_ready_and_Z;
	wire SB_T3_SOUTH_SB_OUT_B1_ready_and_Z;
	wire SB_T3_WEST_SB_OUT_B17_ready_and_Z;
	wire SB_T3_WEST_SB_OUT_B1_ready_and_Z;
	wire SB_T4_EAST_SB_OUT_B17_ready_and_Z;
	wire SB_T4_EAST_SB_OUT_B1_ready_and_Z;
	wire SB_T4_NORTH_SB_OUT_B17_ready_and_Z;
	wire SB_T4_NORTH_SB_OUT_B1_ready_and_Z;
	wire SB_T4_SOUTH_SB_OUT_B17_ready_and_Z;
	wire SB_T4_SOUTH_SB_OUT_B1_ready_and_Z;
	wire SB_T4_WEST_SB_OUT_B17_ready_and_Z;
	wire SB_T4_WEST_SB_OUT_B1_ready_and_Z;
	wire and_inst0_out;
	wire and_inst1_out;
	wire bit_const_1_None_out;
	wire [7:0] const_0_8_out;
	wire [8:0] const_511_9_out;
	wire coreir_eq_16_inst0_out;
	wire [31:0] read_data_mux_O;
	wire [31:0] self_config_config_addr_out;
	wire [339:0] CB_MEM_input_width_17_num_0_I;
	assign CB_MEM_input_width_17_num_0_I[323+:17] = SB_T4_WEST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_0_I[306+:17] = SB_T4_EAST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_0_I[289+:17] = SB_T4_SOUTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_0_I[272+:17] = SB_T4_NORTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_0_I[255+:17] = SB_T3_WEST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_0_I[238+:17] = SB_T3_EAST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_0_I[221+:17] = SB_T3_SOUTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_0_I[204+:17] = SB_T3_NORTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_0_I[187+:17] = SB_T2_WEST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_0_I[170+:17] = SB_T2_EAST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_0_I[153+:17] = SB_T2_SOUTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_0_I[136+:17] = SB_T2_NORTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_0_I[119+:17] = SB_T1_WEST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_0_I[102+:17] = SB_T1_EAST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_0_I[85+:17] = SB_T1_SOUTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_0_I[68+:17] = SB_T1_NORTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_0_I[51+:17] = SB_T0_WEST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_0_I[34+:17] = SB_T0_EAST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_0_I[17+:17] = SB_T0_SOUTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_0_I[0+:17] = SB_T0_NORTH_SB_IN_B17;
	wire [19:0] CB_MEM_input_width_17_num_0_valid_in;
	assign CB_MEM_input_width_17_num_0_valid_in = {SB_T4_WEST_SB_IN_B17_valid, SB_T4_EAST_SB_IN_B17_valid, SB_T4_SOUTH_SB_IN_B17_valid, SB_T4_NORTH_SB_IN_B17_valid, SB_T3_WEST_SB_IN_B17_valid, SB_T3_EAST_SB_IN_B17_valid, SB_T3_SOUTH_SB_IN_B17_valid, SB_T3_NORTH_SB_IN_B17_valid, SB_T2_WEST_SB_IN_B17_valid, SB_T2_EAST_SB_IN_B17_valid, SB_T2_SOUTH_SB_IN_B17_valid, SB_T2_NORTH_SB_IN_B17_valid, SB_T1_WEST_SB_IN_B17_valid, SB_T1_EAST_SB_IN_B17_valid, SB_T1_SOUTH_SB_IN_B17_valid, SB_T1_NORTH_SB_IN_B17_valid, SB_T0_WEST_SB_IN_B17_valid, SB_T0_EAST_SB_IN_B17_valid, SB_T0_SOUTH_SB_IN_B17_valid, SB_T0_NORTH_SB_IN_B17_valid};
	CB_MEM_input_width_17_num_0 CB_MEM_input_width_17_num_0(
		.I(CB_MEM_input_width_17_num_0_I),
		.O(CB_MEM_input_width_17_num_0_O),
		.clk(clk),
		.config_config_addr(self_config_config_addr_out[31:24]),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_3_out),
		.enable(CB_MEM_input_width_17_num_0_enable),
		.out_sel(CB_MEM_input_width_17_num_0_out_sel),
		.read_config_data(CB_MEM_input_width_17_num_0_read_config_data),
		.ready_in(MemCore_inst0_MEM_input_width_17_num_0_ready[0]),
		.ready_out(CB_MEM_input_width_17_num_0_ready_out),
		.reset(reset),
		.valid_in(CB_MEM_input_width_17_num_0_valid_in),
		.valid_out(CB_MEM_input_width_17_num_0_valid_out)
	);
	wire [339:0] CB_MEM_input_width_17_num_1_I;
	assign CB_MEM_input_width_17_num_1_I[323+:17] = SB_T4_WEST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_1_I[306+:17] = SB_T4_EAST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_1_I[289+:17] = SB_T4_SOUTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_1_I[272+:17] = SB_T4_NORTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_1_I[255+:17] = SB_T3_WEST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_1_I[238+:17] = SB_T3_EAST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_1_I[221+:17] = SB_T3_SOUTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_1_I[204+:17] = SB_T3_NORTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_1_I[187+:17] = SB_T2_WEST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_1_I[170+:17] = SB_T2_EAST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_1_I[153+:17] = SB_T2_SOUTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_1_I[136+:17] = SB_T2_NORTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_1_I[119+:17] = SB_T1_WEST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_1_I[102+:17] = SB_T1_EAST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_1_I[85+:17] = SB_T1_SOUTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_1_I[68+:17] = SB_T1_NORTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_1_I[51+:17] = SB_T0_WEST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_1_I[34+:17] = SB_T0_EAST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_1_I[17+:17] = SB_T0_SOUTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_1_I[0+:17] = SB_T0_NORTH_SB_IN_B17;
	wire [19:0] CB_MEM_input_width_17_num_1_valid_in;
	assign CB_MEM_input_width_17_num_1_valid_in = {SB_T4_WEST_SB_IN_B17_valid, SB_T4_EAST_SB_IN_B17_valid, SB_T4_SOUTH_SB_IN_B17_valid, SB_T4_NORTH_SB_IN_B17_valid, SB_T3_WEST_SB_IN_B17_valid, SB_T3_EAST_SB_IN_B17_valid, SB_T3_SOUTH_SB_IN_B17_valid, SB_T3_NORTH_SB_IN_B17_valid, SB_T2_WEST_SB_IN_B17_valid, SB_T2_EAST_SB_IN_B17_valid, SB_T2_SOUTH_SB_IN_B17_valid, SB_T2_NORTH_SB_IN_B17_valid, SB_T1_WEST_SB_IN_B17_valid, SB_T1_EAST_SB_IN_B17_valid, SB_T1_SOUTH_SB_IN_B17_valid, SB_T1_NORTH_SB_IN_B17_valid, SB_T0_WEST_SB_IN_B17_valid, SB_T0_EAST_SB_IN_B17_valid, SB_T0_SOUTH_SB_IN_B17_valid, SB_T0_NORTH_SB_IN_B17_valid};
	CB_MEM_input_width_17_num_1 CB_MEM_input_width_17_num_1(
		.I(CB_MEM_input_width_17_num_1_I),
		.O(CB_MEM_input_width_17_num_1_O),
		.clk(clk),
		.config_config_addr(self_config_config_addr_out[31:24]),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_4_out),
		.enable(CB_MEM_input_width_17_num_1_enable),
		.out_sel(CB_MEM_input_width_17_num_1_out_sel),
		.read_config_data(CB_MEM_input_width_17_num_1_read_config_data),
		.ready_in(MemCore_inst0_MEM_input_width_17_num_1_ready[0]),
		.ready_out(CB_MEM_input_width_17_num_1_ready_out),
		.reset(reset),
		.valid_in(CB_MEM_input_width_17_num_1_valid_in),
		.valid_out(CB_MEM_input_width_17_num_1_valid_out)
	);
	wire [339:0] CB_MEM_input_width_17_num_2_I;
	assign CB_MEM_input_width_17_num_2_I[323+:17] = SB_T4_WEST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_2_I[306+:17] = SB_T4_EAST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_2_I[289+:17] = SB_T4_SOUTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_2_I[272+:17] = SB_T4_NORTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_2_I[255+:17] = SB_T3_WEST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_2_I[238+:17] = SB_T3_EAST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_2_I[221+:17] = SB_T3_SOUTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_2_I[204+:17] = SB_T3_NORTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_2_I[187+:17] = SB_T2_WEST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_2_I[170+:17] = SB_T2_EAST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_2_I[153+:17] = SB_T2_SOUTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_2_I[136+:17] = SB_T2_NORTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_2_I[119+:17] = SB_T1_WEST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_2_I[102+:17] = SB_T1_EAST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_2_I[85+:17] = SB_T1_SOUTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_2_I[68+:17] = SB_T1_NORTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_2_I[51+:17] = SB_T0_WEST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_2_I[34+:17] = SB_T0_EAST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_2_I[17+:17] = SB_T0_SOUTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_2_I[0+:17] = SB_T0_NORTH_SB_IN_B17;
	wire [19:0] CB_MEM_input_width_17_num_2_valid_in;
	assign CB_MEM_input_width_17_num_2_valid_in = {SB_T4_WEST_SB_IN_B17_valid, SB_T4_EAST_SB_IN_B17_valid, SB_T4_SOUTH_SB_IN_B17_valid, SB_T4_NORTH_SB_IN_B17_valid, SB_T3_WEST_SB_IN_B17_valid, SB_T3_EAST_SB_IN_B17_valid, SB_T3_SOUTH_SB_IN_B17_valid, SB_T3_NORTH_SB_IN_B17_valid, SB_T2_WEST_SB_IN_B17_valid, SB_T2_EAST_SB_IN_B17_valid, SB_T2_SOUTH_SB_IN_B17_valid, SB_T2_NORTH_SB_IN_B17_valid, SB_T1_WEST_SB_IN_B17_valid, SB_T1_EAST_SB_IN_B17_valid, SB_T1_SOUTH_SB_IN_B17_valid, SB_T1_NORTH_SB_IN_B17_valid, SB_T0_WEST_SB_IN_B17_valid, SB_T0_EAST_SB_IN_B17_valid, SB_T0_SOUTH_SB_IN_B17_valid, SB_T0_NORTH_SB_IN_B17_valid};
	CB_MEM_input_width_17_num_2 CB_MEM_input_width_17_num_2(
		.I(CB_MEM_input_width_17_num_2_I),
		.O(CB_MEM_input_width_17_num_2_O),
		.clk(clk),
		.config_config_addr(self_config_config_addr_out[31:24]),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_5_out),
		.enable(CB_MEM_input_width_17_num_2_enable),
		.out_sel(CB_MEM_input_width_17_num_2_out_sel),
		.read_config_data(CB_MEM_input_width_17_num_2_read_config_data),
		.ready_in(MemCore_inst0_MEM_input_width_17_num_2_ready[0]),
		.ready_out(CB_MEM_input_width_17_num_2_ready_out),
		.reset(reset),
		.valid_in(CB_MEM_input_width_17_num_2_valid_in),
		.valid_out(CB_MEM_input_width_17_num_2_valid_out)
	);
	wire [339:0] CB_MEM_input_width_17_num_3_I;
	assign CB_MEM_input_width_17_num_3_I[323+:17] = SB_T4_WEST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_3_I[306+:17] = SB_T4_EAST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_3_I[289+:17] = SB_T4_SOUTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_3_I[272+:17] = SB_T4_NORTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_3_I[255+:17] = SB_T3_WEST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_3_I[238+:17] = SB_T3_EAST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_3_I[221+:17] = SB_T3_SOUTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_3_I[204+:17] = SB_T3_NORTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_3_I[187+:17] = SB_T2_WEST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_3_I[170+:17] = SB_T2_EAST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_3_I[153+:17] = SB_T2_SOUTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_3_I[136+:17] = SB_T2_NORTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_3_I[119+:17] = SB_T1_WEST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_3_I[102+:17] = SB_T1_EAST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_3_I[85+:17] = SB_T1_SOUTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_3_I[68+:17] = SB_T1_NORTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_3_I[51+:17] = SB_T0_WEST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_3_I[34+:17] = SB_T0_EAST_SB_IN_B17;
	assign CB_MEM_input_width_17_num_3_I[17+:17] = SB_T0_SOUTH_SB_IN_B17;
	assign CB_MEM_input_width_17_num_3_I[0+:17] = SB_T0_NORTH_SB_IN_B17;
	wire [19:0] CB_MEM_input_width_17_num_3_valid_in;
	assign CB_MEM_input_width_17_num_3_valid_in = {SB_T4_WEST_SB_IN_B17_valid, SB_T4_EAST_SB_IN_B17_valid, SB_T4_SOUTH_SB_IN_B17_valid, SB_T4_NORTH_SB_IN_B17_valid, SB_T3_WEST_SB_IN_B17_valid, SB_T3_EAST_SB_IN_B17_valid, SB_T3_SOUTH_SB_IN_B17_valid, SB_T3_NORTH_SB_IN_B17_valid, SB_T2_WEST_SB_IN_B17_valid, SB_T2_EAST_SB_IN_B17_valid, SB_T2_SOUTH_SB_IN_B17_valid, SB_T2_NORTH_SB_IN_B17_valid, SB_T1_WEST_SB_IN_B17_valid, SB_T1_EAST_SB_IN_B17_valid, SB_T1_SOUTH_SB_IN_B17_valid, SB_T1_NORTH_SB_IN_B17_valid, SB_T0_WEST_SB_IN_B17_valid, SB_T0_EAST_SB_IN_B17_valid, SB_T0_SOUTH_SB_IN_B17_valid, SB_T0_NORTH_SB_IN_B17_valid};
	CB_MEM_input_width_17_num_3 CB_MEM_input_width_17_num_3(
		.I(CB_MEM_input_width_17_num_3_I),
		.O(CB_MEM_input_width_17_num_3_O),
		.clk(clk),
		.config_config_addr(self_config_config_addr_out[31:24]),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_6_out),
		.enable(CB_MEM_input_width_17_num_3_enable),
		.out_sel(CB_MEM_input_width_17_num_3_out_sel),
		.read_config_data(CB_MEM_input_width_17_num_3_read_config_data),
		.ready_in(MemCore_inst0_MEM_input_width_17_num_3_ready[0]),
		.ready_out(CB_MEM_input_width_17_num_3_ready_out),
		.reset(reset),
		.valid_in(CB_MEM_input_width_17_num_3_valid_in),
		.valid_out(CB_MEM_input_width_17_num_3_valid_out)
	);
	wire [19:0] CB_MEM_input_width_1_num_0_I;
	assign CB_MEM_input_width_1_num_0_I[19+:1] = SB_T4_WEST_SB_IN_B1;
	assign CB_MEM_input_width_1_num_0_I[18+:1] = SB_T4_EAST_SB_IN_B1;
	assign CB_MEM_input_width_1_num_0_I[17+:1] = SB_T4_SOUTH_SB_IN_B1;
	assign CB_MEM_input_width_1_num_0_I[16+:1] = SB_T4_NORTH_SB_IN_B1;
	assign CB_MEM_input_width_1_num_0_I[15+:1] = SB_T3_WEST_SB_IN_B1;
	assign CB_MEM_input_width_1_num_0_I[14+:1] = SB_T3_EAST_SB_IN_B1;
	assign CB_MEM_input_width_1_num_0_I[13+:1] = SB_T3_SOUTH_SB_IN_B1;
	assign CB_MEM_input_width_1_num_0_I[12+:1] = SB_T3_NORTH_SB_IN_B1;
	assign CB_MEM_input_width_1_num_0_I[11+:1] = SB_T2_WEST_SB_IN_B1;
	assign CB_MEM_input_width_1_num_0_I[10+:1] = SB_T2_EAST_SB_IN_B1;
	assign CB_MEM_input_width_1_num_0_I[9+:1] = SB_T2_SOUTH_SB_IN_B1;
	assign CB_MEM_input_width_1_num_0_I[8+:1] = SB_T2_NORTH_SB_IN_B1;
	assign CB_MEM_input_width_1_num_0_I[7+:1] = SB_T1_WEST_SB_IN_B1;
	assign CB_MEM_input_width_1_num_0_I[6+:1] = SB_T1_EAST_SB_IN_B1;
	assign CB_MEM_input_width_1_num_0_I[5+:1] = SB_T1_SOUTH_SB_IN_B1;
	assign CB_MEM_input_width_1_num_0_I[4+:1] = SB_T1_NORTH_SB_IN_B1;
	assign CB_MEM_input_width_1_num_0_I[3+:1] = SB_T0_WEST_SB_IN_B1;
	assign CB_MEM_input_width_1_num_0_I[2+:1] = SB_T0_EAST_SB_IN_B1;
	assign CB_MEM_input_width_1_num_0_I[1+:1] = SB_T0_SOUTH_SB_IN_B1;
	assign CB_MEM_input_width_1_num_0_I[0+:1] = SB_T0_NORTH_SB_IN_B1;
	wire [19:0] CB_MEM_input_width_1_num_0_valid_in;
	assign CB_MEM_input_width_1_num_0_valid_in = {SB_T4_WEST_SB_IN_B1_valid, SB_T4_EAST_SB_IN_B1_valid, SB_T4_SOUTH_SB_IN_B1_valid, SB_T4_NORTH_SB_IN_B1_valid, SB_T3_WEST_SB_IN_B1_valid, SB_T3_EAST_SB_IN_B1_valid, SB_T3_SOUTH_SB_IN_B1_valid, SB_T3_NORTH_SB_IN_B1_valid, SB_T2_WEST_SB_IN_B1_valid, SB_T2_EAST_SB_IN_B1_valid, SB_T2_SOUTH_SB_IN_B1_valid, SB_T2_NORTH_SB_IN_B1_valid, SB_T1_WEST_SB_IN_B1_valid, SB_T1_EAST_SB_IN_B1_valid, SB_T1_SOUTH_SB_IN_B1_valid, SB_T1_NORTH_SB_IN_B1_valid, SB_T0_WEST_SB_IN_B1_valid, SB_T0_EAST_SB_IN_B1_valid, SB_T0_SOUTH_SB_IN_B1_valid, SB_T0_NORTH_SB_IN_B1_valid};
	CB_MEM_input_width_1_num_0 CB_MEM_input_width_1_num_0(
		.I(CB_MEM_input_width_1_num_0_I),
		.O(CB_MEM_input_width_1_num_0_O),
		.clk(clk),
		.config_config_addr(self_config_config_addr_out[31:24]),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_7_out),
		.enable(CB_MEM_input_width_1_num_0_enable),
		.out_sel(CB_MEM_input_width_1_num_0_out_sel),
		.read_config_data(CB_MEM_input_width_1_num_0_read_config_data),
		.ready_in(MemCore_inst0_MEM_input_width_1_num_0_ready),
		.ready_out(CB_MEM_input_width_1_num_0_ready_out),
		.reset(reset),
		.valid_in(CB_MEM_input_width_1_num_0_valid_in),
		.valid_out(CB_MEM_input_width_1_num_0_valid_out)
	);
	wire [19:0] CB_MEM_input_width_1_num_1_I;
	assign CB_MEM_input_width_1_num_1_I[19+:1] = SB_T4_WEST_SB_IN_B1;
	assign CB_MEM_input_width_1_num_1_I[18+:1] = SB_T4_EAST_SB_IN_B1;
	assign CB_MEM_input_width_1_num_1_I[17+:1] = SB_T4_SOUTH_SB_IN_B1;
	assign CB_MEM_input_width_1_num_1_I[16+:1] = SB_T4_NORTH_SB_IN_B1;
	assign CB_MEM_input_width_1_num_1_I[15+:1] = SB_T3_WEST_SB_IN_B1;
	assign CB_MEM_input_width_1_num_1_I[14+:1] = SB_T3_EAST_SB_IN_B1;
	assign CB_MEM_input_width_1_num_1_I[13+:1] = SB_T3_SOUTH_SB_IN_B1;
	assign CB_MEM_input_width_1_num_1_I[12+:1] = SB_T3_NORTH_SB_IN_B1;
	assign CB_MEM_input_width_1_num_1_I[11+:1] = SB_T2_WEST_SB_IN_B1;
	assign CB_MEM_input_width_1_num_1_I[10+:1] = SB_T2_EAST_SB_IN_B1;
	assign CB_MEM_input_width_1_num_1_I[9+:1] = SB_T2_SOUTH_SB_IN_B1;
	assign CB_MEM_input_width_1_num_1_I[8+:1] = SB_T2_NORTH_SB_IN_B1;
	assign CB_MEM_input_width_1_num_1_I[7+:1] = SB_T1_WEST_SB_IN_B1;
	assign CB_MEM_input_width_1_num_1_I[6+:1] = SB_T1_EAST_SB_IN_B1;
	assign CB_MEM_input_width_1_num_1_I[5+:1] = SB_T1_SOUTH_SB_IN_B1;
	assign CB_MEM_input_width_1_num_1_I[4+:1] = SB_T1_NORTH_SB_IN_B1;
	assign CB_MEM_input_width_1_num_1_I[3+:1] = SB_T0_WEST_SB_IN_B1;
	assign CB_MEM_input_width_1_num_1_I[2+:1] = SB_T0_EAST_SB_IN_B1;
	assign CB_MEM_input_width_1_num_1_I[1+:1] = SB_T0_SOUTH_SB_IN_B1;
	assign CB_MEM_input_width_1_num_1_I[0+:1] = SB_T0_NORTH_SB_IN_B1;
	wire [19:0] CB_MEM_input_width_1_num_1_valid_in;
	assign CB_MEM_input_width_1_num_1_valid_in = {SB_T4_WEST_SB_IN_B1_valid, SB_T4_EAST_SB_IN_B1_valid, SB_T4_SOUTH_SB_IN_B1_valid, SB_T4_NORTH_SB_IN_B1_valid, SB_T3_WEST_SB_IN_B1_valid, SB_T3_EAST_SB_IN_B1_valid, SB_T3_SOUTH_SB_IN_B1_valid, SB_T3_NORTH_SB_IN_B1_valid, SB_T2_WEST_SB_IN_B1_valid, SB_T2_EAST_SB_IN_B1_valid, SB_T2_SOUTH_SB_IN_B1_valid, SB_T2_NORTH_SB_IN_B1_valid, SB_T1_WEST_SB_IN_B1_valid, SB_T1_EAST_SB_IN_B1_valid, SB_T1_SOUTH_SB_IN_B1_valid, SB_T1_NORTH_SB_IN_B1_valid, SB_T0_WEST_SB_IN_B1_valid, SB_T0_EAST_SB_IN_B1_valid, SB_T0_SOUTH_SB_IN_B1_valid, SB_T0_NORTH_SB_IN_B1_valid};
	CB_MEM_input_width_1_num_1 CB_MEM_input_width_1_num_1(
		.I(CB_MEM_input_width_1_num_1_I),
		.O(CB_MEM_input_width_1_num_1_O),
		.clk(clk),
		.config_config_addr(self_config_config_addr_out[31:24]),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_8_out),
		.enable(CB_MEM_input_width_1_num_1_enable),
		.out_sel(CB_MEM_input_width_1_num_1_out_sel),
		.read_config_data(CB_MEM_input_width_1_num_1_read_config_data),
		.ready_in(MemCore_inst0_MEM_input_width_1_num_1_ready),
		.ready_out(CB_MEM_input_width_1_num_1_ready_out),
		.reset(reset),
		.valid_in(CB_MEM_input_width_1_num_1_valid_in),
		.valid_out(CB_MEM_input_width_1_num_1_valid_out)
	);
	wire [19:0] CB_flush_I;
	assign CB_flush_I[19+:1] = SB_T4_WEST_SB_IN_B1;
	assign CB_flush_I[18+:1] = SB_T4_EAST_SB_IN_B1;
	assign CB_flush_I[17+:1] = SB_T4_SOUTH_SB_IN_B1;
	assign CB_flush_I[16+:1] = SB_T4_NORTH_SB_IN_B1;
	assign CB_flush_I[15+:1] = SB_T3_WEST_SB_IN_B1;
	assign CB_flush_I[14+:1] = SB_T3_EAST_SB_IN_B1;
	assign CB_flush_I[13+:1] = SB_T3_SOUTH_SB_IN_B1;
	assign CB_flush_I[12+:1] = SB_T3_NORTH_SB_IN_B1;
	assign CB_flush_I[11+:1] = SB_T2_WEST_SB_IN_B1;
	assign CB_flush_I[10+:1] = SB_T2_EAST_SB_IN_B1;
	assign CB_flush_I[9+:1] = SB_T2_SOUTH_SB_IN_B1;
	assign CB_flush_I[8+:1] = SB_T2_NORTH_SB_IN_B1;
	assign CB_flush_I[7+:1] = SB_T1_WEST_SB_IN_B1;
	assign CB_flush_I[6+:1] = SB_T1_EAST_SB_IN_B1;
	assign CB_flush_I[5+:1] = SB_T1_SOUTH_SB_IN_B1;
	assign CB_flush_I[4+:1] = SB_T1_NORTH_SB_IN_B1;
	assign CB_flush_I[3+:1] = SB_T0_WEST_SB_IN_B1;
	assign CB_flush_I[2+:1] = SB_T0_EAST_SB_IN_B1;
	assign CB_flush_I[1+:1] = SB_T0_SOUTH_SB_IN_B1;
	assign CB_flush_I[0+:1] = SB_T0_NORTH_SB_IN_B1;
	wire [19:0] CB_flush_valid_in;
	assign CB_flush_valid_in = {SB_T4_WEST_SB_IN_B1_valid, SB_T4_EAST_SB_IN_B1_valid, SB_T4_SOUTH_SB_IN_B1_valid, SB_T4_NORTH_SB_IN_B1_valid, SB_T3_WEST_SB_IN_B1_valid, SB_T3_EAST_SB_IN_B1_valid, SB_T3_SOUTH_SB_IN_B1_valid, SB_T3_NORTH_SB_IN_B1_valid, SB_T2_WEST_SB_IN_B1_valid, SB_T2_EAST_SB_IN_B1_valid, SB_T2_SOUTH_SB_IN_B1_valid, SB_T2_NORTH_SB_IN_B1_valid, SB_T1_WEST_SB_IN_B1_valid, SB_T1_EAST_SB_IN_B1_valid, SB_T1_SOUTH_SB_IN_B1_valid, SB_T1_NORTH_SB_IN_B1_valid, SB_T0_WEST_SB_IN_B1_valid, SB_T0_EAST_SB_IN_B1_valid, SB_T0_SOUTH_SB_IN_B1_valid, SB_T0_NORTH_SB_IN_B1_valid};
	CB_flush CB_flush(
		.I(CB_flush_I),
		.O(CB_flush_O),
		.clk(clk),
		.config_config_addr(self_config_config_addr_out[31:24]),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_9_out),
		.enable(CB_flush_enable),
		.out_sel(CB_flush_out_sel),
		.read_config_data(CB_flush_read_config_data),
		.ready_in(bit_const_1_None_out),
		.ready_out(CB_flush_ready_out),
		.reset(reset),
		.valid_in(CB_flush_valid_in),
		.valid_out(CB_flush_valid_out)
	);
	Decode08 DECODE_FEATURE_0(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_0_O)
	);
	Decode18 DECODE_FEATURE_1(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_1_O)
	);
	Decode108 DECODE_FEATURE_10(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_10_O)
	);
	Decode118 DECODE_FEATURE_11(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_11_O)
	);
	Decode128 DECODE_FEATURE_12(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_12_O)
	);
	Decode28 DECODE_FEATURE_2(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_2_O)
	);
	Decode38 DECODE_FEATURE_3(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_3_O)
	);
	Decode48 DECODE_FEATURE_4(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_4_O)
	);
	Decode58 DECODE_FEATURE_5(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_5_O)
	);
	Decode68 DECODE_FEATURE_6(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_6_O)
	);
	Decode78 DECODE_FEATURE_7(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_7_O)
	);
	Decode88 DECODE_FEATURE_8(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_8_O)
	);
	Decode98 DECODE_FEATURE_9(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_9_O)
	);
	corebit_and FEATURE_AND_0(
		.in0(DECODE_FEATURE_0_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_0_out)
	);
	corebit_and FEATURE_AND_1(
		.in0(DECODE_FEATURE_1_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_1_out)
	);
	corebit_and FEATURE_AND_10(
		.in0(DECODE_FEATURE_10_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_10_out)
	);
	corebit_and FEATURE_AND_11(
		.in0(DECODE_FEATURE_11_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_11_out)
	);
	corebit_and FEATURE_AND_12(
		.in0(DECODE_FEATURE_12_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_12_out)
	);
	corebit_and FEATURE_AND_2(
		.in0(DECODE_FEATURE_2_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_2_out)
	);
	corebit_and FEATURE_AND_3(
		.in0(DECODE_FEATURE_3_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_3_out)
	);
	corebit_and FEATURE_AND_4(
		.in0(DECODE_FEATURE_4_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_4_out)
	);
	corebit_and FEATURE_AND_5(
		.in0(DECODE_FEATURE_5_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_5_out)
	);
	corebit_and FEATURE_AND_6(
		.in0(DECODE_FEATURE_6_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_6_out)
	);
	corebit_and FEATURE_AND_7(
		.in0(DECODE_FEATURE_7_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_7_out)
	);
	corebit_and FEATURE_AND_8(
		.in0(DECODE_FEATURE_8_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_8_out)
	);
	corebit_and FEATURE_AND_9(
		.in0(DECODE_FEATURE_9_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_9_out)
	);
	ReadyValidLoopBack MEM_output_width_17_num_0_loopback(
		.valid_out(MEM_output_width_17_num_0_loopback_valid_out),
		.ready_in(SB_ID0_5TRACKS_B17_MemCore_MEM_output_width_17_num_0_ready_out),
		.valid_in(MemCore_inst0_MEM_output_width_17_num_0_valid)
	);
	ReadyValidLoopBack MEM_output_width_17_num_1_loopback(
		.valid_out(MEM_output_width_17_num_1_loopback_valid_out),
		.ready_in(SB_ID0_5TRACKS_B17_MemCore_MEM_output_width_17_num_1_ready_out),
		.valid_in(MemCore_inst0_MEM_output_width_17_num_1_valid)
	);
	ReadyValidLoopBack MEM_output_width_17_num_2_loopback(
		.valid_out(MEM_output_width_17_num_2_loopback_valid_out),
		.ready_in(SB_ID0_5TRACKS_B17_MemCore_MEM_output_width_17_num_2_ready_out),
		.valid_in(MemCore_inst0_MEM_output_width_17_num_2_valid)
	);
	ReadyValidLoopBack MEM_output_width_1_num_0_loopback(
		.valid_out(MEM_output_width_1_num_0_loopback_valid_out),
		.ready_in(SB_ID0_5TRACKS_B1_MemCore_MEM_output_width_1_num_0_ready_out),
		.valid_in(MemCore_inst0_MEM_output_width_1_num_0_valid)
	);
	ReadyValidLoopBack MEM_output_width_1_num_1_loopback(
		.valid_out(MEM_output_width_1_num_1_loopback_valid_out),
		.ready_in(SB_ID0_5TRACKS_B1_MemCore_MEM_output_width_1_num_1_ready_out),
		.valid_in(MemCore_inst0_MEM_output_width_1_num_1_valid)
	);
	ReadyValidLoopBack MEM_output_width_1_num_2_loopback(
		.valid_out(MEM_output_width_1_num_2_loopback_valid_out),
		.ready_in(SB_ID0_5TRACKS_B1_MemCore_MEM_output_width_1_num_2_ready_out),
		.valid_in(MemCore_inst0_MEM_output_width_1_num_2_valid)
	);
	MemCore MemCore_inst0(
		.MEM_input_width_17_num_0(CB_MEM_input_width_17_num_0_O),
		.MEM_input_width_17_num_0_ready(MemCore_inst0_MEM_input_width_17_num_0_ready),
		.MEM_input_width_17_num_0_valid(CB_MEM_input_width_17_num_0_valid_out),
		.MEM_input_width_17_num_1(CB_MEM_input_width_17_num_1_O),
		.MEM_input_width_17_num_1_ready(MemCore_inst0_MEM_input_width_17_num_1_ready),
		.MEM_input_width_17_num_1_valid(CB_MEM_input_width_17_num_1_valid_out),
		.MEM_input_width_17_num_2(CB_MEM_input_width_17_num_2_O),
		.MEM_input_width_17_num_2_ready(MemCore_inst0_MEM_input_width_17_num_2_ready),
		.MEM_input_width_17_num_2_valid(CB_MEM_input_width_17_num_2_valid_out),
		.MEM_input_width_17_num_3(CB_MEM_input_width_17_num_3_O),
		.MEM_input_width_17_num_3_ready(MemCore_inst0_MEM_input_width_17_num_3_ready),
		.MEM_input_width_17_num_3_valid(CB_MEM_input_width_17_num_3_valid_out),
		.MEM_input_width_1_num_0(CB_MEM_input_width_1_num_0_O),
		.MEM_input_width_1_num_0_ready(MemCore_inst0_MEM_input_width_1_num_0_ready),
		.MEM_input_width_1_num_0_valid(CB_MEM_input_width_1_num_0_valid_out),
		.MEM_input_width_1_num_1(CB_MEM_input_width_1_num_1_O),
		.MEM_input_width_1_num_1_ready(MemCore_inst0_MEM_input_width_1_num_1_ready),
		.MEM_input_width_1_num_1_valid(CB_MEM_input_width_1_num_1_valid_out),
		.MEM_output_width_17_num_0(MemCore_inst0_MEM_output_width_17_num_0),
		.MEM_output_width_17_num_0_ready(SB_ID0_5TRACKS_B17_MemCore_MEM_output_width_17_num_0_ready_out),
		.MEM_output_width_17_num_0_valid(MemCore_inst0_MEM_output_width_17_num_0_valid),
		.MEM_output_width_17_num_1(MemCore_inst0_MEM_output_width_17_num_1),
		.MEM_output_width_17_num_1_ready(SB_ID0_5TRACKS_B17_MemCore_MEM_output_width_17_num_1_ready_out),
		.MEM_output_width_17_num_1_valid(MemCore_inst0_MEM_output_width_17_num_1_valid),
		.MEM_output_width_17_num_2(MemCore_inst0_MEM_output_width_17_num_2),
		.MEM_output_width_17_num_2_ready(SB_ID0_5TRACKS_B17_MemCore_MEM_output_width_17_num_2_ready_out),
		.MEM_output_width_17_num_2_valid(MemCore_inst0_MEM_output_width_17_num_2_valid),
		.MEM_output_width_1_num_0(MemCore_inst0_MEM_output_width_1_num_0),
		.MEM_output_width_1_num_0_ready(SB_ID0_5TRACKS_B1_MemCore_MEM_output_width_1_num_0_ready_out),
		.MEM_output_width_1_num_0_valid(MemCore_inst0_MEM_output_width_1_num_0_valid),
		.MEM_output_width_1_num_1(MemCore_inst0_MEM_output_width_1_num_1),
		.MEM_output_width_1_num_1_ready(SB_ID0_5TRACKS_B1_MemCore_MEM_output_width_1_num_1_ready_out),
		.MEM_output_width_1_num_1_valid(MemCore_inst0_MEM_output_width_1_num_1_valid),
		.MEM_output_width_1_num_2(MemCore_inst0_MEM_output_width_1_num_2),
		.MEM_output_width_1_num_2_ready(SB_ID0_5TRACKS_B1_MemCore_MEM_output_width_1_num_2_ready_out),
		.MEM_output_width_1_num_2_valid(MemCore_inst0_MEM_output_width_1_num_2_valid),
		.clk(clk),
		.config_1_config_addr(self_config_config_addr_out[31:24]),
		.config_1_config_data(config_config_data),
		.config_1_read(config_read),
		.config_1_write(FEATURE_AND_1_out),
		.config_2_config_addr(self_config_config_addr_out[31:24]),
		.config_2_config_data(config_config_data),
		.config_2_read(config_read),
		.config_2_write(FEATURE_AND_2_out),
		.config_config_addr(self_config_config_addr_out[31:24]),
		.config_config_data(config_config_data),
		.config_en_0(DECODE_FEATURE_1_O),
		.config_en_1(DECODE_FEATURE_2_O),
		.config_read(config_read),
		.config_write(FEATURE_AND_0_out),
		.flush(CB_flush_O),
		.flush_core(flush),
		.read_config_data(MemCore_inst0_read_config_data),
		.read_config_data_1(MemCore_inst0_read_config_data_1),
		.read_config_data_2(MemCore_inst0_read_config_data_2),
		.reset(reset),
		.stall(stall)
	);
	PowerDomainConfigReg PowerDomainConfigReg_inst0(
		.clk(clk),
		.config_config_addr(self_config_config_addr_out[31:24]),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_12_out),
		.ps_en_out(PowerDomainConfigReg_inst0_ps_en_out),
		.read_config_data(PowerDomainConfigReg_inst0_read_config_data),
		.reset(reset)
	);
	PowerDomainOR PowerDomainOR(
		.I0(read_data_mux_O),
		.I1(read_config_data_in),
		.O(PowerDomainOR_O),
		.I_not(PowerDomainConfigReg_inst0_ps_en_out)
	);
	SB_ID0_5TRACKS_B17_MemCore SB_ID0_5TRACKS_B17_MemCore(
		.MEM_input_width_17_num_0_enable(CB_MEM_input_width_17_num_0_enable),
		.MEM_input_width_17_num_0_out_sel(CB_MEM_input_width_17_num_0_out_sel),
		.MEM_input_width_17_num_0_ready(CB_MEM_input_width_17_num_0_ready_out),
		.MEM_input_width_17_num_1_enable(CB_MEM_input_width_17_num_1_enable),
		.MEM_input_width_17_num_1_out_sel(CB_MEM_input_width_17_num_1_out_sel),
		.MEM_input_width_17_num_1_ready(CB_MEM_input_width_17_num_1_ready_out),
		.MEM_input_width_17_num_2_enable(CB_MEM_input_width_17_num_2_enable),
		.MEM_input_width_17_num_2_out_sel(CB_MEM_input_width_17_num_2_out_sel),
		.MEM_input_width_17_num_2_ready(CB_MEM_input_width_17_num_2_ready_out),
		.MEM_input_width_17_num_3_enable(CB_MEM_input_width_17_num_3_enable),
		.MEM_input_width_17_num_3_out_sel(CB_MEM_input_width_17_num_3_out_sel),
		.MEM_input_width_17_num_3_ready(CB_MEM_input_width_17_num_3_ready_out),
		.MEM_output_width_17_num_0(MemCore_inst0_MEM_output_width_17_num_0),
		.MEM_output_width_17_num_0_ready_out(SB_ID0_5TRACKS_B17_MemCore_MEM_output_width_17_num_0_ready_out),
		.MEM_output_width_17_num_0_valid(MEM_output_width_17_num_0_loopback_valid_out[0]),
		.MEM_output_width_17_num_1(MemCore_inst0_MEM_output_width_17_num_1),
		.MEM_output_width_17_num_1_ready_out(SB_ID0_5TRACKS_B17_MemCore_MEM_output_width_17_num_1_ready_out),
		.MEM_output_width_17_num_1_valid(MEM_output_width_17_num_1_loopback_valid_out[0]),
		.MEM_output_width_17_num_2(MemCore_inst0_MEM_output_width_17_num_2),
		.MEM_output_width_17_num_2_ready_out(SB_ID0_5TRACKS_B17_MemCore_MEM_output_width_17_num_2_ready_out),
		.MEM_output_width_17_num_2_valid(MEM_output_width_17_num_2_loopback_valid_out[0]),
		.SB_T0_EAST_SB_IN_B17(SB_T0_EAST_SB_IN_B17),
		.SB_T0_EAST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T0_EAST_SB_IN_B17_enable),
		.SB_T0_EAST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T0_EAST_SB_IN_B17_ready_out),
		.SB_T0_EAST_SB_IN_B17_valid_in(SB_T0_EAST_SB_IN_B17_valid),
		.SB_T0_EAST_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_EAST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T0_EAST_SB_OUT_B17_enable),
		.SB_T0_EAST_SB_OUT_B17_ready_in(SB_T0_EAST_SB_OUT_B17_ready_and_Z),
		.SB_T0_EAST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T0_EAST_SB_OUT_B17_valid_out),
		.SB_T0_NORTH_SB_IN_B17(SB_T0_NORTH_SB_IN_B17),
		.SB_T0_NORTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T0_NORTH_SB_IN_B17_enable),
		.SB_T0_NORTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T0_NORTH_SB_IN_B17_ready_out),
		.SB_T0_NORTH_SB_IN_B17_valid_in(SB_T0_NORTH_SB_IN_B17_valid),
		.SB_T0_NORTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T0_NORTH_SB_OUT_B17_enable),
		.SB_T0_NORTH_SB_OUT_B17_ready_in(SB_T0_NORTH_SB_OUT_B17_ready_and_Z),
		.SB_T0_NORTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T0_NORTH_SB_OUT_B17_valid_out),
		.SB_T0_SOUTH_SB_IN_B17(SB_T0_SOUTH_SB_IN_B17),
		.SB_T0_SOUTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T0_SOUTH_SB_IN_B17_enable),
		.SB_T0_SOUTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T0_SOUTH_SB_IN_B17_ready_out),
		.SB_T0_SOUTH_SB_IN_B17_valid_in(SB_T0_SOUTH_SB_IN_B17_valid),
		.SB_T0_SOUTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T0_SOUTH_SB_OUT_B17_enable),
		.SB_T0_SOUTH_SB_OUT_B17_ready_in(SB_T0_SOUTH_SB_OUT_B17_ready_and_Z),
		.SB_T0_SOUTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T0_SOUTH_SB_OUT_B17_valid_out),
		.SB_T0_WEST_SB_IN_B17(SB_T0_WEST_SB_IN_B17),
		.SB_T0_WEST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T0_WEST_SB_IN_B17_enable),
		.SB_T0_WEST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T0_WEST_SB_IN_B17_ready_out),
		.SB_T0_WEST_SB_IN_B17_valid_in(SB_T0_WEST_SB_IN_B17_valid),
		.SB_T0_WEST_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_WEST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T0_WEST_SB_OUT_B17_enable),
		.SB_T0_WEST_SB_OUT_B17_ready_in(SB_T0_WEST_SB_OUT_B17_ready_and_Z),
		.SB_T0_WEST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T0_WEST_SB_OUT_B17_valid_out),
		.SB_T1_EAST_SB_IN_B17(SB_T1_EAST_SB_IN_B17),
		.SB_T1_EAST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T1_EAST_SB_IN_B17_enable),
		.SB_T1_EAST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T1_EAST_SB_IN_B17_ready_out),
		.SB_T1_EAST_SB_IN_B17_valid_in(SB_T1_EAST_SB_IN_B17_valid),
		.SB_T1_EAST_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_EAST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T1_EAST_SB_OUT_B17_enable),
		.SB_T1_EAST_SB_OUT_B17_ready_in(SB_T1_EAST_SB_OUT_B17_ready_and_Z),
		.SB_T1_EAST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T1_EAST_SB_OUT_B17_valid_out),
		.SB_T1_NORTH_SB_IN_B17(SB_T1_NORTH_SB_IN_B17),
		.SB_T1_NORTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T1_NORTH_SB_IN_B17_enable),
		.SB_T1_NORTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T1_NORTH_SB_IN_B17_ready_out),
		.SB_T1_NORTH_SB_IN_B17_valid_in(SB_T1_NORTH_SB_IN_B17_valid),
		.SB_T1_NORTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T1_NORTH_SB_OUT_B17_enable),
		.SB_T1_NORTH_SB_OUT_B17_ready_in(SB_T1_NORTH_SB_OUT_B17_ready_and_Z),
		.SB_T1_NORTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T1_NORTH_SB_OUT_B17_valid_out),
		.SB_T1_SOUTH_SB_IN_B17(SB_T1_SOUTH_SB_IN_B17),
		.SB_T1_SOUTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T1_SOUTH_SB_IN_B17_enable),
		.SB_T1_SOUTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T1_SOUTH_SB_IN_B17_ready_out),
		.SB_T1_SOUTH_SB_IN_B17_valid_in(SB_T1_SOUTH_SB_IN_B17_valid),
		.SB_T1_SOUTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T1_SOUTH_SB_OUT_B17_enable),
		.SB_T1_SOUTH_SB_OUT_B17_ready_in(SB_T1_SOUTH_SB_OUT_B17_ready_and_Z),
		.SB_T1_SOUTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T1_SOUTH_SB_OUT_B17_valid_out),
		.SB_T1_WEST_SB_IN_B17(SB_T1_WEST_SB_IN_B17),
		.SB_T1_WEST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T1_WEST_SB_IN_B17_enable),
		.SB_T1_WEST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T1_WEST_SB_IN_B17_ready_out),
		.SB_T1_WEST_SB_IN_B17_valid_in(SB_T1_WEST_SB_IN_B17_valid),
		.SB_T1_WEST_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_WEST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T1_WEST_SB_OUT_B17_enable),
		.SB_T1_WEST_SB_OUT_B17_ready_in(SB_T1_WEST_SB_OUT_B17_ready_and_Z),
		.SB_T1_WEST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T1_WEST_SB_OUT_B17_valid_out),
		.SB_T2_EAST_SB_IN_B17(SB_T2_EAST_SB_IN_B17),
		.SB_T2_EAST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T2_EAST_SB_IN_B17_enable),
		.SB_T2_EAST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T2_EAST_SB_IN_B17_ready_out),
		.SB_T2_EAST_SB_IN_B17_valid_in(SB_T2_EAST_SB_IN_B17_valid),
		.SB_T2_EAST_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_EAST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T2_EAST_SB_OUT_B17_enable),
		.SB_T2_EAST_SB_OUT_B17_ready_in(SB_T2_EAST_SB_OUT_B17_ready_and_Z),
		.SB_T2_EAST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T2_EAST_SB_OUT_B17_valid_out),
		.SB_T2_NORTH_SB_IN_B17(SB_T2_NORTH_SB_IN_B17),
		.SB_T2_NORTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T2_NORTH_SB_IN_B17_enable),
		.SB_T2_NORTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T2_NORTH_SB_IN_B17_ready_out),
		.SB_T2_NORTH_SB_IN_B17_valid_in(SB_T2_NORTH_SB_IN_B17_valid),
		.SB_T2_NORTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T2_NORTH_SB_OUT_B17_enable),
		.SB_T2_NORTH_SB_OUT_B17_ready_in(SB_T2_NORTH_SB_OUT_B17_ready_and_Z),
		.SB_T2_NORTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T2_NORTH_SB_OUT_B17_valid_out),
		.SB_T2_SOUTH_SB_IN_B17(SB_T2_SOUTH_SB_IN_B17),
		.SB_T2_SOUTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T2_SOUTH_SB_IN_B17_enable),
		.SB_T2_SOUTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T2_SOUTH_SB_IN_B17_ready_out),
		.SB_T2_SOUTH_SB_IN_B17_valid_in(SB_T2_SOUTH_SB_IN_B17_valid),
		.SB_T2_SOUTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T2_SOUTH_SB_OUT_B17_enable),
		.SB_T2_SOUTH_SB_OUT_B17_ready_in(SB_T2_SOUTH_SB_OUT_B17_ready_and_Z),
		.SB_T2_SOUTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T2_SOUTH_SB_OUT_B17_valid_out),
		.SB_T2_WEST_SB_IN_B17(SB_T2_WEST_SB_IN_B17),
		.SB_T2_WEST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T2_WEST_SB_IN_B17_enable),
		.SB_T2_WEST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T2_WEST_SB_IN_B17_ready_out),
		.SB_T2_WEST_SB_IN_B17_valid_in(SB_T2_WEST_SB_IN_B17_valid),
		.SB_T2_WEST_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_WEST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T2_WEST_SB_OUT_B17_enable),
		.SB_T2_WEST_SB_OUT_B17_ready_in(SB_T2_WEST_SB_OUT_B17_ready_and_Z),
		.SB_T2_WEST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T2_WEST_SB_OUT_B17_valid_out),
		.SB_T3_EAST_SB_IN_B17(SB_T3_EAST_SB_IN_B17),
		.SB_T3_EAST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T3_EAST_SB_IN_B17_enable),
		.SB_T3_EAST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T3_EAST_SB_IN_B17_ready_out),
		.SB_T3_EAST_SB_IN_B17_valid_in(SB_T3_EAST_SB_IN_B17_valid),
		.SB_T3_EAST_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_EAST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T3_EAST_SB_OUT_B17_enable),
		.SB_T3_EAST_SB_OUT_B17_ready_in(SB_T3_EAST_SB_OUT_B17_ready_and_Z),
		.SB_T3_EAST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T3_EAST_SB_OUT_B17_valid_out),
		.SB_T3_NORTH_SB_IN_B17(SB_T3_NORTH_SB_IN_B17),
		.SB_T3_NORTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T3_NORTH_SB_IN_B17_enable),
		.SB_T3_NORTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T3_NORTH_SB_IN_B17_ready_out),
		.SB_T3_NORTH_SB_IN_B17_valid_in(SB_T3_NORTH_SB_IN_B17_valid),
		.SB_T3_NORTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T3_NORTH_SB_OUT_B17_enable),
		.SB_T3_NORTH_SB_OUT_B17_ready_in(SB_T3_NORTH_SB_OUT_B17_ready_and_Z),
		.SB_T3_NORTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T3_NORTH_SB_OUT_B17_valid_out),
		.SB_T3_SOUTH_SB_IN_B17(SB_T3_SOUTH_SB_IN_B17),
		.SB_T3_SOUTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T3_SOUTH_SB_IN_B17_enable),
		.SB_T3_SOUTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T3_SOUTH_SB_IN_B17_ready_out),
		.SB_T3_SOUTH_SB_IN_B17_valid_in(SB_T3_SOUTH_SB_IN_B17_valid),
		.SB_T3_SOUTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T3_SOUTH_SB_OUT_B17_enable),
		.SB_T3_SOUTH_SB_OUT_B17_ready_in(SB_T3_SOUTH_SB_OUT_B17_ready_and_Z),
		.SB_T3_SOUTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T3_SOUTH_SB_OUT_B17_valid_out),
		.SB_T3_WEST_SB_IN_B17(SB_T3_WEST_SB_IN_B17),
		.SB_T3_WEST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T3_WEST_SB_IN_B17_enable),
		.SB_T3_WEST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T3_WEST_SB_IN_B17_ready_out),
		.SB_T3_WEST_SB_IN_B17_valid_in(SB_T3_WEST_SB_IN_B17_valid),
		.SB_T3_WEST_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_WEST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T3_WEST_SB_OUT_B17_enable),
		.SB_T3_WEST_SB_OUT_B17_ready_in(SB_T3_WEST_SB_OUT_B17_ready_and_Z),
		.SB_T3_WEST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T3_WEST_SB_OUT_B17_valid_out),
		.SB_T4_EAST_SB_IN_B17(SB_T4_EAST_SB_IN_B17),
		.SB_T4_EAST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T4_EAST_SB_IN_B17_enable),
		.SB_T4_EAST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T4_EAST_SB_IN_B17_ready_out),
		.SB_T4_EAST_SB_IN_B17_valid_in(SB_T4_EAST_SB_IN_B17_valid),
		.SB_T4_EAST_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_EAST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T4_EAST_SB_OUT_B17_enable),
		.SB_T4_EAST_SB_OUT_B17_ready_in(SB_T4_EAST_SB_OUT_B17_ready_and_Z),
		.SB_T4_EAST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T4_EAST_SB_OUT_B17_valid_out),
		.SB_T4_NORTH_SB_IN_B17(SB_T4_NORTH_SB_IN_B17),
		.SB_T4_NORTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T4_NORTH_SB_IN_B17_enable),
		.SB_T4_NORTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T4_NORTH_SB_IN_B17_ready_out),
		.SB_T4_NORTH_SB_IN_B17_valid_in(SB_T4_NORTH_SB_IN_B17_valid),
		.SB_T4_NORTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T4_NORTH_SB_OUT_B17_enable),
		.SB_T4_NORTH_SB_OUT_B17_ready_in(SB_T4_NORTH_SB_OUT_B17_ready_and_Z),
		.SB_T4_NORTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T4_NORTH_SB_OUT_B17_valid_out),
		.SB_T4_SOUTH_SB_IN_B17(SB_T4_SOUTH_SB_IN_B17),
		.SB_T4_SOUTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T4_SOUTH_SB_IN_B17_enable),
		.SB_T4_SOUTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T4_SOUTH_SB_IN_B17_ready_out),
		.SB_T4_SOUTH_SB_IN_B17_valid_in(SB_T4_SOUTH_SB_IN_B17_valid),
		.SB_T4_SOUTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T4_SOUTH_SB_OUT_B17_enable),
		.SB_T4_SOUTH_SB_OUT_B17_ready_in(SB_T4_SOUTH_SB_OUT_B17_ready_and_Z),
		.SB_T4_SOUTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T4_SOUTH_SB_OUT_B17_valid_out),
		.SB_T4_WEST_SB_IN_B17(SB_T4_WEST_SB_IN_B17),
		.SB_T4_WEST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T4_WEST_SB_IN_B17_enable),
		.SB_T4_WEST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T4_WEST_SB_IN_B17_ready_out),
		.SB_T4_WEST_SB_IN_B17_valid_in(SB_T4_WEST_SB_IN_B17_valid),
		.SB_T4_WEST_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_WEST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T4_WEST_SB_OUT_B17_enable),
		.SB_T4_WEST_SB_OUT_B17_ready_in(SB_T4_WEST_SB_OUT_B17_ready_and_Z),
		.SB_T4_WEST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T4_WEST_SB_OUT_B17_valid_out),
		.clk(clk),
		.config_config_addr(self_config_config_addr_out[31:24]),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_11_out),
		.read_config_data(SB_ID0_5TRACKS_B17_MemCore_read_config_data),
		.reset(reset),
		.stall(stall)
	);
	SB_ID0_5TRACKS_B1_MemCore SB_ID0_5TRACKS_B1_MemCore(
		.MEM_input_width_1_num_0_enable(CB_MEM_input_width_1_num_0_enable),
		.MEM_input_width_1_num_0_out_sel(CB_MEM_input_width_1_num_0_out_sel),
		.MEM_input_width_1_num_0_ready(CB_MEM_input_width_1_num_0_ready_out),
		.MEM_input_width_1_num_1_enable(CB_MEM_input_width_1_num_1_enable),
		.MEM_input_width_1_num_1_out_sel(CB_MEM_input_width_1_num_1_out_sel),
		.MEM_input_width_1_num_1_ready(CB_MEM_input_width_1_num_1_ready_out),
		.MEM_output_width_1_num_0(MemCore_inst0_MEM_output_width_1_num_0),
		.MEM_output_width_1_num_0_ready_out(SB_ID0_5TRACKS_B1_MemCore_MEM_output_width_1_num_0_ready_out),
		.MEM_output_width_1_num_0_valid(MEM_output_width_1_num_0_loopback_valid_out[0]),
		.MEM_output_width_1_num_1(MemCore_inst0_MEM_output_width_1_num_1),
		.MEM_output_width_1_num_1_ready_out(SB_ID0_5TRACKS_B1_MemCore_MEM_output_width_1_num_1_ready_out),
		.MEM_output_width_1_num_1_valid(MEM_output_width_1_num_1_loopback_valid_out[0]),
		.MEM_output_width_1_num_2(MemCore_inst0_MEM_output_width_1_num_2),
		.MEM_output_width_1_num_2_ready_out(SB_ID0_5TRACKS_B1_MemCore_MEM_output_width_1_num_2_ready_out),
		.MEM_output_width_1_num_2_valid(MEM_output_width_1_num_2_loopback_valid_out[0]),
		.SB_T0_EAST_SB_IN_B1(SB_T0_EAST_SB_IN_B1),
		.SB_T0_EAST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_IN_B1_enable),
		.SB_T0_EAST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_IN_B1_ready_out),
		.SB_T0_EAST_SB_IN_B1_valid_in(SB_T0_EAST_SB_IN_B1_valid),
		.SB_T0_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_EAST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_OUT_B1_enable),
		.SB_T0_EAST_SB_OUT_B1_ready_in(SB_T0_EAST_SB_OUT_B1_ready_and_Z),
		.SB_T0_EAST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_OUT_B1_valid_out),
		.SB_T0_NORTH_SB_IN_B1(SB_T0_NORTH_SB_IN_B1),
		.SB_T0_NORTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_IN_B1_enable),
		.SB_T0_NORTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_IN_B1_ready_out),
		.SB_T0_NORTH_SB_IN_B1_valid_in(SB_T0_NORTH_SB_IN_B1_valid),
		.SB_T0_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_OUT_B1_enable),
		.SB_T0_NORTH_SB_OUT_B1_ready_in(SB_T0_NORTH_SB_OUT_B1_ready_and_Z),
		.SB_T0_NORTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_OUT_B1_valid_out),
		.SB_T0_SOUTH_SB_IN_B1(SB_T0_SOUTH_SB_IN_B1),
		.SB_T0_SOUTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_IN_B1_enable),
		.SB_T0_SOUTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_IN_B1_ready_out),
		.SB_T0_SOUTH_SB_IN_B1_valid_in(SB_T0_SOUTH_SB_IN_B1_valid),
		.SB_T0_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_OUT_B1_enable),
		.SB_T0_SOUTH_SB_OUT_B1_ready_in(SB_T0_SOUTH_SB_OUT_B1_ready_and_Z),
		.SB_T0_SOUTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_OUT_B1_valid_out),
		.SB_T0_WEST_SB_IN_B1(SB_T0_WEST_SB_IN_B1),
		.SB_T0_WEST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_IN_B1_enable),
		.SB_T0_WEST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_IN_B1_ready_out),
		.SB_T0_WEST_SB_IN_B1_valid_in(SB_T0_WEST_SB_IN_B1_valid),
		.SB_T0_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_WEST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_OUT_B1_enable),
		.SB_T0_WEST_SB_OUT_B1_ready_in(SB_T0_WEST_SB_OUT_B1_ready_and_Z),
		.SB_T0_WEST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_OUT_B1_valid_out),
		.SB_T1_EAST_SB_IN_B1(SB_T1_EAST_SB_IN_B1),
		.SB_T1_EAST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_IN_B1_enable),
		.SB_T1_EAST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_IN_B1_ready_out),
		.SB_T1_EAST_SB_IN_B1_valid_in(SB_T1_EAST_SB_IN_B1_valid),
		.SB_T1_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_EAST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_OUT_B1_enable),
		.SB_T1_EAST_SB_OUT_B1_ready_in(SB_T1_EAST_SB_OUT_B1_ready_and_Z),
		.SB_T1_EAST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_OUT_B1_valid_out),
		.SB_T1_NORTH_SB_IN_B1(SB_T1_NORTH_SB_IN_B1),
		.SB_T1_NORTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_IN_B1_enable),
		.SB_T1_NORTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_IN_B1_ready_out),
		.SB_T1_NORTH_SB_IN_B1_valid_in(SB_T1_NORTH_SB_IN_B1_valid),
		.SB_T1_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_OUT_B1_enable),
		.SB_T1_NORTH_SB_OUT_B1_ready_in(SB_T1_NORTH_SB_OUT_B1_ready_and_Z),
		.SB_T1_NORTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_OUT_B1_valid_out),
		.SB_T1_SOUTH_SB_IN_B1(SB_T1_SOUTH_SB_IN_B1),
		.SB_T1_SOUTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_IN_B1_enable),
		.SB_T1_SOUTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_IN_B1_ready_out),
		.SB_T1_SOUTH_SB_IN_B1_valid_in(SB_T1_SOUTH_SB_IN_B1_valid),
		.SB_T1_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_OUT_B1_enable),
		.SB_T1_SOUTH_SB_OUT_B1_ready_in(SB_T1_SOUTH_SB_OUT_B1_ready_and_Z),
		.SB_T1_SOUTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_OUT_B1_valid_out),
		.SB_T1_WEST_SB_IN_B1(SB_T1_WEST_SB_IN_B1),
		.SB_T1_WEST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_IN_B1_enable),
		.SB_T1_WEST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_IN_B1_ready_out),
		.SB_T1_WEST_SB_IN_B1_valid_in(SB_T1_WEST_SB_IN_B1_valid),
		.SB_T1_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_WEST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_OUT_B1_enable),
		.SB_T1_WEST_SB_OUT_B1_ready_in(SB_T1_WEST_SB_OUT_B1_ready_and_Z),
		.SB_T1_WEST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_OUT_B1_valid_out),
		.SB_T2_EAST_SB_IN_B1(SB_T2_EAST_SB_IN_B1),
		.SB_T2_EAST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_IN_B1_enable),
		.SB_T2_EAST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_IN_B1_ready_out),
		.SB_T2_EAST_SB_IN_B1_valid_in(SB_T2_EAST_SB_IN_B1_valid),
		.SB_T2_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_EAST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_OUT_B1_enable),
		.SB_T2_EAST_SB_OUT_B1_ready_in(SB_T2_EAST_SB_OUT_B1_ready_and_Z),
		.SB_T2_EAST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_OUT_B1_valid_out),
		.SB_T2_NORTH_SB_IN_B1(SB_T2_NORTH_SB_IN_B1),
		.SB_T2_NORTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_IN_B1_enable),
		.SB_T2_NORTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_IN_B1_ready_out),
		.SB_T2_NORTH_SB_IN_B1_valid_in(SB_T2_NORTH_SB_IN_B1_valid),
		.SB_T2_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_OUT_B1_enable),
		.SB_T2_NORTH_SB_OUT_B1_ready_in(SB_T2_NORTH_SB_OUT_B1_ready_and_Z),
		.SB_T2_NORTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_OUT_B1_valid_out),
		.SB_T2_SOUTH_SB_IN_B1(SB_T2_SOUTH_SB_IN_B1),
		.SB_T2_SOUTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_IN_B1_enable),
		.SB_T2_SOUTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_IN_B1_ready_out),
		.SB_T2_SOUTH_SB_IN_B1_valid_in(SB_T2_SOUTH_SB_IN_B1_valid),
		.SB_T2_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_OUT_B1_enable),
		.SB_T2_SOUTH_SB_OUT_B1_ready_in(SB_T2_SOUTH_SB_OUT_B1_ready_and_Z),
		.SB_T2_SOUTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_OUT_B1_valid_out),
		.SB_T2_WEST_SB_IN_B1(SB_T2_WEST_SB_IN_B1),
		.SB_T2_WEST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_IN_B1_enable),
		.SB_T2_WEST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_IN_B1_ready_out),
		.SB_T2_WEST_SB_IN_B1_valid_in(SB_T2_WEST_SB_IN_B1_valid),
		.SB_T2_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_WEST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_OUT_B1_enable),
		.SB_T2_WEST_SB_OUT_B1_ready_in(SB_T2_WEST_SB_OUT_B1_ready_and_Z),
		.SB_T2_WEST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_OUT_B1_valid_out),
		.SB_T3_EAST_SB_IN_B1(SB_T3_EAST_SB_IN_B1),
		.SB_T3_EAST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_IN_B1_enable),
		.SB_T3_EAST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_IN_B1_ready_out),
		.SB_T3_EAST_SB_IN_B1_valid_in(SB_T3_EAST_SB_IN_B1_valid),
		.SB_T3_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_EAST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_OUT_B1_enable),
		.SB_T3_EAST_SB_OUT_B1_ready_in(SB_T3_EAST_SB_OUT_B1_ready_and_Z),
		.SB_T3_EAST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_OUT_B1_valid_out),
		.SB_T3_NORTH_SB_IN_B1(SB_T3_NORTH_SB_IN_B1),
		.SB_T3_NORTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_IN_B1_enable),
		.SB_T3_NORTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_IN_B1_ready_out),
		.SB_T3_NORTH_SB_IN_B1_valid_in(SB_T3_NORTH_SB_IN_B1_valid),
		.SB_T3_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_OUT_B1_enable),
		.SB_T3_NORTH_SB_OUT_B1_ready_in(SB_T3_NORTH_SB_OUT_B1_ready_and_Z),
		.SB_T3_NORTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_OUT_B1_valid_out),
		.SB_T3_SOUTH_SB_IN_B1(SB_T3_SOUTH_SB_IN_B1),
		.SB_T3_SOUTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_IN_B1_enable),
		.SB_T3_SOUTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_IN_B1_ready_out),
		.SB_T3_SOUTH_SB_IN_B1_valid_in(SB_T3_SOUTH_SB_IN_B1_valid),
		.SB_T3_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_OUT_B1_enable),
		.SB_T3_SOUTH_SB_OUT_B1_ready_in(SB_T3_SOUTH_SB_OUT_B1_ready_and_Z),
		.SB_T3_SOUTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_OUT_B1_valid_out),
		.SB_T3_WEST_SB_IN_B1(SB_T3_WEST_SB_IN_B1),
		.SB_T3_WEST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_IN_B1_enable),
		.SB_T3_WEST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_IN_B1_ready_out),
		.SB_T3_WEST_SB_IN_B1_valid_in(SB_T3_WEST_SB_IN_B1_valid),
		.SB_T3_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_WEST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_OUT_B1_enable),
		.SB_T3_WEST_SB_OUT_B1_ready_in(SB_T3_WEST_SB_OUT_B1_ready_and_Z),
		.SB_T3_WEST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_OUT_B1_valid_out),
		.SB_T4_EAST_SB_IN_B1(SB_T4_EAST_SB_IN_B1),
		.SB_T4_EAST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_IN_B1_enable),
		.SB_T4_EAST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_IN_B1_ready_out),
		.SB_T4_EAST_SB_IN_B1_valid_in(SB_T4_EAST_SB_IN_B1_valid),
		.SB_T4_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_EAST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_OUT_B1_enable),
		.SB_T4_EAST_SB_OUT_B1_ready_in(SB_T4_EAST_SB_OUT_B1_ready_and_Z),
		.SB_T4_EAST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_OUT_B1_valid_out),
		.SB_T4_NORTH_SB_IN_B1(SB_T4_NORTH_SB_IN_B1),
		.SB_T4_NORTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_IN_B1_enable),
		.SB_T4_NORTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_IN_B1_ready_out),
		.SB_T4_NORTH_SB_IN_B1_valid_in(SB_T4_NORTH_SB_IN_B1_valid),
		.SB_T4_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_OUT_B1_enable),
		.SB_T4_NORTH_SB_OUT_B1_ready_in(SB_T4_NORTH_SB_OUT_B1_ready_and_Z),
		.SB_T4_NORTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_OUT_B1_valid_out),
		.SB_T4_SOUTH_SB_IN_B1(SB_T4_SOUTH_SB_IN_B1),
		.SB_T4_SOUTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_IN_B1_enable),
		.SB_T4_SOUTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_IN_B1_ready_out),
		.SB_T4_SOUTH_SB_IN_B1_valid_in(SB_T4_SOUTH_SB_IN_B1_valid),
		.SB_T4_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_OUT_B1_enable),
		.SB_T4_SOUTH_SB_OUT_B1_ready_in(SB_T4_SOUTH_SB_OUT_B1_ready_and_Z),
		.SB_T4_SOUTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_OUT_B1_valid_out),
		.SB_T4_WEST_SB_IN_B1(SB_T4_WEST_SB_IN_B1),
		.SB_T4_WEST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_IN_B1_enable),
		.SB_T4_WEST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_IN_B1_ready_out),
		.SB_T4_WEST_SB_IN_B1_valid_in(SB_T4_WEST_SB_IN_B1_valid),
		.SB_T4_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_WEST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_OUT_B1_enable),
		.SB_T4_WEST_SB_OUT_B1_ready_in(SB_T4_WEST_SB_OUT_B1_ready_and_Z),
		.SB_T4_WEST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_OUT_B1_valid_out),
		.clk(clk),
		.config_config_addr(self_config_config_addr_out[31:24]),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_10_out),
		.read_config_data(SB_ID0_5TRACKS_B1_MemCore_read_config_data),
		.reset(reset),
		.stall(stall)
	);
	and_cell SB_T0_EAST_SB_OUT_B17_ready_and(
		.A(SB_T0_EAST_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_MemCore_SB_T0_EAST_SB_OUT_B17_enable),
		.Z(SB_T0_EAST_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T0_EAST_SB_OUT_B1_ready_and(
		.A(SB_T0_EAST_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_OUT_B1_enable),
		.Z(SB_T0_EAST_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T0_NORTH_SB_OUT_B17_ready_and(
		.A(SB_T0_NORTH_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_MemCore_SB_T0_NORTH_SB_OUT_B17_enable),
		.Z(SB_T0_NORTH_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T0_NORTH_SB_OUT_B1_ready_and(
		.A(SB_T0_NORTH_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_OUT_B1_enable),
		.Z(SB_T0_NORTH_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T0_SOUTH_SB_OUT_B17_ready_and(
		.A(SB_T0_SOUTH_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_MemCore_SB_T0_SOUTH_SB_OUT_B17_enable),
		.Z(SB_T0_SOUTH_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T0_SOUTH_SB_OUT_B1_ready_and(
		.A(SB_T0_SOUTH_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_OUT_B1_enable),
		.Z(SB_T0_SOUTH_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T0_WEST_SB_OUT_B17_ready_and(
		.A(SB_T0_WEST_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_MemCore_SB_T0_WEST_SB_OUT_B17_enable),
		.Z(SB_T0_WEST_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T0_WEST_SB_OUT_B1_ready_and(
		.A(SB_T0_WEST_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_OUT_B1_enable),
		.Z(SB_T0_WEST_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T1_EAST_SB_OUT_B17_ready_and(
		.A(SB_T1_EAST_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_MemCore_SB_T1_EAST_SB_OUT_B17_enable),
		.Z(SB_T1_EAST_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T1_EAST_SB_OUT_B1_ready_and(
		.A(SB_T1_EAST_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_OUT_B1_enable),
		.Z(SB_T1_EAST_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T1_NORTH_SB_OUT_B17_ready_and(
		.A(SB_T1_NORTH_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_MemCore_SB_T1_NORTH_SB_OUT_B17_enable),
		.Z(SB_T1_NORTH_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T1_NORTH_SB_OUT_B1_ready_and(
		.A(SB_T1_NORTH_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_OUT_B1_enable),
		.Z(SB_T1_NORTH_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T1_SOUTH_SB_OUT_B17_ready_and(
		.A(SB_T1_SOUTH_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_MemCore_SB_T1_SOUTH_SB_OUT_B17_enable),
		.Z(SB_T1_SOUTH_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T1_SOUTH_SB_OUT_B1_ready_and(
		.A(SB_T1_SOUTH_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_OUT_B1_enable),
		.Z(SB_T1_SOUTH_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T1_WEST_SB_OUT_B17_ready_and(
		.A(SB_T1_WEST_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_MemCore_SB_T1_WEST_SB_OUT_B17_enable),
		.Z(SB_T1_WEST_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T1_WEST_SB_OUT_B1_ready_and(
		.A(SB_T1_WEST_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_OUT_B1_enable),
		.Z(SB_T1_WEST_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T2_EAST_SB_OUT_B17_ready_and(
		.A(SB_T2_EAST_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_MemCore_SB_T2_EAST_SB_OUT_B17_enable),
		.Z(SB_T2_EAST_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T2_EAST_SB_OUT_B1_ready_and(
		.A(SB_T2_EAST_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_OUT_B1_enable),
		.Z(SB_T2_EAST_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T2_NORTH_SB_OUT_B17_ready_and(
		.A(SB_T2_NORTH_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_MemCore_SB_T2_NORTH_SB_OUT_B17_enable),
		.Z(SB_T2_NORTH_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T2_NORTH_SB_OUT_B1_ready_and(
		.A(SB_T2_NORTH_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_OUT_B1_enable),
		.Z(SB_T2_NORTH_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T2_SOUTH_SB_OUT_B17_ready_and(
		.A(SB_T2_SOUTH_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_MemCore_SB_T2_SOUTH_SB_OUT_B17_enable),
		.Z(SB_T2_SOUTH_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T2_SOUTH_SB_OUT_B1_ready_and(
		.A(SB_T2_SOUTH_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_OUT_B1_enable),
		.Z(SB_T2_SOUTH_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T2_WEST_SB_OUT_B17_ready_and(
		.A(SB_T2_WEST_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_MemCore_SB_T2_WEST_SB_OUT_B17_enable),
		.Z(SB_T2_WEST_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T2_WEST_SB_OUT_B1_ready_and(
		.A(SB_T2_WEST_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_OUT_B1_enable),
		.Z(SB_T2_WEST_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T3_EAST_SB_OUT_B17_ready_and(
		.A(SB_T3_EAST_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_MemCore_SB_T3_EAST_SB_OUT_B17_enable),
		.Z(SB_T3_EAST_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T3_EAST_SB_OUT_B1_ready_and(
		.A(SB_T3_EAST_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_OUT_B1_enable),
		.Z(SB_T3_EAST_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T3_NORTH_SB_OUT_B17_ready_and(
		.A(SB_T3_NORTH_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_MemCore_SB_T3_NORTH_SB_OUT_B17_enable),
		.Z(SB_T3_NORTH_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T3_NORTH_SB_OUT_B1_ready_and(
		.A(SB_T3_NORTH_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_OUT_B1_enable),
		.Z(SB_T3_NORTH_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T3_SOUTH_SB_OUT_B17_ready_and(
		.A(SB_T3_SOUTH_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_MemCore_SB_T3_SOUTH_SB_OUT_B17_enable),
		.Z(SB_T3_SOUTH_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T3_SOUTH_SB_OUT_B1_ready_and(
		.A(SB_T3_SOUTH_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_OUT_B1_enable),
		.Z(SB_T3_SOUTH_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T3_WEST_SB_OUT_B17_ready_and(
		.A(SB_T3_WEST_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_MemCore_SB_T3_WEST_SB_OUT_B17_enable),
		.Z(SB_T3_WEST_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T3_WEST_SB_OUT_B1_ready_and(
		.A(SB_T3_WEST_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_OUT_B1_enable),
		.Z(SB_T3_WEST_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T4_EAST_SB_OUT_B17_ready_and(
		.A(SB_T4_EAST_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_MemCore_SB_T4_EAST_SB_OUT_B17_enable),
		.Z(SB_T4_EAST_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T4_EAST_SB_OUT_B1_ready_and(
		.A(SB_T4_EAST_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_OUT_B1_enable),
		.Z(SB_T4_EAST_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T4_NORTH_SB_OUT_B17_ready_and(
		.A(SB_T4_NORTH_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_MemCore_SB_T4_NORTH_SB_OUT_B17_enable),
		.Z(SB_T4_NORTH_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T4_NORTH_SB_OUT_B1_ready_and(
		.A(SB_T4_NORTH_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_OUT_B1_enable),
		.Z(SB_T4_NORTH_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T4_SOUTH_SB_OUT_B17_ready_and(
		.A(SB_T4_SOUTH_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_MemCore_SB_T4_SOUTH_SB_OUT_B17_enable),
		.Z(SB_T4_SOUTH_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T4_SOUTH_SB_OUT_B1_ready_and(
		.A(SB_T4_SOUTH_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_OUT_B1_enable),
		.Z(SB_T4_SOUTH_SB_OUT_B1_ready_and_Z)
	);
	and_cell SB_T4_WEST_SB_OUT_B17_ready_and(
		.A(SB_T4_WEST_SB_OUT_B17_ready),
		.B(SB_ID0_5TRACKS_B17_MemCore_SB_T4_WEST_SB_OUT_B17_enable),
		.Z(SB_T4_WEST_SB_OUT_B17_ready_and_Z)
	);
	and_cell SB_T4_WEST_SB_OUT_B1_ready_and(
		.A(SB_T4_WEST_SB_OUT_B1_ready),
		.B(SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_OUT_B1_enable),
		.Z(SB_T4_WEST_SB_OUT_B1_ready_and_Z)
	);
	corebit_and and_inst0(
		.in0(coreir_eq_16_inst0_out),
		.in1(config_read[0]),
		.out(and_inst0_out)
	);
	corebit_and and_inst1(
		.in0(coreir_eq_16_inst0_out),
		.in1(config_write[0]),
		.out(and_inst1_out)
	);
	corebit_const #(.value(1'b1)) bit_const_1_None(.out(bit_const_1_None_out));
	coreir_const #(
		.value(8'h00),
		.width(8)
	) const_0_8(.out(const_0_8_out));
	coreir_const #(
		.value(9'h1ff),
		.width(9)
	) const_511_9(.out(const_511_9_out));
	coreir_eq #(.width(16)) coreir_eq_16_inst0(
		.in0(tile_id),
		.in1(self_config_config_addr_out[15:0]),
		.out(coreir_eq_16_inst0_out)
	);
	wire [415:0] read_data_mux_I;
	assign read_data_mux_I[384+:32] = PowerDomainConfigReg_inst0_read_config_data;
	assign read_data_mux_I[352+:32] = SB_ID0_5TRACKS_B17_MemCore_read_config_data;
	assign read_data_mux_I[320+:32] = SB_ID0_5TRACKS_B1_MemCore_read_config_data;
	assign read_data_mux_I[288+:32] = CB_flush_read_config_data;
	assign read_data_mux_I[256+:32] = CB_MEM_input_width_1_num_1_read_config_data;
	assign read_data_mux_I[224+:32] = CB_MEM_input_width_1_num_0_read_config_data;
	assign read_data_mux_I[192+:32] = CB_MEM_input_width_17_num_3_read_config_data;
	assign read_data_mux_I[160+:32] = CB_MEM_input_width_17_num_2_read_config_data;
	assign read_data_mux_I[128+:32] = CB_MEM_input_width_17_num_1_read_config_data;
	assign read_data_mux_I[96+:32] = CB_MEM_input_width_17_num_0_read_config_data;
	assign read_data_mux_I[64+:32] = MemCore_inst0_read_config_data_2;
	assign read_data_mux_I[32+:32] = MemCore_inst0_read_config_data_1;
	assign read_data_mux_I[0+:32] = MemCore_inst0_read_config_data;
	MuxWithDefaultWrapper_13_32_8_0 read_data_mux(
		.I(read_data_mux_I),
		.S(self_config_config_addr_out[23:16]),
		.EN(and_inst0_out),
		.O(read_data_mux_O)
	);
	mantle_wire__typeBit32 self_config_config_addr(
		.in(config_config_addr),
		.out(self_config_config_addr_out)
	);
	assign SB_T0_EAST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T0_EAST_SB_IN_B17_ready_out;
	assign SB_T0_EAST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_IN_B1_ready_out;
	assign SB_T0_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_OUT_B1;
	assign SB_T0_EAST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T0_EAST_SB_OUT_B17;
	assign SB_T0_EAST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T0_EAST_SB_OUT_B17_valid_out;
	assign SB_T0_EAST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_OUT_B1_valid_out;
	assign SB_T0_NORTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T0_NORTH_SB_IN_B17_ready_out;
	assign SB_T0_NORTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_IN_B1_ready_out;
	assign SB_T0_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_OUT_B1;
	assign SB_T0_NORTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T0_NORTH_SB_OUT_B17;
	assign SB_T0_NORTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T0_NORTH_SB_OUT_B17_valid_out;
	assign SB_T0_NORTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_OUT_B1_valid_out;
	assign SB_T0_SOUTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T0_SOUTH_SB_IN_B17_ready_out;
	assign SB_T0_SOUTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_IN_B1_ready_out;
	assign SB_T0_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_OUT_B1;
	assign SB_T0_SOUTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T0_SOUTH_SB_OUT_B17;
	assign SB_T0_SOUTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T0_SOUTH_SB_OUT_B17_valid_out;
	assign SB_T0_SOUTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_OUT_B1_valid_out;
	assign SB_T0_WEST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T0_WEST_SB_IN_B17_ready_out;
	assign SB_T0_WEST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_IN_B1_ready_out;
	assign SB_T0_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_OUT_B1;
	assign SB_T0_WEST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T0_WEST_SB_OUT_B17;
	assign SB_T0_WEST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T0_WEST_SB_OUT_B17_valid_out;
	assign SB_T0_WEST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_OUT_B1_valid_out;
	assign SB_T1_EAST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T1_EAST_SB_IN_B17_ready_out;
	assign SB_T1_EAST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_IN_B1_ready_out;
	assign SB_T1_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_OUT_B1;
	assign SB_T1_EAST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T1_EAST_SB_OUT_B17;
	assign SB_T1_EAST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T1_EAST_SB_OUT_B17_valid_out;
	assign SB_T1_EAST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_OUT_B1_valid_out;
	assign SB_T1_NORTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T1_NORTH_SB_IN_B17_ready_out;
	assign SB_T1_NORTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_IN_B1_ready_out;
	assign SB_T1_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_OUT_B1;
	assign SB_T1_NORTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T1_NORTH_SB_OUT_B17;
	assign SB_T1_NORTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T1_NORTH_SB_OUT_B17_valid_out;
	assign SB_T1_NORTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_OUT_B1_valid_out;
	assign SB_T1_SOUTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T1_SOUTH_SB_IN_B17_ready_out;
	assign SB_T1_SOUTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_IN_B1_ready_out;
	assign SB_T1_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_OUT_B1;
	assign SB_T1_SOUTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T1_SOUTH_SB_OUT_B17;
	assign SB_T1_SOUTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T1_SOUTH_SB_OUT_B17_valid_out;
	assign SB_T1_SOUTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_OUT_B1_valid_out;
	assign SB_T1_WEST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T1_WEST_SB_IN_B17_ready_out;
	assign SB_T1_WEST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_IN_B1_ready_out;
	assign SB_T1_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_OUT_B1;
	assign SB_T1_WEST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T1_WEST_SB_OUT_B17;
	assign SB_T1_WEST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T1_WEST_SB_OUT_B17_valid_out;
	assign SB_T1_WEST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_OUT_B1_valid_out;
	assign SB_T2_EAST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T2_EAST_SB_IN_B17_ready_out;
	assign SB_T2_EAST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_IN_B1_ready_out;
	assign SB_T2_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_OUT_B1;
	assign SB_T2_EAST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T2_EAST_SB_OUT_B17;
	assign SB_T2_EAST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T2_EAST_SB_OUT_B17_valid_out;
	assign SB_T2_EAST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_OUT_B1_valid_out;
	assign SB_T2_NORTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T2_NORTH_SB_IN_B17_ready_out;
	assign SB_T2_NORTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_IN_B1_ready_out;
	assign SB_T2_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_OUT_B1;
	assign SB_T2_NORTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T2_NORTH_SB_OUT_B17;
	assign SB_T2_NORTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T2_NORTH_SB_OUT_B17_valid_out;
	assign SB_T2_NORTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_OUT_B1_valid_out;
	assign SB_T2_SOUTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T2_SOUTH_SB_IN_B17_ready_out;
	assign SB_T2_SOUTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_IN_B1_ready_out;
	assign SB_T2_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_OUT_B1;
	assign SB_T2_SOUTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T2_SOUTH_SB_OUT_B17;
	assign SB_T2_SOUTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T2_SOUTH_SB_OUT_B17_valid_out;
	assign SB_T2_SOUTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_OUT_B1_valid_out;
	assign SB_T2_WEST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T2_WEST_SB_IN_B17_ready_out;
	assign SB_T2_WEST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_IN_B1_ready_out;
	assign SB_T2_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_OUT_B1;
	assign SB_T2_WEST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T2_WEST_SB_OUT_B17;
	assign SB_T2_WEST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T2_WEST_SB_OUT_B17_valid_out;
	assign SB_T2_WEST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_OUT_B1_valid_out;
	assign SB_T3_EAST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T3_EAST_SB_IN_B17_ready_out;
	assign SB_T3_EAST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_IN_B1_ready_out;
	assign SB_T3_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_OUT_B1;
	assign SB_T3_EAST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T3_EAST_SB_OUT_B17;
	assign SB_T3_EAST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T3_EAST_SB_OUT_B17_valid_out;
	assign SB_T3_EAST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_OUT_B1_valid_out;
	assign SB_T3_NORTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T3_NORTH_SB_IN_B17_ready_out;
	assign SB_T3_NORTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_IN_B1_ready_out;
	assign SB_T3_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_OUT_B1;
	assign SB_T3_NORTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T3_NORTH_SB_OUT_B17;
	assign SB_T3_NORTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T3_NORTH_SB_OUT_B17_valid_out;
	assign SB_T3_NORTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_OUT_B1_valid_out;
	assign SB_T3_SOUTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T3_SOUTH_SB_IN_B17_ready_out;
	assign SB_T3_SOUTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_IN_B1_ready_out;
	assign SB_T3_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_OUT_B1;
	assign SB_T3_SOUTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T3_SOUTH_SB_OUT_B17;
	assign SB_T3_SOUTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T3_SOUTH_SB_OUT_B17_valid_out;
	assign SB_T3_SOUTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_OUT_B1_valid_out;
	assign SB_T3_WEST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T3_WEST_SB_IN_B17_ready_out;
	assign SB_T3_WEST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_IN_B1_ready_out;
	assign SB_T3_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_OUT_B1;
	assign SB_T3_WEST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T3_WEST_SB_OUT_B17;
	assign SB_T3_WEST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T3_WEST_SB_OUT_B17_valid_out;
	assign SB_T3_WEST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_OUT_B1_valid_out;
	assign SB_T4_EAST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T4_EAST_SB_IN_B17_ready_out;
	assign SB_T4_EAST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_IN_B1_ready_out;
	assign SB_T4_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_OUT_B1;
	assign SB_T4_EAST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T4_EAST_SB_OUT_B17;
	assign SB_T4_EAST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T4_EAST_SB_OUT_B17_valid_out;
	assign SB_T4_EAST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_OUT_B1_valid_out;
	assign SB_T4_NORTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T4_NORTH_SB_IN_B17_ready_out;
	assign SB_T4_NORTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_IN_B1_ready_out;
	assign SB_T4_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_OUT_B1;
	assign SB_T4_NORTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T4_NORTH_SB_OUT_B17;
	assign SB_T4_NORTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T4_NORTH_SB_OUT_B17_valid_out;
	assign SB_T4_NORTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_OUT_B1_valid_out;
	assign SB_T4_SOUTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T4_SOUTH_SB_IN_B17_ready_out;
	assign SB_T4_SOUTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_IN_B1_ready_out;
	assign SB_T4_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_OUT_B1;
	assign SB_T4_SOUTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T4_SOUTH_SB_OUT_B17;
	assign SB_T4_SOUTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T4_SOUTH_SB_OUT_B17_valid_out;
	assign SB_T4_SOUTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_OUT_B1_valid_out;
	assign SB_T4_WEST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T4_WEST_SB_IN_B17_ready_out;
	assign SB_T4_WEST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_IN_B1_ready_out;
	assign SB_T4_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_OUT_B1;
	assign SB_T4_WEST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T4_WEST_SB_OUT_B17;
	assign SB_T4_WEST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T4_WEST_SB_OUT_B17_valid_out;
	assign SB_T4_WEST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_OUT_B1_valid_out;
	assign clk_out = clk;
	assign config_out_config_addr = config_config_addr;
	assign config_out_config_data = config_config_data;
	assign config_out_read = config_read;
	assign config_out_write = config_write;
	assign flush_out = flush;
	assign hi = const_511_9_out;
	assign lo = const_0_8_out;
	assign read_config_data = PowerDomainOR_O;
	assign reset_out = reset;
	assign stall_out = stall;
endmodule
module Interconnect (
	clk,
	config_0_config_addr,
	config_0_config_data,
	config_0_read,
	config_0_write,
	config_1_config_addr,
	config_1_config_data,
	config_1_read,
	config_1_write,
	config_2_config_addr,
	config_2_config_data,
	config_2_read,
	config_2_write,
	config_3_config_addr,
	config_3_config_data,
	config_3_read,
	config_3_write,
	flush,
	glb2io_17_X00_Y00,
	glb2io_17_X00_Y00_ready,
	glb2io_17_X00_Y00_valid,
	glb2io_17_X01_Y00,
	glb2io_17_X01_Y00_ready,
	glb2io_17_X01_Y00_valid,
	glb2io_17_X02_Y00,
	glb2io_17_X02_Y00_ready,
	glb2io_17_X02_Y00_valid,
	glb2io_17_X03_Y00,
	glb2io_17_X03_Y00_ready,
	glb2io_17_X03_Y00_valid,
	glb2io_1_X00_Y00,
	glb2io_1_X00_Y00_ready,
	glb2io_1_X00_Y00_valid,
	glb2io_1_X01_Y00,
	glb2io_1_X01_Y00_ready,
	glb2io_1_X01_Y00_valid,
	glb2io_1_X02_Y00,
	glb2io_1_X02_Y00_ready,
	glb2io_1_X02_Y00_valid,
	glb2io_1_X03_Y00,
	glb2io_1_X03_Y00_ready,
	glb2io_1_X03_Y00_valid,
	io2glb_17_X00_Y00,
	io2glb_17_X00_Y00_ready,
	io2glb_17_X00_Y00_valid,
	io2glb_17_X01_Y00,
	io2glb_17_X01_Y00_ready,
	io2glb_17_X01_Y00_valid,
	io2glb_17_X02_Y00,
	io2glb_17_X02_Y00_ready,
	io2glb_17_X02_Y00_valid,
	io2glb_17_X03_Y00,
	io2glb_17_X03_Y00_ready,
	io2glb_17_X03_Y00_valid,
	io2glb_1_X00_Y00,
	io2glb_1_X00_Y00_ready,
	io2glb_1_X00_Y00_valid,
	io2glb_1_X01_Y00,
	io2glb_1_X01_Y00_ready,
	io2glb_1_X01_Y00_valid,
	io2glb_1_X02_Y00,
	io2glb_1_X02_Y00_ready,
	io2glb_1_X02_Y00_valid,
	io2glb_1_X03_Y00,
	io2glb_1_X03_Y00_ready,
	io2glb_1_X03_Y00_valid,
	read_config_data,
	reset,
	stall
);
	input clk;
	input [31:0] config_0_config_addr;
	input [31:0] config_0_config_data;
	input [0:0] config_0_read;
	input [0:0] config_0_write;
	input [31:0] config_1_config_addr;
	input [31:0] config_1_config_data;
	input [0:0] config_1_read;
	input [0:0] config_1_write;
	input [31:0] config_2_config_addr;
	input [31:0] config_2_config_data;
	input [0:0] config_2_read;
	input [0:0] config_2_write;
	input [31:0] config_3_config_addr;
	input [31:0] config_3_config_data;
	input [0:0] config_3_read;
	input [0:0] config_3_write;
	input [0:0] flush;
	input [16:0] glb2io_17_X00_Y00;
	output wire glb2io_17_X00_Y00_ready;
	input glb2io_17_X00_Y00_valid;
	input [16:0] glb2io_17_X01_Y00;
	output wire glb2io_17_X01_Y00_ready;
	input glb2io_17_X01_Y00_valid;
	input [16:0] glb2io_17_X02_Y00;
	output wire glb2io_17_X02_Y00_ready;
	input glb2io_17_X02_Y00_valid;
	input [16:0] glb2io_17_X03_Y00;
	output wire glb2io_17_X03_Y00_ready;
	input glb2io_17_X03_Y00_valid;
	input [0:0] glb2io_1_X00_Y00;
	output wire glb2io_1_X00_Y00_ready;
	input glb2io_1_X00_Y00_valid;
	input [0:0] glb2io_1_X01_Y00;
	output wire glb2io_1_X01_Y00_ready;
	input glb2io_1_X01_Y00_valid;
	input [0:0] glb2io_1_X02_Y00;
	output wire glb2io_1_X02_Y00_ready;
	input glb2io_1_X02_Y00_valid;
	input [0:0] glb2io_1_X03_Y00;
	output wire glb2io_1_X03_Y00_ready;
	input glb2io_1_X03_Y00_valid;
	output wire [16:0] io2glb_17_X00_Y00;
	input io2glb_17_X00_Y00_ready;
	output wire io2glb_17_X00_Y00_valid;
	output wire [16:0] io2glb_17_X01_Y00;
	input io2glb_17_X01_Y00_ready;
	output wire io2glb_17_X01_Y00_valid;
	output wire [16:0] io2glb_17_X02_Y00;
	input io2glb_17_X02_Y00_ready;
	output wire io2glb_17_X02_Y00_valid;
	output wire [16:0] io2glb_17_X03_Y00;
	input io2glb_17_X03_Y00_ready;
	output wire io2glb_17_X03_Y00_valid;
	output wire [0:0] io2glb_1_X00_Y00;
	input io2glb_1_X00_Y00_ready;
	output wire io2glb_1_X00_Y00_valid;
	output wire [0:0] io2glb_1_X01_Y00;
	input io2glb_1_X01_Y00_ready;
	output wire io2glb_1_X01_Y00_valid;
	output wire [0:0] io2glb_1_X02_Y00;
	input io2glb_1_X02_Y00_ready;
	output wire io2glb_1_X02_Y00_valid;
	output wire [0:0] io2glb_1_X03_Y00;
	input io2glb_1_X03_Y00_ready;
	output wire io2glb_1_X03_Y00_valid;
	output wire [31:0] read_config_data;
	input reset;
	input [3:0] stall;
	wire [0:0] PipelineRegister_inst0$Register_inst0$reg_P1_inst0_out;
	wire [0:0] PipelineRegister_inst1$Register_inst0$reg_P1_inst0_out;
	wire [0:0] PipelineRegister_inst2$Register_inst0$reg_P1_inst0_out;
	wire [0:0] PipelineRegister_inst3$Register_inst0$reg_P1_inst0_out;
	wire [65:0] PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out;
	wire [65:0] PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out;
	wire [65:0] PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out;
	wire [65:0] PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out;
	wire Tile_X00_Y00_clk_out;
	wire [31:0] Tile_X00_Y00_config_out_config_addr;
	wire [31:0] Tile_X00_Y00_config_out_config_data;
	wire [0:0] Tile_X00_Y00_config_out_read;
	wire [0:0] Tile_X00_Y00_config_out_write;
	wire Tile_X00_Y00_f2io_17_ready;
	wire Tile_X00_Y00_f2io_1_ready;
	wire [0:0] Tile_X00_Y00_flush_out;
	wire Tile_X00_Y00_glb2io_17_ready;
	wire Tile_X00_Y00_glb2io_1_ready;
	wire [8:0] Tile_X00_Y00_hi;
	wire [0:0] Tile_X00_Y00_io2f_1;
	wire [16:0] Tile_X00_Y00_io2f_17;
	wire Tile_X00_Y00_io2f_17_valid;
	wire Tile_X00_Y00_io2f_1_valid;
	wire [0:0] Tile_X00_Y00_io2glb_1;
	wire [16:0] Tile_X00_Y00_io2glb_17;
	wire Tile_X00_Y00_io2glb_17_valid;
	wire Tile_X00_Y00_io2glb_1_valid;
	wire [7:0] Tile_X00_Y00_lo;
	wire [31:0] Tile_X00_Y00_read_config_data;
	wire Tile_X00_Y00_reset_out;
	wire [0:0] Tile_X00_Y00_stall_out;
	wire Tile_X00_Y01_SB_T0_EAST_SB_IN_B17_ready;
	wire Tile_X00_Y01_SB_T0_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y01_SB_T0_EAST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y01_SB_T0_EAST_SB_OUT_B17;
	wire Tile_X00_Y01_SB_T0_EAST_SB_OUT_B17_valid;
	wire Tile_X00_Y01_SB_T0_EAST_SB_OUT_B1_valid;
	wire Tile_X00_Y01_SB_T0_NORTH_SB_IN_B17_ready;
	wire Tile_X00_Y01_SB_T0_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B17;
	wire Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B17_valid;
	wire Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B1_valid;
	wire Tile_X00_Y01_SB_T0_SOUTH_SB_IN_B17_ready;
	wire Tile_X00_Y01_SB_T0_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B17;
	wire Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B17_valid;
	wire Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B1_valid;
	wire Tile_X00_Y01_SB_T0_WEST_SB_IN_B17_ready;
	wire Tile_X00_Y01_SB_T0_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y01_SB_T0_WEST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y01_SB_T0_WEST_SB_OUT_B17;
	wire Tile_X00_Y01_SB_T0_WEST_SB_OUT_B17_valid;
	wire Tile_X00_Y01_SB_T0_WEST_SB_OUT_B1_valid;
	wire Tile_X00_Y01_SB_T1_EAST_SB_IN_B17_ready;
	wire Tile_X00_Y01_SB_T1_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y01_SB_T1_EAST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y01_SB_T1_EAST_SB_OUT_B17;
	wire Tile_X00_Y01_SB_T1_EAST_SB_OUT_B17_valid;
	wire Tile_X00_Y01_SB_T1_EAST_SB_OUT_B1_valid;
	wire Tile_X00_Y01_SB_T1_NORTH_SB_IN_B17_ready;
	wire Tile_X00_Y01_SB_T1_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y01_SB_T1_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y01_SB_T1_NORTH_SB_OUT_B17;
	wire Tile_X00_Y01_SB_T1_NORTH_SB_OUT_B17_valid;
	wire Tile_X00_Y01_SB_T1_NORTH_SB_OUT_B1_valid;
	wire Tile_X00_Y01_SB_T1_SOUTH_SB_IN_B17_ready;
	wire Tile_X00_Y01_SB_T1_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B17;
	wire Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B17_valid;
	wire Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B1_valid;
	wire Tile_X00_Y01_SB_T1_WEST_SB_IN_B17_ready;
	wire Tile_X00_Y01_SB_T1_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y01_SB_T1_WEST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y01_SB_T1_WEST_SB_OUT_B17;
	wire Tile_X00_Y01_SB_T1_WEST_SB_OUT_B17_valid;
	wire Tile_X00_Y01_SB_T1_WEST_SB_OUT_B1_valid;
	wire Tile_X00_Y01_SB_T2_EAST_SB_IN_B17_ready;
	wire Tile_X00_Y01_SB_T2_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y01_SB_T2_EAST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y01_SB_T2_EAST_SB_OUT_B17;
	wire Tile_X00_Y01_SB_T2_EAST_SB_OUT_B17_valid;
	wire Tile_X00_Y01_SB_T2_EAST_SB_OUT_B1_valid;
	wire Tile_X00_Y01_SB_T2_NORTH_SB_IN_B17_ready;
	wire Tile_X00_Y01_SB_T2_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y01_SB_T2_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y01_SB_T2_NORTH_SB_OUT_B17;
	wire Tile_X00_Y01_SB_T2_NORTH_SB_OUT_B17_valid;
	wire Tile_X00_Y01_SB_T2_NORTH_SB_OUT_B1_valid;
	wire Tile_X00_Y01_SB_T2_SOUTH_SB_IN_B17_ready;
	wire Tile_X00_Y01_SB_T2_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B17;
	wire Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B17_valid;
	wire Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B1_valid;
	wire Tile_X00_Y01_SB_T2_WEST_SB_IN_B17_ready;
	wire Tile_X00_Y01_SB_T2_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y01_SB_T2_WEST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y01_SB_T2_WEST_SB_OUT_B17;
	wire Tile_X00_Y01_SB_T2_WEST_SB_OUT_B17_valid;
	wire Tile_X00_Y01_SB_T2_WEST_SB_OUT_B1_valid;
	wire Tile_X00_Y01_SB_T3_EAST_SB_IN_B17_ready;
	wire Tile_X00_Y01_SB_T3_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y01_SB_T3_EAST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y01_SB_T3_EAST_SB_OUT_B17;
	wire Tile_X00_Y01_SB_T3_EAST_SB_OUT_B17_valid;
	wire Tile_X00_Y01_SB_T3_EAST_SB_OUT_B1_valid;
	wire Tile_X00_Y01_SB_T3_NORTH_SB_IN_B17_ready;
	wire Tile_X00_Y01_SB_T3_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y01_SB_T3_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y01_SB_T3_NORTH_SB_OUT_B17;
	wire Tile_X00_Y01_SB_T3_NORTH_SB_OUT_B17_valid;
	wire Tile_X00_Y01_SB_T3_NORTH_SB_OUT_B1_valid;
	wire Tile_X00_Y01_SB_T3_SOUTH_SB_IN_B17_ready;
	wire Tile_X00_Y01_SB_T3_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B17;
	wire Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B17_valid;
	wire Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B1_valid;
	wire Tile_X00_Y01_SB_T3_WEST_SB_IN_B17_ready;
	wire Tile_X00_Y01_SB_T3_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y01_SB_T3_WEST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y01_SB_T3_WEST_SB_OUT_B17;
	wire Tile_X00_Y01_SB_T3_WEST_SB_OUT_B17_valid;
	wire Tile_X00_Y01_SB_T3_WEST_SB_OUT_B1_valid;
	wire Tile_X00_Y01_SB_T4_EAST_SB_IN_B17_ready;
	wire Tile_X00_Y01_SB_T4_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y01_SB_T4_EAST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y01_SB_T4_EAST_SB_OUT_B17;
	wire Tile_X00_Y01_SB_T4_EAST_SB_OUT_B17_valid;
	wire Tile_X00_Y01_SB_T4_EAST_SB_OUT_B1_valid;
	wire Tile_X00_Y01_SB_T4_NORTH_SB_IN_B17_ready;
	wire Tile_X00_Y01_SB_T4_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y01_SB_T4_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y01_SB_T4_NORTH_SB_OUT_B17;
	wire Tile_X00_Y01_SB_T4_NORTH_SB_OUT_B17_valid;
	wire Tile_X00_Y01_SB_T4_NORTH_SB_OUT_B1_valid;
	wire Tile_X00_Y01_SB_T4_SOUTH_SB_IN_B17_ready;
	wire Tile_X00_Y01_SB_T4_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B17;
	wire Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B17_valid;
	wire Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B1_valid;
	wire Tile_X00_Y01_SB_T4_WEST_SB_IN_B17_ready;
	wire Tile_X00_Y01_SB_T4_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y01_SB_T4_WEST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y01_SB_T4_WEST_SB_OUT_B17;
	wire Tile_X00_Y01_SB_T4_WEST_SB_OUT_B17_valid;
	wire Tile_X00_Y01_SB_T4_WEST_SB_OUT_B1_valid;
	wire Tile_X00_Y01_clk_out;
	wire Tile_X00_Y01_clk_pass_through_out_bot;
	wire Tile_X00_Y01_clk_pass_through_out_right;
	wire [31:0] Tile_X00_Y01_config_out_config_addr;
	wire [31:0] Tile_X00_Y01_config_out_config_data;
	wire [0:0] Tile_X00_Y01_config_out_read;
	wire [0:0] Tile_X00_Y01_config_out_write;
	wire [0:0] Tile_X00_Y01_flush_out;
	wire [8:0] Tile_X00_Y01_hi;
	wire [7:0] Tile_X00_Y01_lo;
	wire [31:0] Tile_X00_Y01_read_config_data;
	wire Tile_X00_Y01_reset_out;
	wire [0:0] Tile_X00_Y01_stall_out;
	wire Tile_X00_Y02_SB_T0_EAST_SB_IN_B17_ready;
	wire Tile_X00_Y02_SB_T0_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y02_SB_T0_EAST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y02_SB_T0_EAST_SB_OUT_B17;
	wire Tile_X00_Y02_SB_T0_EAST_SB_OUT_B17_valid;
	wire Tile_X00_Y02_SB_T0_EAST_SB_OUT_B1_valid;
	wire Tile_X00_Y02_SB_T0_NORTH_SB_IN_B17_ready;
	wire Tile_X00_Y02_SB_T0_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B17;
	wire Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B17_valid;
	wire Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B1_valid;
	wire Tile_X00_Y02_SB_T0_SOUTH_SB_IN_B17_ready;
	wire Tile_X00_Y02_SB_T0_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B17;
	wire Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B17_valid;
	wire Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B1_valid;
	wire Tile_X00_Y02_SB_T0_WEST_SB_IN_B17_ready;
	wire Tile_X00_Y02_SB_T0_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y02_SB_T0_WEST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y02_SB_T0_WEST_SB_OUT_B17;
	wire Tile_X00_Y02_SB_T0_WEST_SB_OUT_B17_valid;
	wire Tile_X00_Y02_SB_T0_WEST_SB_OUT_B1_valid;
	wire Tile_X00_Y02_SB_T1_EAST_SB_IN_B17_ready;
	wire Tile_X00_Y02_SB_T1_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y02_SB_T1_EAST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y02_SB_T1_EAST_SB_OUT_B17;
	wire Tile_X00_Y02_SB_T1_EAST_SB_OUT_B17_valid;
	wire Tile_X00_Y02_SB_T1_EAST_SB_OUT_B1_valid;
	wire Tile_X00_Y02_SB_T1_NORTH_SB_IN_B17_ready;
	wire Tile_X00_Y02_SB_T1_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B17;
	wire Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B17_valid;
	wire Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B1_valid;
	wire Tile_X00_Y02_SB_T1_SOUTH_SB_IN_B17_ready;
	wire Tile_X00_Y02_SB_T1_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B17;
	wire Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B17_valid;
	wire Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B1_valid;
	wire Tile_X00_Y02_SB_T1_WEST_SB_IN_B17_ready;
	wire Tile_X00_Y02_SB_T1_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y02_SB_T1_WEST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y02_SB_T1_WEST_SB_OUT_B17;
	wire Tile_X00_Y02_SB_T1_WEST_SB_OUT_B17_valid;
	wire Tile_X00_Y02_SB_T1_WEST_SB_OUT_B1_valid;
	wire Tile_X00_Y02_SB_T2_EAST_SB_IN_B17_ready;
	wire Tile_X00_Y02_SB_T2_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y02_SB_T2_EAST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y02_SB_T2_EAST_SB_OUT_B17;
	wire Tile_X00_Y02_SB_T2_EAST_SB_OUT_B17_valid;
	wire Tile_X00_Y02_SB_T2_EAST_SB_OUT_B1_valid;
	wire Tile_X00_Y02_SB_T2_NORTH_SB_IN_B17_ready;
	wire Tile_X00_Y02_SB_T2_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B17;
	wire Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B17_valid;
	wire Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B1_valid;
	wire Tile_X00_Y02_SB_T2_SOUTH_SB_IN_B17_ready;
	wire Tile_X00_Y02_SB_T2_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B17;
	wire Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B17_valid;
	wire Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B1_valid;
	wire Tile_X00_Y02_SB_T2_WEST_SB_IN_B17_ready;
	wire Tile_X00_Y02_SB_T2_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y02_SB_T2_WEST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y02_SB_T2_WEST_SB_OUT_B17;
	wire Tile_X00_Y02_SB_T2_WEST_SB_OUT_B17_valid;
	wire Tile_X00_Y02_SB_T2_WEST_SB_OUT_B1_valid;
	wire Tile_X00_Y02_SB_T3_EAST_SB_IN_B17_ready;
	wire Tile_X00_Y02_SB_T3_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y02_SB_T3_EAST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y02_SB_T3_EAST_SB_OUT_B17;
	wire Tile_X00_Y02_SB_T3_EAST_SB_OUT_B17_valid;
	wire Tile_X00_Y02_SB_T3_EAST_SB_OUT_B1_valid;
	wire Tile_X00_Y02_SB_T3_NORTH_SB_IN_B17_ready;
	wire Tile_X00_Y02_SB_T3_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B17;
	wire Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B17_valid;
	wire Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B1_valid;
	wire Tile_X00_Y02_SB_T3_SOUTH_SB_IN_B17_ready;
	wire Tile_X00_Y02_SB_T3_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B17;
	wire Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B17_valid;
	wire Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B1_valid;
	wire Tile_X00_Y02_SB_T3_WEST_SB_IN_B17_ready;
	wire Tile_X00_Y02_SB_T3_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y02_SB_T3_WEST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y02_SB_T3_WEST_SB_OUT_B17;
	wire Tile_X00_Y02_SB_T3_WEST_SB_OUT_B17_valid;
	wire Tile_X00_Y02_SB_T3_WEST_SB_OUT_B1_valid;
	wire Tile_X00_Y02_SB_T4_EAST_SB_IN_B17_ready;
	wire Tile_X00_Y02_SB_T4_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y02_SB_T4_EAST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y02_SB_T4_EAST_SB_OUT_B17;
	wire Tile_X00_Y02_SB_T4_EAST_SB_OUT_B17_valid;
	wire Tile_X00_Y02_SB_T4_EAST_SB_OUT_B1_valid;
	wire Tile_X00_Y02_SB_T4_NORTH_SB_IN_B17_ready;
	wire Tile_X00_Y02_SB_T4_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B17;
	wire Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B17_valid;
	wire Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B1_valid;
	wire Tile_X00_Y02_SB_T4_SOUTH_SB_IN_B17_ready;
	wire Tile_X00_Y02_SB_T4_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B17;
	wire Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B17_valid;
	wire Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B1_valid;
	wire Tile_X00_Y02_SB_T4_WEST_SB_IN_B17_ready;
	wire Tile_X00_Y02_SB_T4_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y02_SB_T4_WEST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y02_SB_T4_WEST_SB_OUT_B17;
	wire Tile_X00_Y02_SB_T4_WEST_SB_OUT_B17_valid;
	wire Tile_X00_Y02_SB_T4_WEST_SB_OUT_B1_valid;
	wire Tile_X00_Y02_clk_out;
	wire Tile_X00_Y02_clk_pass_through_out_bot;
	wire Tile_X00_Y02_clk_pass_through_out_right;
	wire [31:0] Tile_X00_Y02_config_out_config_addr;
	wire [31:0] Tile_X00_Y02_config_out_config_data;
	wire [0:0] Tile_X00_Y02_config_out_read;
	wire [0:0] Tile_X00_Y02_config_out_write;
	wire [0:0] Tile_X00_Y02_flush_out;
	wire [8:0] Tile_X00_Y02_hi;
	wire [7:0] Tile_X00_Y02_lo;
	wire [31:0] Tile_X00_Y02_read_config_data;
	wire Tile_X00_Y02_reset_out;
	wire [0:0] Tile_X00_Y02_stall_out;
	wire Tile_X00_Y03_SB_T0_EAST_SB_IN_B17_ready;
	wire Tile_X00_Y03_SB_T0_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y03_SB_T0_EAST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y03_SB_T0_EAST_SB_OUT_B17;
	wire Tile_X00_Y03_SB_T0_EAST_SB_OUT_B17_valid;
	wire Tile_X00_Y03_SB_T0_EAST_SB_OUT_B1_valid;
	wire Tile_X00_Y03_SB_T0_NORTH_SB_IN_B17_ready;
	wire Tile_X00_Y03_SB_T0_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B17;
	wire Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B17_valid;
	wire Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B1_valid;
	wire Tile_X00_Y03_SB_T0_SOUTH_SB_IN_B17_ready;
	wire Tile_X00_Y03_SB_T0_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B17;
	wire Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B17_valid;
	wire Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B1_valid;
	wire Tile_X00_Y03_SB_T0_WEST_SB_IN_B17_ready;
	wire Tile_X00_Y03_SB_T0_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y03_SB_T0_WEST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y03_SB_T0_WEST_SB_OUT_B17;
	wire Tile_X00_Y03_SB_T0_WEST_SB_OUT_B17_valid;
	wire Tile_X00_Y03_SB_T0_WEST_SB_OUT_B1_valid;
	wire Tile_X00_Y03_SB_T1_EAST_SB_IN_B17_ready;
	wire Tile_X00_Y03_SB_T1_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y03_SB_T1_EAST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y03_SB_T1_EAST_SB_OUT_B17;
	wire Tile_X00_Y03_SB_T1_EAST_SB_OUT_B17_valid;
	wire Tile_X00_Y03_SB_T1_EAST_SB_OUT_B1_valid;
	wire Tile_X00_Y03_SB_T1_NORTH_SB_IN_B17_ready;
	wire Tile_X00_Y03_SB_T1_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B17;
	wire Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B17_valid;
	wire Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B1_valid;
	wire Tile_X00_Y03_SB_T1_SOUTH_SB_IN_B17_ready;
	wire Tile_X00_Y03_SB_T1_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B17;
	wire Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B17_valid;
	wire Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B1_valid;
	wire Tile_X00_Y03_SB_T1_WEST_SB_IN_B17_ready;
	wire Tile_X00_Y03_SB_T1_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y03_SB_T1_WEST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y03_SB_T1_WEST_SB_OUT_B17;
	wire Tile_X00_Y03_SB_T1_WEST_SB_OUT_B17_valid;
	wire Tile_X00_Y03_SB_T1_WEST_SB_OUT_B1_valid;
	wire Tile_X00_Y03_SB_T2_EAST_SB_IN_B17_ready;
	wire Tile_X00_Y03_SB_T2_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y03_SB_T2_EAST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y03_SB_T2_EAST_SB_OUT_B17;
	wire Tile_X00_Y03_SB_T2_EAST_SB_OUT_B17_valid;
	wire Tile_X00_Y03_SB_T2_EAST_SB_OUT_B1_valid;
	wire Tile_X00_Y03_SB_T2_NORTH_SB_IN_B17_ready;
	wire Tile_X00_Y03_SB_T2_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B17;
	wire Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B17_valid;
	wire Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B1_valid;
	wire Tile_X00_Y03_SB_T2_SOUTH_SB_IN_B17_ready;
	wire Tile_X00_Y03_SB_T2_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B17;
	wire Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B17_valid;
	wire Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B1_valid;
	wire Tile_X00_Y03_SB_T2_WEST_SB_IN_B17_ready;
	wire Tile_X00_Y03_SB_T2_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y03_SB_T2_WEST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y03_SB_T2_WEST_SB_OUT_B17;
	wire Tile_X00_Y03_SB_T2_WEST_SB_OUT_B17_valid;
	wire Tile_X00_Y03_SB_T2_WEST_SB_OUT_B1_valid;
	wire Tile_X00_Y03_SB_T3_EAST_SB_IN_B17_ready;
	wire Tile_X00_Y03_SB_T3_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y03_SB_T3_EAST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y03_SB_T3_EAST_SB_OUT_B17;
	wire Tile_X00_Y03_SB_T3_EAST_SB_OUT_B17_valid;
	wire Tile_X00_Y03_SB_T3_EAST_SB_OUT_B1_valid;
	wire Tile_X00_Y03_SB_T3_NORTH_SB_IN_B17_ready;
	wire Tile_X00_Y03_SB_T3_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B17;
	wire Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B17_valid;
	wire Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B1_valid;
	wire Tile_X00_Y03_SB_T3_SOUTH_SB_IN_B17_ready;
	wire Tile_X00_Y03_SB_T3_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B17;
	wire Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B17_valid;
	wire Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B1_valid;
	wire Tile_X00_Y03_SB_T3_WEST_SB_IN_B17_ready;
	wire Tile_X00_Y03_SB_T3_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y03_SB_T3_WEST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y03_SB_T3_WEST_SB_OUT_B17;
	wire Tile_X00_Y03_SB_T3_WEST_SB_OUT_B17_valid;
	wire Tile_X00_Y03_SB_T3_WEST_SB_OUT_B1_valid;
	wire Tile_X00_Y03_SB_T4_EAST_SB_IN_B17_ready;
	wire Tile_X00_Y03_SB_T4_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y03_SB_T4_EAST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y03_SB_T4_EAST_SB_OUT_B17;
	wire Tile_X00_Y03_SB_T4_EAST_SB_OUT_B17_valid;
	wire Tile_X00_Y03_SB_T4_EAST_SB_OUT_B1_valid;
	wire Tile_X00_Y03_SB_T4_NORTH_SB_IN_B17_ready;
	wire Tile_X00_Y03_SB_T4_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B17;
	wire Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B17_valid;
	wire Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B1_valid;
	wire Tile_X00_Y03_SB_T4_SOUTH_SB_IN_B17_ready;
	wire Tile_X00_Y03_SB_T4_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B17;
	wire Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B17_valid;
	wire Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B1_valid;
	wire Tile_X00_Y03_SB_T4_WEST_SB_IN_B17_ready;
	wire Tile_X00_Y03_SB_T4_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y03_SB_T4_WEST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y03_SB_T4_WEST_SB_OUT_B17;
	wire Tile_X00_Y03_SB_T4_WEST_SB_OUT_B17_valid;
	wire Tile_X00_Y03_SB_T4_WEST_SB_OUT_B1_valid;
	wire Tile_X00_Y03_clk_out;
	wire Tile_X00_Y03_clk_pass_through_out_bot;
	wire Tile_X00_Y03_clk_pass_through_out_right;
	wire [31:0] Tile_X00_Y03_config_out_config_addr;
	wire [31:0] Tile_X00_Y03_config_out_config_data;
	wire [0:0] Tile_X00_Y03_config_out_read;
	wire [0:0] Tile_X00_Y03_config_out_write;
	wire [0:0] Tile_X00_Y03_flush_out;
	wire [8:0] Tile_X00_Y03_hi;
	wire [7:0] Tile_X00_Y03_lo;
	wire [31:0] Tile_X00_Y03_read_config_data;
	wire Tile_X00_Y03_reset_out;
	wire [0:0] Tile_X00_Y03_stall_out;
	wire Tile_X00_Y04_SB_T0_EAST_SB_IN_B17_ready;
	wire Tile_X00_Y04_SB_T0_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y04_SB_T0_EAST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y04_SB_T0_EAST_SB_OUT_B17;
	wire Tile_X00_Y04_SB_T0_EAST_SB_OUT_B17_valid;
	wire Tile_X00_Y04_SB_T0_EAST_SB_OUT_B1_valid;
	wire Tile_X00_Y04_SB_T0_NORTH_SB_IN_B17_ready;
	wire Tile_X00_Y04_SB_T0_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B17;
	wire Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B17_valid;
	wire Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B1_valid;
	wire Tile_X00_Y04_SB_T0_SOUTH_SB_IN_B17_ready;
	wire Tile_X00_Y04_SB_T0_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B17;
	wire Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B17_valid;
	wire Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B1_valid;
	wire Tile_X00_Y04_SB_T0_WEST_SB_IN_B17_ready;
	wire Tile_X00_Y04_SB_T0_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y04_SB_T0_WEST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y04_SB_T0_WEST_SB_OUT_B17;
	wire Tile_X00_Y04_SB_T0_WEST_SB_OUT_B17_valid;
	wire Tile_X00_Y04_SB_T0_WEST_SB_OUT_B1_valid;
	wire Tile_X00_Y04_SB_T1_EAST_SB_IN_B17_ready;
	wire Tile_X00_Y04_SB_T1_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y04_SB_T1_EAST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y04_SB_T1_EAST_SB_OUT_B17;
	wire Tile_X00_Y04_SB_T1_EAST_SB_OUT_B17_valid;
	wire Tile_X00_Y04_SB_T1_EAST_SB_OUT_B1_valid;
	wire Tile_X00_Y04_SB_T1_NORTH_SB_IN_B17_ready;
	wire Tile_X00_Y04_SB_T1_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B17;
	wire Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B17_valid;
	wire Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B1_valid;
	wire Tile_X00_Y04_SB_T1_SOUTH_SB_IN_B17_ready;
	wire Tile_X00_Y04_SB_T1_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B17;
	wire Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B17_valid;
	wire Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B1_valid;
	wire Tile_X00_Y04_SB_T1_WEST_SB_IN_B17_ready;
	wire Tile_X00_Y04_SB_T1_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y04_SB_T1_WEST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y04_SB_T1_WEST_SB_OUT_B17;
	wire Tile_X00_Y04_SB_T1_WEST_SB_OUT_B17_valid;
	wire Tile_X00_Y04_SB_T1_WEST_SB_OUT_B1_valid;
	wire Tile_X00_Y04_SB_T2_EAST_SB_IN_B17_ready;
	wire Tile_X00_Y04_SB_T2_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y04_SB_T2_EAST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y04_SB_T2_EAST_SB_OUT_B17;
	wire Tile_X00_Y04_SB_T2_EAST_SB_OUT_B17_valid;
	wire Tile_X00_Y04_SB_T2_EAST_SB_OUT_B1_valid;
	wire Tile_X00_Y04_SB_T2_NORTH_SB_IN_B17_ready;
	wire Tile_X00_Y04_SB_T2_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B17;
	wire Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B17_valid;
	wire Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B1_valid;
	wire Tile_X00_Y04_SB_T2_SOUTH_SB_IN_B17_ready;
	wire Tile_X00_Y04_SB_T2_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B17;
	wire Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B17_valid;
	wire Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B1_valid;
	wire Tile_X00_Y04_SB_T2_WEST_SB_IN_B17_ready;
	wire Tile_X00_Y04_SB_T2_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y04_SB_T2_WEST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y04_SB_T2_WEST_SB_OUT_B17;
	wire Tile_X00_Y04_SB_T2_WEST_SB_OUT_B17_valid;
	wire Tile_X00_Y04_SB_T2_WEST_SB_OUT_B1_valid;
	wire Tile_X00_Y04_SB_T3_EAST_SB_IN_B17_ready;
	wire Tile_X00_Y04_SB_T3_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y04_SB_T3_EAST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y04_SB_T3_EAST_SB_OUT_B17;
	wire Tile_X00_Y04_SB_T3_EAST_SB_OUT_B17_valid;
	wire Tile_X00_Y04_SB_T3_EAST_SB_OUT_B1_valid;
	wire Tile_X00_Y04_SB_T3_NORTH_SB_IN_B17_ready;
	wire Tile_X00_Y04_SB_T3_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B17;
	wire Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B17_valid;
	wire Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B1_valid;
	wire Tile_X00_Y04_SB_T3_SOUTH_SB_IN_B17_ready;
	wire Tile_X00_Y04_SB_T3_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y04_SB_T3_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y04_SB_T3_SOUTH_SB_OUT_B17;
	wire Tile_X00_Y04_SB_T3_SOUTH_SB_OUT_B17_valid;
	wire Tile_X00_Y04_SB_T3_SOUTH_SB_OUT_B1_valid;
	wire Tile_X00_Y04_SB_T3_WEST_SB_IN_B17_ready;
	wire Tile_X00_Y04_SB_T3_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y04_SB_T3_WEST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y04_SB_T3_WEST_SB_OUT_B17;
	wire Tile_X00_Y04_SB_T3_WEST_SB_OUT_B17_valid;
	wire Tile_X00_Y04_SB_T3_WEST_SB_OUT_B1_valid;
	wire Tile_X00_Y04_SB_T4_EAST_SB_IN_B17_ready;
	wire Tile_X00_Y04_SB_T4_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y04_SB_T4_EAST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y04_SB_T4_EAST_SB_OUT_B17;
	wire Tile_X00_Y04_SB_T4_EAST_SB_OUT_B17_valid;
	wire Tile_X00_Y04_SB_T4_EAST_SB_OUT_B1_valid;
	wire Tile_X00_Y04_SB_T4_NORTH_SB_IN_B17_ready;
	wire Tile_X00_Y04_SB_T4_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B17;
	wire Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B17_valid;
	wire Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B1_valid;
	wire Tile_X00_Y04_SB_T4_SOUTH_SB_IN_B17_ready;
	wire Tile_X00_Y04_SB_T4_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y04_SB_T4_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X00_Y04_SB_T4_SOUTH_SB_OUT_B17;
	wire Tile_X00_Y04_SB_T4_SOUTH_SB_OUT_B17_valid;
	wire Tile_X00_Y04_SB_T4_SOUTH_SB_OUT_B1_valid;
	wire Tile_X00_Y04_SB_T4_WEST_SB_IN_B17_ready;
	wire Tile_X00_Y04_SB_T4_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X00_Y04_SB_T4_WEST_SB_OUT_B1;
	wire [16:0] Tile_X00_Y04_SB_T4_WEST_SB_OUT_B17;
	wire Tile_X00_Y04_SB_T4_WEST_SB_OUT_B17_valid;
	wire Tile_X00_Y04_SB_T4_WEST_SB_OUT_B1_valid;
	wire Tile_X00_Y04_clk_out;
	wire Tile_X00_Y04_clk_pass_through_out_bot;
	wire Tile_X00_Y04_clk_pass_through_out_right;
	wire [31:0] Tile_X00_Y04_config_out_config_addr;
	wire [31:0] Tile_X00_Y04_config_out_config_data;
	wire [0:0] Tile_X00_Y04_config_out_read;
	wire [0:0] Tile_X00_Y04_config_out_write;
	wire [0:0] Tile_X00_Y04_flush_out;
	wire [8:0] Tile_X00_Y04_hi;
	wire [7:0] Tile_X00_Y04_lo;
	wire [31:0] Tile_X00_Y04_read_config_data;
	wire Tile_X00_Y04_reset_out;
	wire [0:0] Tile_X00_Y04_stall_out;
	wire Tile_X01_Y00_clk_out;
	wire [31:0] Tile_X01_Y00_config_out_config_addr;
	wire [31:0] Tile_X01_Y00_config_out_config_data;
	wire [0:0] Tile_X01_Y00_config_out_read;
	wire [0:0] Tile_X01_Y00_config_out_write;
	wire Tile_X01_Y00_f2io_17_ready;
	wire Tile_X01_Y00_f2io_1_ready;
	wire [0:0] Tile_X01_Y00_flush_out;
	wire Tile_X01_Y00_glb2io_17_ready;
	wire Tile_X01_Y00_glb2io_1_ready;
	wire [8:0] Tile_X01_Y00_hi;
	wire [0:0] Tile_X01_Y00_io2f_1;
	wire [16:0] Tile_X01_Y00_io2f_17;
	wire Tile_X01_Y00_io2f_17_valid;
	wire Tile_X01_Y00_io2f_1_valid;
	wire [0:0] Tile_X01_Y00_io2glb_1;
	wire [16:0] Tile_X01_Y00_io2glb_17;
	wire Tile_X01_Y00_io2glb_17_valid;
	wire Tile_X01_Y00_io2glb_1_valid;
	wire [7:0] Tile_X01_Y00_lo;
	wire [31:0] Tile_X01_Y00_read_config_data;
	wire Tile_X01_Y00_reset_out;
	wire [0:0] Tile_X01_Y00_stall_out;
	wire Tile_X01_Y01_SB_T0_EAST_SB_IN_B17_ready;
	wire Tile_X01_Y01_SB_T0_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y01_SB_T0_EAST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y01_SB_T0_EAST_SB_OUT_B17;
	wire Tile_X01_Y01_SB_T0_EAST_SB_OUT_B17_valid;
	wire Tile_X01_Y01_SB_T0_EAST_SB_OUT_B1_valid;
	wire Tile_X01_Y01_SB_T0_NORTH_SB_IN_B17_ready;
	wire Tile_X01_Y01_SB_T0_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B17;
	wire Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B17_valid;
	wire Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B1_valid;
	wire Tile_X01_Y01_SB_T0_SOUTH_SB_IN_B17_ready;
	wire Tile_X01_Y01_SB_T0_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B17;
	wire Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B17_valid;
	wire Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B1_valid;
	wire Tile_X01_Y01_SB_T0_WEST_SB_IN_B17_ready;
	wire Tile_X01_Y01_SB_T0_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y01_SB_T0_WEST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y01_SB_T0_WEST_SB_OUT_B17;
	wire Tile_X01_Y01_SB_T0_WEST_SB_OUT_B17_valid;
	wire Tile_X01_Y01_SB_T0_WEST_SB_OUT_B1_valid;
	wire Tile_X01_Y01_SB_T1_EAST_SB_IN_B17_ready;
	wire Tile_X01_Y01_SB_T1_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y01_SB_T1_EAST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y01_SB_T1_EAST_SB_OUT_B17;
	wire Tile_X01_Y01_SB_T1_EAST_SB_OUT_B17_valid;
	wire Tile_X01_Y01_SB_T1_EAST_SB_OUT_B1_valid;
	wire Tile_X01_Y01_SB_T1_NORTH_SB_IN_B17_ready;
	wire Tile_X01_Y01_SB_T1_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y01_SB_T1_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y01_SB_T1_NORTH_SB_OUT_B17;
	wire Tile_X01_Y01_SB_T1_NORTH_SB_OUT_B17_valid;
	wire Tile_X01_Y01_SB_T1_NORTH_SB_OUT_B1_valid;
	wire Tile_X01_Y01_SB_T1_SOUTH_SB_IN_B17_ready;
	wire Tile_X01_Y01_SB_T1_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B17;
	wire Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B17_valid;
	wire Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B1_valid;
	wire Tile_X01_Y01_SB_T1_WEST_SB_IN_B17_ready;
	wire Tile_X01_Y01_SB_T1_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y01_SB_T1_WEST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y01_SB_T1_WEST_SB_OUT_B17;
	wire Tile_X01_Y01_SB_T1_WEST_SB_OUT_B17_valid;
	wire Tile_X01_Y01_SB_T1_WEST_SB_OUT_B1_valid;
	wire Tile_X01_Y01_SB_T2_EAST_SB_IN_B17_ready;
	wire Tile_X01_Y01_SB_T2_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y01_SB_T2_EAST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y01_SB_T2_EAST_SB_OUT_B17;
	wire Tile_X01_Y01_SB_T2_EAST_SB_OUT_B17_valid;
	wire Tile_X01_Y01_SB_T2_EAST_SB_OUT_B1_valid;
	wire Tile_X01_Y01_SB_T2_NORTH_SB_IN_B17_ready;
	wire Tile_X01_Y01_SB_T2_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y01_SB_T2_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y01_SB_T2_NORTH_SB_OUT_B17;
	wire Tile_X01_Y01_SB_T2_NORTH_SB_OUT_B17_valid;
	wire Tile_X01_Y01_SB_T2_NORTH_SB_OUT_B1_valid;
	wire Tile_X01_Y01_SB_T2_SOUTH_SB_IN_B17_ready;
	wire Tile_X01_Y01_SB_T2_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B17;
	wire Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B17_valid;
	wire Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B1_valid;
	wire Tile_X01_Y01_SB_T2_WEST_SB_IN_B17_ready;
	wire Tile_X01_Y01_SB_T2_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y01_SB_T2_WEST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y01_SB_T2_WEST_SB_OUT_B17;
	wire Tile_X01_Y01_SB_T2_WEST_SB_OUT_B17_valid;
	wire Tile_X01_Y01_SB_T2_WEST_SB_OUT_B1_valid;
	wire Tile_X01_Y01_SB_T3_EAST_SB_IN_B17_ready;
	wire Tile_X01_Y01_SB_T3_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y01_SB_T3_EAST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y01_SB_T3_EAST_SB_OUT_B17;
	wire Tile_X01_Y01_SB_T3_EAST_SB_OUT_B17_valid;
	wire Tile_X01_Y01_SB_T3_EAST_SB_OUT_B1_valid;
	wire Tile_X01_Y01_SB_T3_NORTH_SB_IN_B17_ready;
	wire Tile_X01_Y01_SB_T3_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y01_SB_T3_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y01_SB_T3_NORTH_SB_OUT_B17;
	wire Tile_X01_Y01_SB_T3_NORTH_SB_OUT_B17_valid;
	wire Tile_X01_Y01_SB_T3_NORTH_SB_OUT_B1_valid;
	wire Tile_X01_Y01_SB_T3_SOUTH_SB_IN_B17_ready;
	wire Tile_X01_Y01_SB_T3_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B17;
	wire Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B17_valid;
	wire Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B1_valid;
	wire Tile_X01_Y01_SB_T3_WEST_SB_IN_B17_ready;
	wire Tile_X01_Y01_SB_T3_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y01_SB_T3_WEST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y01_SB_T3_WEST_SB_OUT_B17;
	wire Tile_X01_Y01_SB_T3_WEST_SB_OUT_B17_valid;
	wire Tile_X01_Y01_SB_T3_WEST_SB_OUT_B1_valid;
	wire Tile_X01_Y01_SB_T4_EAST_SB_IN_B17_ready;
	wire Tile_X01_Y01_SB_T4_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y01_SB_T4_EAST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y01_SB_T4_EAST_SB_OUT_B17;
	wire Tile_X01_Y01_SB_T4_EAST_SB_OUT_B17_valid;
	wire Tile_X01_Y01_SB_T4_EAST_SB_OUT_B1_valid;
	wire Tile_X01_Y01_SB_T4_NORTH_SB_IN_B17_ready;
	wire Tile_X01_Y01_SB_T4_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y01_SB_T4_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y01_SB_T4_NORTH_SB_OUT_B17;
	wire Tile_X01_Y01_SB_T4_NORTH_SB_OUT_B17_valid;
	wire Tile_X01_Y01_SB_T4_NORTH_SB_OUT_B1_valid;
	wire Tile_X01_Y01_SB_T4_SOUTH_SB_IN_B17_ready;
	wire Tile_X01_Y01_SB_T4_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B17;
	wire Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B17_valid;
	wire Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B1_valid;
	wire Tile_X01_Y01_SB_T4_WEST_SB_IN_B17_ready;
	wire Tile_X01_Y01_SB_T4_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y01_SB_T4_WEST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y01_SB_T4_WEST_SB_OUT_B17;
	wire Tile_X01_Y01_SB_T4_WEST_SB_OUT_B17_valid;
	wire Tile_X01_Y01_SB_T4_WEST_SB_OUT_B1_valid;
	wire Tile_X01_Y01_clk_out;
	wire Tile_X01_Y01_clk_pass_through_out_bot;
	wire Tile_X01_Y01_clk_pass_through_out_right;
	wire [31:0] Tile_X01_Y01_config_out_config_addr;
	wire [31:0] Tile_X01_Y01_config_out_config_data;
	wire [0:0] Tile_X01_Y01_config_out_read;
	wire [0:0] Tile_X01_Y01_config_out_write;
	wire [0:0] Tile_X01_Y01_flush_out;
	wire [8:0] Tile_X01_Y01_hi;
	wire [7:0] Tile_X01_Y01_lo;
	wire [31:0] Tile_X01_Y01_read_config_data;
	wire Tile_X01_Y01_reset_out;
	wire [0:0] Tile_X01_Y01_stall_out;
	wire Tile_X01_Y02_SB_T0_EAST_SB_IN_B17_ready;
	wire Tile_X01_Y02_SB_T0_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y02_SB_T0_EAST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y02_SB_T0_EAST_SB_OUT_B17;
	wire Tile_X01_Y02_SB_T0_EAST_SB_OUT_B17_valid;
	wire Tile_X01_Y02_SB_T0_EAST_SB_OUT_B1_valid;
	wire Tile_X01_Y02_SB_T0_NORTH_SB_IN_B17_ready;
	wire Tile_X01_Y02_SB_T0_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B17;
	wire Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B17_valid;
	wire Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B1_valid;
	wire Tile_X01_Y02_SB_T0_SOUTH_SB_IN_B17_ready;
	wire Tile_X01_Y02_SB_T0_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B17;
	wire Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B17_valid;
	wire Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B1_valid;
	wire Tile_X01_Y02_SB_T0_WEST_SB_IN_B17_ready;
	wire Tile_X01_Y02_SB_T0_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y02_SB_T0_WEST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y02_SB_T0_WEST_SB_OUT_B17;
	wire Tile_X01_Y02_SB_T0_WEST_SB_OUT_B17_valid;
	wire Tile_X01_Y02_SB_T0_WEST_SB_OUT_B1_valid;
	wire Tile_X01_Y02_SB_T1_EAST_SB_IN_B17_ready;
	wire Tile_X01_Y02_SB_T1_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y02_SB_T1_EAST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y02_SB_T1_EAST_SB_OUT_B17;
	wire Tile_X01_Y02_SB_T1_EAST_SB_OUT_B17_valid;
	wire Tile_X01_Y02_SB_T1_EAST_SB_OUT_B1_valid;
	wire Tile_X01_Y02_SB_T1_NORTH_SB_IN_B17_ready;
	wire Tile_X01_Y02_SB_T1_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B17;
	wire Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B17_valid;
	wire Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B1_valid;
	wire Tile_X01_Y02_SB_T1_SOUTH_SB_IN_B17_ready;
	wire Tile_X01_Y02_SB_T1_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B17;
	wire Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B17_valid;
	wire Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B1_valid;
	wire Tile_X01_Y02_SB_T1_WEST_SB_IN_B17_ready;
	wire Tile_X01_Y02_SB_T1_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y02_SB_T1_WEST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y02_SB_T1_WEST_SB_OUT_B17;
	wire Tile_X01_Y02_SB_T1_WEST_SB_OUT_B17_valid;
	wire Tile_X01_Y02_SB_T1_WEST_SB_OUT_B1_valid;
	wire Tile_X01_Y02_SB_T2_EAST_SB_IN_B17_ready;
	wire Tile_X01_Y02_SB_T2_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y02_SB_T2_EAST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y02_SB_T2_EAST_SB_OUT_B17;
	wire Tile_X01_Y02_SB_T2_EAST_SB_OUT_B17_valid;
	wire Tile_X01_Y02_SB_T2_EAST_SB_OUT_B1_valid;
	wire Tile_X01_Y02_SB_T2_NORTH_SB_IN_B17_ready;
	wire Tile_X01_Y02_SB_T2_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B17;
	wire Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B17_valid;
	wire Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B1_valid;
	wire Tile_X01_Y02_SB_T2_SOUTH_SB_IN_B17_ready;
	wire Tile_X01_Y02_SB_T2_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B17;
	wire Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B17_valid;
	wire Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B1_valid;
	wire Tile_X01_Y02_SB_T2_WEST_SB_IN_B17_ready;
	wire Tile_X01_Y02_SB_T2_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y02_SB_T2_WEST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y02_SB_T2_WEST_SB_OUT_B17;
	wire Tile_X01_Y02_SB_T2_WEST_SB_OUT_B17_valid;
	wire Tile_X01_Y02_SB_T2_WEST_SB_OUT_B1_valid;
	wire Tile_X01_Y02_SB_T3_EAST_SB_IN_B17_ready;
	wire Tile_X01_Y02_SB_T3_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y02_SB_T3_EAST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y02_SB_T3_EAST_SB_OUT_B17;
	wire Tile_X01_Y02_SB_T3_EAST_SB_OUT_B17_valid;
	wire Tile_X01_Y02_SB_T3_EAST_SB_OUT_B1_valid;
	wire Tile_X01_Y02_SB_T3_NORTH_SB_IN_B17_ready;
	wire Tile_X01_Y02_SB_T3_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B17;
	wire Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B17_valid;
	wire Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B1_valid;
	wire Tile_X01_Y02_SB_T3_SOUTH_SB_IN_B17_ready;
	wire Tile_X01_Y02_SB_T3_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B17;
	wire Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B17_valid;
	wire Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B1_valid;
	wire Tile_X01_Y02_SB_T3_WEST_SB_IN_B17_ready;
	wire Tile_X01_Y02_SB_T3_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y02_SB_T3_WEST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y02_SB_T3_WEST_SB_OUT_B17;
	wire Tile_X01_Y02_SB_T3_WEST_SB_OUT_B17_valid;
	wire Tile_X01_Y02_SB_T3_WEST_SB_OUT_B1_valid;
	wire Tile_X01_Y02_SB_T4_EAST_SB_IN_B17_ready;
	wire Tile_X01_Y02_SB_T4_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y02_SB_T4_EAST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y02_SB_T4_EAST_SB_OUT_B17;
	wire Tile_X01_Y02_SB_T4_EAST_SB_OUT_B17_valid;
	wire Tile_X01_Y02_SB_T4_EAST_SB_OUT_B1_valid;
	wire Tile_X01_Y02_SB_T4_NORTH_SB_IN_B17_ready;
	wire Tile_X01_Y02_SB_T4_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B17;
	wire Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B17_valid;
	wire Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B1_valid;
	wire Tile_X01_Y02_SB_T4_SOUTH_SB_IN_B17_ready;
	wire Tile_X01_Y02_SB_T4_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B17;
	wire Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B17_valid;
	wire Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B1_valid;
	wire Tile_X01_Y02_SB_T4_WEST_SB_IN_B17_ready;
	wire Tile_X01_Y02_SB_T4_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y02_SB_T4_WEST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y02_SB_T4_WEST_SB_OUT_B17;
	wire Tile_X01_Y02_SB_T4_WEST_SB_OUT_B17_valid;
	wire Tile_X01_Y02_SB_T4_WEST_SB_OUT_B1_valid;
	wire Tile_X01_Y02_clk_out;
	wire Tile_X01_Y02_clk_pass_through_out_bot;
	wire Tile_X01_Y02_clk_pass_through_out_right;
	wire [31:0] Tile_X01_Y02_config_out_config_addr;
	wire [31:0] Tile_X01_Y02_config_out_config_data;
	wire [0:0] Tile_X01_Y02_config_out_read;
	wire [0:0] Tile_X01_Y02_config_out_write;
	wire [0:0] Tile_X01_Y02_flush_out;
	wire [8:0] Tile_X01_Y02_hi;
	wire [7:0] Tile_X01_Y02_lo;
	wire [31:0] Tile_X01_Y02_read_config_data;
	wire Tile_X01_Y02_reset_out;
	wire [0:0] Tile_X01_Y02_stall_out;
	wire Tile_X01_Y03_SB_T0_EAST_SB_IN_B17_ready;
	wire Tile_X01_Y03_SB_T0_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y03_SB_T0_EAST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y03_SB_T0_EAST_SB_OUT_B17;
	wire Tile_X01_Y03_SB_T0_EAST_SB_OUT_B17_valid;
	wire Tile_X01_Y03_SB_T0_EAST_SB_OUT_B1_valid;
	wire Tile_X01_Y03_SB_T0_NORTH_SB_IN_B17_ready;
	wire Tile_X01_Y03_SB_T0_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B17;
	wire Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B17_valid;
	wire Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B1_valid;
	wire Tile_X01_Y03_SB_T0_SOUTH_SB_IN_B17_ready;
	wire Tile_X01_Y03_SB_T0_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B17;
	wire Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B17_valid;
	wire Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B1_valid;
	wire Tile_X01_Y03_SB_T0_WEST_SB_IN_B17_ready;
	wire Tile_X01_Y03_SB_T0_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y03_SB_T0_WEST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y03_SB_T0_WEST_SB_OUT_B17;
	wire Tile_X01_Y03_SB_T0_WEST_SB_OUT_B17_valid;
	wire Tile_X01_Y03_SB_T0_WEST_SB_OUT_B1_valid;
	wire Tile_X01_Y03_SB_T1_EAST_SB_IN_B17_ready;
	wire Tile_X01_Y03_SB_T1_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y03_SB_T1_EAST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y03_SB_T1_EAST_SB_OUT_B17;
	wire Tile_X01_Y03_SB_T1_EAST_SB_OUT_B17_valid;
	wire Tile_X01_Y03_SB_T1_EAST_SB_OUT_B1_valid;
	wire Tile_X01_Y03_SB_T1_NORTH_SB_IN_B17_ready;
	wire Tile_X01_Y03_SB_T1_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B17;
	wire Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B17_valid;
	wire Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B1_valid;
	wire Tile_X01_Y03_SB_T1_SOUTH_SB_IN_B17_ready;
	wire Tile_X01_Y03_SB_T1_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B17;
	wire Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B17_valid;
	wire Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B1_valid;
	wire Tile_X01_Y03_SB_T1_WEST_SB_IN_B17_ready;
	wire Tile_X01_Y03_SB_T1_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y03_SB_T1_WEST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y03_SB_T1_WEST_SB_OUT_B17;
	wire Tile_X01_Y03_SB_T1_WEST_SB_OUT_B17_valid;
	wire Tile_X01_Y03_SB_T1_WEST_SB_OUT_B1_valid;
	wire Tile_X01_Y03_SB_T2_EAST_SB_IN_B17_ready;
	wire Tile_X01_Y03_SB_T2_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y03_SB_T2_EAST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y03_SB_T2_EAST_SB_OUT_B17;
	wire Tile_X01_Y03_SB_T2_EAST_SB_OUT_B17_valid;
	wire Tile_X01_Y03_SB_T2_EAST_SB_OUT_B1_valid;
	wire Tile_X01_Y03_SB_T2_NORTH_SB_IN_B17_ready;
	wire Tile_X01_Y03_SB_T2_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B17;
	wire Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B17_valid;
	wire Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B1_valid;
	wire Tile_X01_Y03_SB_T2_SOUTH_SB_IN_B17_ready;
	wire Tile_X01_Y03_SB_T2_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B17;
	wire Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B17_valid;
	wire Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B1_valid;
	wire Tile_X01_Y03_SB_T2_WEST_SB_IN_B17_ready;
	wire Tile_X01_Y03_SB_T2_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y03_SB_T2_WEST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y03_SB_T2_WEST_SB_OUT_B17;
	wire Tile_X01_Y03_SB_T2_WEST_SB_OUT_B17_valid;
	wire Tile_X01_Y03_SB_T2_WEST_SB_OUT_B1_valid;
	wire Tile_X01_Y03_SB_T3_EAST_SB_IN_B17_ready;
	wire Tile_X01_Y03_SB_T3_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y03_SB_T3_EAST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y03_SB_T3_EAST_SB_OUT_B17;
	wire Tile_X01_Y03_SB_T3_EAST_SB_OUT_B17_valid;
	wire Tile_X01_Y03_SB_T3_EAST_SB_OUT_B1_valid;
	wire Tile_X01_Y03_SB_T3_NORTH_SB_IN_B17_ready;
	wire Tile_X01_Y03_SB_T3_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B17;
	wire Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B17_valid;
	wire Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B1_valid;
	wire Tile_X01_Y03_SB_T3_SOUTH_SB_IN_B17_ready;
	wire Tile_X01_Y03_SB_T3_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B17;
	wire Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B17_valid;
	wire Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B1_valid;
	wire Tile_X01_Y03_SB_T3_WEST_SB_IN_B17_ready;
	wire Tile_X01_Y03_SB_T3_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y03_SB_T3_WEST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y03_SB_T3_WEST_SB_OUT_B17;
	wire Tile_X01_Y03_SB_T3_WEST_SB_OUT_B17_valid;
	wire Tile_X01_Y03_SB_T3_WEST_SB_OUT_B1_valid;
	wire Tile_X01_Y03_SB_T4_EAST_SB_IN_B17_ready;
	wire Tile_X01_Y03_SB_T4_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y03_SB_T4_EAST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y03_SB_T4_EAST_SB_OUT_B17;
	wire Tile_X01_Y03_SB_T4_EAST_SB_OUT_B17_valid;
	wire Tile_X01_Y03_SB_T4_EAST_SB_OUT_B1_valid;
	wire Tile_X01_Y03_SB_T4_NORTH_SB_IN_B17_ready;
	wire Tile_X01_Y03_SB_T4_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B17;
	wire Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B17_valid;
	wire Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B1_valid;
	wire Tile_X01_Y03_SB_T4_SOUTH_SB_IN_B17_ready;
	wire Tile_X01_Y03_SB_T4_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B17;
	wire Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B17_valid;
	wire Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B1_valid;
	wire Tile_X01_Y03_SB_T4_WEST_SB_IN_B17_ready;
	wire Tile_X01_Y03_SB_T4_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y03_SB_T4_WEST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y03_SB_T4_WEST_SB_OUT_B17;
	wire Tile_X01_Y03_SB_T4_WEST_SB_OUT_B17_valid;
	wire Tile_X01_Y03_SB_T4_WEST_SB_OUT_B1_valid;
	wire Tile_X01_Y03_clk_out;
	wire Tile_X01_Y03_clk_pass_through_out_bot;
	wire Tile_X01_Y03_clk_pass_through_out_right;
	wire [31:0] Tile_X01_Y03_config_out_config_addr;
	wire [31:0] Tile_X01_Y03_config_out_config_data;
	wire [0:0] Tile_X01_Y03_config_out_read;
	wire [0:0] Tile_X01_Y03_config_out_write;
	wire [0:0] Tile_X01_Y03_flush_out;
	wire [8:0] Tile_X01_Y03_hi;
	wire [7:0] Tile_X01_Y03_lo;
	wire [31:0] Tile_X01_Y03_read_config_data;
	wire Tile_X01_Y03_reset_out;
	wire [0:0] Tile_X01_Y03_stall_out;
	wire Tile_X01_Y04_SB_T0_EAST_SB_IN_B17_ready;
	wire Tile_X01_Y04_SB_T0_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y04_SB_T0_EAST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y04_SB_T0_EAST_SB_OUT_B17;
	wire Tile_X01_Y04_SB_T0_EAST_SB_OUT_B17_valid;
	wire Tile_X01_Y04_SB_T0_EAST_SB_OUT_B1_valid;
	wire Tile_X01_Y04_SB_T0_NORTH_SB_IN_B17_ready;
	wire Tile_X01_Y04_SB_T0_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B17;
	wire Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B17_valid;
	wire Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B1_valid;
	wire Tile_X01_Y04_SB_T0_SOUTH_SB_IN_B17_ready;
	wire Tile_X01_Y04_SB_T0_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B17;
	wire Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B17_valid;
	wire Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B1_valid;
	wire Tile_X01_Y04_SB_T0_WEST_SB_IN_B17_ready;
	wire Tile_X01_Y04_SB_T0_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y04_SB_T0_WEST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y04_SB_T0_WEST_SB_OUT_B17;
	wire Tile_X01_Y04_SB_T0_WEST_SB_OUT_B17_valid;
	wire Tile_X01_Y04_SB_T0_WEST_SB_OUT_B1_valid;
	wire Tile_X01_Y04_SB_T1_EAST_SB_IN_B17_ready;
	wire Tile_X01_Y04_SB_T1_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y04_SB_T1_EAST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y04_SB_T1_EAST_SB_OUT_B17;
	wire Tile_X01_Y04_SB_T1_EAST_SB_OUT_B17_valid;
	wire Tile_X01_Y04_SB_T1_EAST_SB_OUT_B1_valid;
	wire Tile_X01_Y04_SB_T1_NORTH_SB_IN_B17_ready;
	wire Tile_X01_Y04_SB_T1_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B17;
	wire Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B17_valid;
	wire Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B1_valid;
	wire Tile_X01_Y04_SB_T1_SOUTH_SB_IN_B17_ready;
	wire Tile_X01_Y04_SB_T1_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B17;
	wire Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B17_valid;
	wire Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B1_valid;
	wire Tile_X01_Y04_SB_T1_WEST_SB_IN_B17_ready;
	wire Tile_X01_Y04_SB_T1_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y04_SB_T1_WEST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y04_SB_T1_WEST_SB_OUT_B17;
	wire Tile_X01_Y04_SB_T1_WEST_SB_OUT_B17_valid;
	wire Tile_X01_Y04_SB_T1_WEST_SB_OUT_B1_valid;
	wire Tile_X01_Y04_SB_T2_EAST_SB_IN_B17_ready;
	wire Tile_X01_Y04_SB_T2_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y04_SB_T2_EAST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y04_SB_T2_EAST_SB_OUT_B17;
	wire Tile_X01_Y04_SB_T2_EAST_SB_OUT_B17_valid;
	wire Tile_X01_Y04_SB_T2_EAST_SB_OUT_B1_valid;
	wire Tile_X01_Y04_SB_T2_NORTH_SB_IN_B17_ready;
	wire Tile_X01_Y04_SB_T2_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B17;
	wire Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B17_valid;
	wire Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B1_valid;
	wire Tile_X01_Y04_SB_T2_SOUTH_SB_IN_B17_ready;
	wire Tile_X01_Y04_SB_T2_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B17;
	wire Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B17_valid;
	wire Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B1_valid;
	wire Tile_X01_Y04_SB_T2_WEST_SB_IN_B17_ready;
	wire Tile_X01_Y04_SB_T2_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y04_SB_T2_WEST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y04_SB_T2_WEST_SB_OUT_B17;
	wire Tile_X01_Y04_SB_T2_WEST_SB_OUT_B17_valid;
	wire Tile_X01_Y04_SB_T2_WEST_SB_OUT_B1_valid;
	wire Tile_X01_Y04_SB_T3_EAST_SB_IN_B17_ready;
	wire Tile_X01_Y04_SB_T3_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y04_SB_T3_EAST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y04_SB_T3_EAST_SB_OUT_B17;
	wire Tile_X01_Y04_SB_T3_EAST_SB_OUT_B17_valid;
	wire Tile_X01_Y04_SB_T3_EAST_SB_OUT_B1_valid;
	wire Tile_X01_Y04_SB_T3_NORTH_SB_IN_B17_ready;
	wire Tile_X01_Y04_SB_T3_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B17;
	wire Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B17_valid;
	wire Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B1_valid;
	wire Tile_X01_Y04_SB_T3_SOUTH_SB_IN_B17_ready;
	wire Tile_X01_Y04_SB_T3_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y04_SB_T3_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y04_SB_T3_SOUTH_SB_OUT_B17;
	wire Tile_X01_Y04_SB_T3_SOUTH_SB_OUT_B17_valid;
	wire Tile_X01_Y04_SB_T3_SOUTH_SB_OUT_B1_valid;
	wire Tile_X01_Y04_SB_T3_WEST_SB_IN_B17_ready;
	wire Tile_X01_Y04_SB_T3_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y04_SB_T3_WEST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y04_SB_T3_WEST_SB_OUT_B17;
	wire Tile_X01_Y04_SB_T3_WEST_SB_OUT_B17_valid;
	wire Tile_X01_Y04_SB_T3_WEST_SB_OUT_B1_valid;
	wire Tile_X01_Y04_SB_T4_EAST_SB_IN_B17_ready;
	wire Tile_X01_Y04_SB_T4_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y04_SB_T4_EAST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y04_SB_T4_EAST_SB_OUT_B17;
	wire Tile_X01_Y04_SB_T4_EAST_SB_OUT_B17_valid;
	wire Tile_X01_Y04_SB_T4_EAST_SB_OUT_B1_valid;
	wire Tile_X01_Y04_SB_T4_NORTH_SB_IN_B17_ready;
	wire Tile_X01_Y04_SB_T4_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B17;
	wire Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B17_valid;
	wire Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B1_valid;
	wire Tile_X01_Y04_SB_T4_SOUTH_SB_IN_B17_ready;
	wire Tile_X01_Y04_SB_T4_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y04_SB_T4_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X01_Y04_SB_T4_SOUTH_SB_OUT_B17;
	wire Tile_X01_Y04_SB_T4_SOUTH_SB_OUT_B17_valid;
	wire Tile_X01_Y04_SB_T4_SOUTH_SB_OUT_B1_valid;
	wire Tile_X01_Y04_SB_T4_WEST_SB_IN_B17_ready;
	wire Tile_X01_Y04_SB_T4_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X01_Y04_SB_T4_WEST_SB_OUT_B1;
	wire [16:0] Tile_X01_Y04_SB_T4_WEST_SB_OUT_B17;
	wire Tile_X01_Y04_SB_T4_WEST_SB_OUT_B17_valid;
	wire Tile_X01_Y04_SB_T4_WEST_SB_OUT_B1_valid;
	wire Tile_X01_Y04_clk_out;
	wire Tile_X01_Y04_clk_pass_through_out_bot;
	wire Tile_X01_Y04_clk_pass_through_out_right;
	wire [31:0] Tile_X01_Y04_config_out_config_addr;
	wire [31:0] Tile_X01_Y04_config_out_config_data;
	wire [0:0] Tile_X01_Y04_config_out_read;
	wire [0:0] Tile_X01_Y04_config_out_write;
	wire [0:0] Tile_X01_Y04_flush_out;
	wire [8:0] Tile_X01_Y04_hi;
	wire [7:0] Tile_X01_Y04_lo;
	wire [31:0] Tile_X01_Y04_read_config_data;
	wire Tile_X01_Y04_reset_out;
	wire [0:0] Tile_X01_Y04_stall_out;
	wire Tile_X02_Y00_clk_out;
	wire [31:0] Tile_X02_Y00_config_out_config_addr;
	wire [31:0] Tile_X02_Y00_config_out_config_data;
	wire [0:0] Tile_X02_Y00_config_out_read;
	wire [0:0] Tile_X02_Y00_config_out_write;
	wire Tile_X02_Y00_f2io_17_ready;
	wire Tile_X02_Y00_f2io_1_ready;
	wire [0:0] Tile_X02_Y00_flush_out;
	wire Tile_X02_Y00_glb2io_17_ready;
	wire Tile_X02_Y00_glb2io_1_ready;
	wire [8:0] Tile_X02_Y00_hi;
	wire [0:0] Tile_X02_Y00_io2f_1;
	wire [16:0] Tile_X02_Y00_io2f_17;
	wire Tile_X02_Y00_io2f_17_valid;
	wire Tile_X02_Y00_io2f_1_valid;
	wire [0:0] Tile_X02_Y00_io2glb_1;
	wire [16:0] Tile_X02_Y00_io2glb_17;
	wire Tile_X02_Y00_io2glb_17_valid;
	wire Tile_X02_Y00_io2glb_1_valid;
	wire [7:0] Tile_X02_Y00_lo;
	wire [31:0] Tile_X02_Y00_read_config_data;
	wire Tile_X02_Y00_reset_out;
	wire [0:0] Tile_X02_Y00_stall_out;
	wire Tile_X02_Y01_SB_T0_EAST_SB_IN_B17_ready;
	wire Tile_X02_Y01_SB_T0_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y01_SB_T0_EAST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y01_SB_T0_EAST_SB_OUT_B17;
	wire Tile_X02_Y01_SB_T0_EAST_SB_OUT_B17_valid;
	wire Tile_X02_Y01_SB_T0_EAST_SB_OUT_B1_valid;
	wire Tile_X02_Y01_SB_T0_NORTH_SB_IN_B17_ready;
	wire Tile_X02_Y01_SB_T0_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B17;
	wire Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B17_valid;
	wire Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B1_valid;
	wire Tile_X02_Y01_SB_T0_SOUTH_SB_IN_B17_ready;
	wire Tile_X02_Y01_SB_T0_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B17;
	wire Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B17_valid;
	wire Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B1_valid;
	wire Tile_X02_Y01_SB_T0_WEST_SB_IN_B17_ready;
	wire Tile_X02_Y01_SB_T0_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y01_SB_T0_WEST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y01_SB_T0_WEST_SB_OUT_B17;
	wire Tile_X02_Y01_SB_T0_WEST_SB_OUT_B17_valid;
	wire Tile_X02_Y01_SB_T0_WEST_SB_OUT_B1_valid;
	wire Tile_X02_Y01_SB_T1_EAST_SB_IN_B17_ready;
	wire Tile_X02_Y01_SB_T1_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y01_SB_T1_EAST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y01_SB_T1_EAST_SB_OUT_B17;
	wire Tile_X02_Y01_SB_T1_EAST_SB_OUT_B17_valid;
	wire Tile_X02_Y01_SB_T1_EAST_SB_OUT_B1_valid;
	wire Tile_X02_Y01_SB_T1_NORTH_SB_IN_B17_ready;
	wire Tile_X02_Y01_SB_T1_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y01_SB_T1_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y01_SB_T1_NORTH_SB_OUT_B17;
	wire Tile_X02_Y01_SB_T1_NORTH_SB_OUT_B17_valid;
	wire Tile_X02_Y01_SB_T1_NORTH_SB_OUT_B1_valid;
	wire Tile_X02_Y01_SB_T1_SOUTH_SB_IN_B17_ready;
	wire Tile_X02_Y01_SB_T1_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B17;
	wire Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B17_valid;
	wire Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B1_valid;
	wire Tile_X02_Y01_SB_T1_WEST_SB_IN_B17_ready;
	wire Tile_X02_Y01_SB_T1_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y01_SB_T1_WEST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y01_SB_T1_WEST_SB_OUT_B17;
	wire Tile_X02_Y01_SB_T1_WEST_SB_OUT_B17_valid;
	wire Tile_X02_Y01_SB_T1_WEST_SB_OUT_B1_valid;
	wire Tile_X02_Y01_SB_T2_EAST_SB_IN_B17_ready;
	wire Tile_X02_Y01_SB_T2_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y01_SB_T2_EAST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y01_SB_T2_EAST_SB_OUT_B17;
	wire Tile_X02_Y01_SB_T2_EAST_SB_OUT_B17_valid;
	wire Tile_X02_Y01_SB_T2_EAST_SB_OUT_B1_valid;
	wire Tile_X02_Y01_SB_T2_NORTH_SB_IN_B17_ready;
	wire Tile_X02_Y01_SB_T2_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y01_SB_T2_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y01_SB_T2_NORTH_SB_OUT_B17;
	wire Tile_X02_Y01_SB_T2_NORTH_SB_OUT_B17_valid;
	wire Tile_X02_Y01_SB_T2_NORTH_SB_OUT_B1_valid;
	wire Tile_X02_Y01_SB_T2_SOUTH_SB_IN_B17_ready;
	wire Tile_X02_Y01_SB_T2_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B17;
	wire Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B17_valid;
	wire Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B1_valid;
	wire Tile_X02_Y01_SB_T2_WEST_SB_IN_B17_ready;
	wire Tile_X02_Y01_SB_T2_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y01_SB_T2_WEST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y01_SB_T2_WEST_SB_OUT_B17;
	wire Tile_X02_Y01_SB_T2_WEST_SB_OUT_B17_valid;
	wire Tile_X02_Y01_SB_T2_WEST_SB_OUT_B1_valid;
	wire Tile_X02_Y01_SB_T3_EAST_SB_IN_B17_ready;
	wire Tile_X02_Y01_SB_T3_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y01_SB_T3_EAST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y01_SB_T3_EAST_SB_OUT_B17;
	wire Tile_X02_Y01_SB_T3_EAST_SB_OUT_B17_valid;
	wire Tile_X02_Y01_SB_T3_EAST_SB_OUT_B1_valid;
	wire Tile_X02_Y01_SB_T3_NORTH_SB_IN_B17_ready;
	wire Tile_X02_Y01_SB_T3_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y01_SB_T3_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y01_SB_T3_NORTH_SB_OUT_B17;
	wire Tile_X02_Y01_SB_T3_NORTH_SB_OUT_B17_valid;
	wire Tile_X02_Y01_SB_T3_NORTH_SB_OUT_B1_valid;
	wire Tile_X02_Y01_SB_T3_SOUTH_SB_IN_B17_ready;
	wire Tile_X02_Y01_SB_T3_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B17;
	wire Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B17_valid;
	wire Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B1_valid;
	wire Tile_X02_Y01_SB_T3_WEST_SB_IN_B17_ready;
	wire Tile_X02_Y01_SB_T3_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y01_SB_T3_WEST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y01_SB_T3_WEST_SB_OUT_B17;
	wire Tile_X02_Y01_SB_T3_WEST_SB_OUT_B17_valid;
	wire Tile_X02_Y01_SB_T3_WEST_SB_OUT_B1_valid;
	wire Tile_X02_Y01_SB_T4_EAST_SB_IN_B17_ready;
	wire Tile_X02_Y01_SB_T4_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y01_SB_T4_EAST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y01_SB_T4_EAST_SB_OUT_B17;
	wire Tile_X02_Y01_SB_T4_EAST_SB_OUT_B17_valid;
	wire Tile_X02_Y01_SB_T4_EAST_SB_OUT_B1_valid;
	wire Tile_X02_Y01_SB_T4_NORTH_SB_IN_B17_ready;
	wire Tile_X02_Y01_SB_T4_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y01_SB_T4_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y01_SB_T4_NORTH_SB_OUT_B17;
	wire Tile_X02_Y01_SB_T4_NORTH_SB_OUT_B17_valid;
	wire Tile_X02_Y01_SB_T4_NORTH_SB_OUT_B1_valid;
	wire Tile_X02_Y01_SB_T4_SOUTH_SB_IN_B17_ready;
	wire Tile_X02_Y01_SB_T4_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B17;
	wire Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B17_valid;
	wire Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B1_valid;
	wire Tile_X02_Y01_SB_T4_WEST_SB_IN_B17_ready;
	wire Tile_X02_Y01_SB_T4_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y01_SB_T4_WEST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y01_SB_T4_WEST_SB_OUT_B17;
	wire Tile_X02_Y01_SB_T4_WEST_SB_OUT_B17_valid;
	wire Tile_X02_Y01_SB_T4_WEST_SB_OUT_B1_valid;
	wire Tile_X02_Y01_clk_out;
	wire Tile_X02_Y01_clk_pass_through_out_bot;
	wire Tile_X02_Y01_clk_pass_through_out_right;
	wire [31:0] Tile_X02_Y01_config_out_config_addr;
	wire [31:0] Tile_X02_Y01_config_out_config_data;
	wire [0:0] Tile_X02_Y01_config_out_read;
	wire [0:0] Tile_X02_Y01_config_out_write;
	wire [0:0] Tile_X02_Y01_flush_out;
	wire [8:0] Tile_X02_Y01_hi;
	wire [7:0] Tile_X02_Y01_lo;
	wire [31:0] Tile_X02_Y01_read_config_data;
	wire Tile_X02_Y01_reset_out;
	wire [0:0] Tile_X02_Y01_stall_out;
	wire Tile_X02_Y02_SB_T0_EAST_SB_IN_B17_ready;
	wire Tile_X02_Y02_SB_T0_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y02_SB_T0_EAST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y02_SB_T0_EAST_SB_OUT_B17;
	wire Tile_X02_Y02_SB_T0_EAST_SB_OUT_B17_valid;
	wire Tile_X02_Y02_SB_T0_EAST_SB_OUT_B1_valid;
	wire Tile_X02_Y02_SB_T0_NORTH_SB_IN_B17_ready;
	wire Tile_X02_Y02_SB_T0_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B17;
	wire Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B17_valid;
	wire Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B1_valid;
	wire Tile_X02_Y02_SB_T0_SOUTH_SB_IN_B17_ready;
	wire Tile_X02_Y02_SB_T0_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B17;
	wire Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B17_valid;
	wire Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B1_valid;
	wire Tile_X02_Y02_SB_T0_WEST_SB_IN_B17_ready;
	wire Tile_X02_Y02_SB_T0_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y02_SB_T0_WEST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y02_SB_T0_WEST_SB_OUT_B17;
	wire Tile_X02_Y02_SB_T0_WEST_SB_OUT_B17_valid;
	wire Tile_X02_Y02_SB_T0_WEST_SB_OUT_B1_valid;
	wire Tile_X02_Y02_SB_T1_EAST_SB_IN_B17_ready;
	wire Tile_X02_Y02_SB_T1_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y02_SB_T1_EAST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y02_SB_T1_EAST_SB_OUT_B17;
	wire Tile_X02_Y02_SB_T1_EAST_SB_OUT_B17_valid;
	wire Tile_X02_Y02_SB_T1_EAST_SB_OUT_B1_valid;
	wire Tile_X02_Y02_SB_T1_NORTH_SB_IN_B17_ready;
	wire Tile_X02_Y02_SB_T1_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B17;
	wire Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B17_valid;
	wire Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B1_valid;
	wire Tile_X02_Y02_SB_T1_SOUTH_SB_IN_B17_ready;
	wire Tile_X02_Y02_SB_T1_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B17;
	wire Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B17_valid;
	wire Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B1_valid;
	wire Tile_X02_Y02_SB_T1_WEST_SB_IN_B17_ready;
	wire Tile_X02_Y02_SB_T1_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y02_SB_T1_WEST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y02_SB_T1_WEST_SB_OUT_B17;
	wire Tile_X02_Y02_SB_T1_WEST_SB_OUT_B17_valid;
	wire Tile_X02_Y02_SB_T1_WEST_SB_OUT_B1_valid;
	wire Tile_X02_Y02_SB_T2_EAST_SB_IN_B17_ready;
	wire Tile_X02_Y02_SB_T2_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y02_SB_T2_EAST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y02_SB_T2_EAST_SB_OUT_B17;
	wire Tile_X02_Y02_SB_T2_EAST_SB_OUT_B17_valid;
	wire Tile_X02_Y02_SB_T2_EAST_SB_OUT_B1_valid;
	wire Tile_X02_Y02_SB_T2_NORTH_SB_IN_B17_ready;
	wire Tile_X02_Y02_SB_T2_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B17;
	wire Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B17_valid;
	wire Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B1_valid;
	wire Tile_X02_Y02_SB_T2_SOUTH_SB_IN_B17_ready;
	wire Tile_X02_Y02_SB_T2_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B17;
	wire Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B17_valid;
	wire Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B1_valid;
	wire Tile_X02_Y02_SB_T2_WEST_SB_IN_B17_ready;
	wire Tile_X02_Y02_SB_T2_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y02_SB_T2_WEST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y02_SB_T2_WEST_SB_OUT_B17;
	wire Tile_X02_Y02_SB_T2_WEST_SB_OUT_B17_valid;
	wire Tile_X02_Y02_SB_T2_WEST_SB_OUT_B1_valid;
	wire Tile_X02_Y02_SB_T3_EAST_SB_IN_B17_ready;
	wire Tile_X02_Y02_SB_T3_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y02_SB_T3_EAST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y02_SB_T3_EAST_SB_OUT_B17;
	wire Tile_X02_Y02_SB_T3_EAST_SB_OUT_B17_valid;
	wire Tile_X02_Y02_SB_T3_EAST_SB_OUT_B1_valid;
	wire Tile_X02_Y02_SB_T3_NORTH_SB_IN_B17_ready;
	wire Tile_X02_Y02_SB_T3_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B17;
	wire Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B17_valid;
	wire Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B1_valid;
	wire Tile_X02_Y02_SB_T3_SOUTH_SB_IN_B17_ready;
	wire Tile_X02_Y02_SB_T3_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B17;
	wire Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B17_valid;
	wire Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B1_valid;
	wire Tile_X02_Y02_SB_T3_WEST_SB_IN_B17_ready;
	wire Tile_X02_Y02_SB_T3_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y02_SB_T3_WEST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y02_SB_T3_WEST_SB_OUT_B17;
	wire Tile_X02_Y02_SB_T3_WEST_SB_OUT_B17_valid;
	wire Tile_X02_Y02_SB_T3_WEST_SB_OUT_B1_valid;
	wire Tile_X02_Y02_SB_T4_EAST_SB_IN_B17_ready;
	wire Tile_X02_Y02_SB_T4_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y02_SB_T4_EAST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y02_SB_T4_EAST_SB_OUT_B17;
	wire Tile_X02_Y02_SB_T4_EAST_SB_OUT_B17_valid;
	wire Tile_X02_Y02_SB_T4_EAST_SB_OUT_B1_valid;
	wire Tile_X02_Y02_SB_T4_NORTH_SB_IN_B17_ready;
	wire Tile_X02_Y02_SB_T4_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B17;
	wire Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B17_valid;
	wire Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B1_valid;
	wire Tile_X02_Y02_SB_T4_SOUTH_SB_IN_B17_ready;
	wire Tile_X02_Y02_SB_T4_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B17;
	wire Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B17_valid;
	wire Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B1_valid;
	wire Tile_X02_Y02_SB_T4_WEST_SB_IN_B17_ready;
	wire Tile_X02_Y02_SB_T4_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y02_SB_T4_WEST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y02_SB_T4_WEST_SB_OUT_B17;
	wire Tile_X02_Y02_SB_T4_WEST_SB_OUT_B17_valid;
	wire Tile_X02_Y02_SB_T4_WEST_SB_OUT_B1_valid;
	wire Tile_X02_Y02_clk_out;
	wire Tile_X02_Y02_clk_pass_through_out_bot;
	wire Tile_X02_Y02_clk_pass_through_out_right;
	wire [31:0] Tile_X02_Y02_config_out_config_addr;
	wire [31:0] Tile_X02_Y02_config_out_config_data;
	wire [0:0] Tile_X02_Y02_config_out_read;
	wire [0:0] Tile_X02_Y02_config_out_write;
	wire [0:0] Tile_X02_Y02_flush_out;
	wire [8:0] Tile_X02_Y02_hi;
	wire [7:0] Tile_X02_Y02_lo;
	wire [31:0] Tile_X02_Y02_read_config_data;
	wire Tile_X02_Y02_reset_out;
	wire [0:0] Tile_X02_Y02_stall_out;
	wire Tile_X02_Y03_SB_T0_EAST_SB_IN_B17_ready;
	wire Tile_X02_Y03_SB_T0_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y03_SB_T0_EAST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y03_SB_T0_EAST_SB_OUT_B17;
	wire Tile_X02_Y03_SB_T0_EAST_SB_OUT_B17_valid;
	wire Tile_X02_Y03_SB_T0_EAST_SB_OUT_B1_valid;
	wire Tile_X02_Y03_SB_T0_NORTH_SB_IN_B17_ready;
	wire Tile_X02_Y03_SB_T0_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B17;
	wire Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B17_valid;
	wire Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B1_valid;
	wire Tile_X02_Y03_SB_T0_SOUTH_SB_IN_B17_ready;
	wire Tile_X02_Y03_SB_T0_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B17;
	wire Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B17_valid;
	wire Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B1_valid;
	wire Tile_X02_Y03_SB_T0_WEST_SB_IN_B17_ready;
	wire Tile_X02_Y03_SB_T0_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y03_SB_T0_WEST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y03_SB_T0_WEST_SB_OUT_B17;
	wire Tile_X02_Y03_SB_T0_WEST_SB_OUT_B17_valid;
	wire Tile_X02_Y03_SB_T0_WEST_SB_OUT_B1_valid;
	wire Tile_X02_Y03_SB_T1_EAST_SB_IN_B17_ready;
	wire Tile_X02_Y03_SB_T1_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y03_SB_T1_EAST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y03_SB_T1_EAST_SB_OUT_B17;
	wire Tile_X02_Y03_SB_T1_EAST_SB_OUT_B17_valid;
	wire Tile_X02_Y03_SB_T1_EAST_SB_OUT_B1_valid;
	wire Tile_X02_Y03_SB_T1_NORTH_SB_IN_B17_ready;
	wire Tile_X02_Y03_SB_T1_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B17;
	wire Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B17_valid;
	wire Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B1_valid;
	wire Tile_X02_Y03_SB_T1_SOUTH_SB_IN_B17_ready;
	wire Tile_X02_Y03_SB_T1_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B17;
	wire Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B17_valid;
	wire Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B1_valid;
	wire Tile_X02_Y03_SB_T1_WEST_SB_IN_B17_ready;
	wire Tile_X02_Y03_SB_T1_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y03_SB_T1_WEST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y03_SB_T1_WEST_SB_OUT_B17;
	wire Tile_X02_Y03_SB_T1_WEST_SB_OUT_B17_valid;
	wire Tile_X02_Y03_SB_T1_WEST_SB_OUT_B1_valid;
	wire Tile_X02_Y03_SB_T2_EAST_SB_IN_B17_ready;
	wire Tile_X02_Y03_SB_T2_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y03_SB_T2_EAST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y03_SB_T2_EAST_SB_OUT_B17;
	wire Tile_X02_Y03_SB_T2_EAST_SB_OUT_B17_valid;
	wire Tile_X02_Y03_SB_T2_EAST_SB_OUT_B1_valid;
	wire Tile_X02_Y03_SB_T2_NORTH_SB_IN_B17_ready;
	wire Tile_X02_Y03_SB_T2_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B17;
	wire Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B17_valid;
	wire Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B1_valid;
	wire Tile_X02_Y03_SB_T2_SOUTH_SB_IN_B17_ready;
	wire Tile_X02_Y03_SB_T2_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B17;
	wire Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B17_valid;
	wire Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B1_valid;
	wire Tile_X02_Y03_SB_T2_WEST_SB_IN_B17_ready;
	wire Tile_X02_Y03_SB_T2_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y03_SB_T2_WEST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y03_SB_T2_WEST_SB_OUT_B17;
	wire Tile_X02_Y03_SB_T2_WEST_SB_OUT_B17_valid;
	wire Tile_X02_Y03_SB_T2_WEST_SB_OUT_B1_valid;
	wire Tile_X02_Y03_SB_T3_EAST_SB_IN_B17_ready;
	wire Tile_X02_Y03_SB_T3_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y03_SB_T3_EAST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y03_SB_T3_EAST_SB_OUT_B17;
	wire Tile_X02_Y03_SB_T3_EAST_SB_OUT_B17_valid;
	wire Tile_X02_Y03_SB_T3_EAST_SB_OUT_B1_valid;
	wire Tile_X02_Y03_SB_T3_NORTH_SB_IN_B17_ready;
	wire Tile_X02_Y03_SB_T3_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B17;
	wire Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B17_valid;
	wire Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B1_valid;
	wire Tile_X02_Y03_SB_T3_SOUTH_SB_IN_B17_ready;
	wire Tile_X02_Y03_SB_T3_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B17;
	wire Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B17_valid;
	wire Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B1_valid;
	wire Tile_X02_Y03_SB_T3_WEST_SB_IN_B17_ready;
	wire Tile_X02_Y03_SB_T3_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y03_SB_T3_WEST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y03_SB_T3_WEST_SB_OUT_B17;
	wire Tile_X02_Y03_SB_T3_WEST_SB_OUT_B17_valid;
	wire Tile_X02_Y03_SB_T3_WEST_SB_OUT_B1_valid;
	wire Tile_X02_Y03_SB_T4_EAST_SB_IN_B17_ready;
	wire Tile_X02_Y03_SB_T4_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y03_SB_T4_EAST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y03_SB_T4_EAST_SB_OUT_B17;
	wire Tile_X02_Y03_SB_T4_EAST_SB_OUT_B17_valid;
	wire Tile_X02_Y03_SB_T4_EAST_SB_OUT_B1_valid;
	wire Tile_X02_Y03_SB_T4_NORTH_SB_IN_B17_ready;
	wire Tile_X02_Y03_SB_T4_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B17;
	wire Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B17_valid;
	wire Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B1_valid;
	wire Tile_X02_Y03_SB_T4_SOUTH_SB_IN_B17_ready;
	wire Tile_X02_Y03_SB_T4_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B17;
	wire Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B17_valid;
	wire Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B1_valid;
	wire Tile_X02_Y03_SB_T4_WEST_SB_IN_B17_ready;
	wire Tile_X02_Y03_SB_T4_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y03_SB_T4_WEST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y03_SB_T4_WEST_SB_OUT_B17;
	wire Tile_X02_Y03_SB_T4_WEST_SB_OUT_B17_valid;
	wire Tile_X02_Y03_SB_T4_WEST_SB_OUT_B1_valid;
	wire Tile_X02_Y03_clk_out;
	wire Tile_X02_Y03_clk_pass_through_out_bot;
	wire Tile_X02_Y03_clk_pass_through_out_right;
	wire [31:0] Tile_X02_Y03_config_out_config_addr;
	wire [31:0] Tile_X02_Y03_config_out_config_data;
	wire [0:0] Tile_X02_Y03_config_out_read;
	wire [0:0] Tile_X02_Y03_config_out_write;
	wire [0:0] Tile_X02_Y03_flush_out;
	wire [8:0] Tile_X02_Y03_hi;
	wire [7:0] Tile_X02_Y03_lo;
	wire [31:0] Tile_X02_Y03_read_config_data;
	wire Tile_X02_Y03_reset_out;
	wire [0:0] Tile_X02_Y03_stall_out;
	wire Tile_X02_Y04_SB_T0_EAST_SB_IN_B17_ready;
	wire Tile_X02_Y04_SB_T0_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y04_SB_T0_EAST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y04_SB_T0_EAST_SB_OUT_B17;
	wire Tile_X02_Y04_SB_T0_EAST_SB_OUT_B17_valid;
	wire Tile_X02_Y04_SB_T0_EAST_SB_OUT_B1_valid;
	wire Tile_X02_Y04_SB_T0_NORTH_SB_IN_B17_ready;
	wire Tile_X02_Y04_SB_T0_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B17;
	wire Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B17_valid;
	wire Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B1_valid;
	wire Tile_X02_Y04_SB_T0_SOUTH_SB_IN_B17_ready;
	wire Tile_X02_Y04_SB_T0_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B17;
	wire Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B17_valid;
	wire Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B1_valid;
	wire Tile_X02_Y04_SB_T0_WEST_SB_IN_B17_ready;
	wire Tile_X02_Y04_SB_T0_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y04_SB_T0_WEST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y04_SB_T0_WEST_SB_OUT_B17;
	wire Tile_X02_Y04_SB_T0_WEST_SB_OUT_B17_valid;
	wire Tile_X02_Y04_SB_T0_WEST_SB_OUT_B1_valid;
	wire Tile_X02_Y04_SB_T1_EAST_SB_IN_B17_ready;
	wire Tile_X02_Y04_SB_T1_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y04_SB_T1_EAST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y04_SB_T1_EAST_SB_OUT_B17;
	wire Tile_X02_Y04_SB_T1_EAST_SB_OUT_B17_valid;
	wire Tile_X02_Y04_SB_T1_EAST_SB_OUT_B1_valid;
	wire Tile_X02_Y04_SB_T1_NORTH_SB_IN_B17_ready;
	wire Tile_X02_Y04_SB_T1_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B17;
	wire Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B17_valid;
	wire Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B1_valid;
	wire Tile_X02_Y04_SB_T1_SOUTH_SB_IN_B17_ready;
	wire Tile_X02_Y04_SB_T1_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B17;
	wire Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B17_valid;
	wire Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B1_valid;
	wire Tile_X02_Y04_SB_T1_WEST_SB_IN_B17_ready;
	wire Tile_X02_Y04_SB_T1_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y04_SB_T1_WEST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y04_SB_T1_WEST_SB_OUT_B17;
	wire Tile_X02_Y04_SB_T1_WEST_SB_OUT_B17_valid;
	wire Tile_X02_Y04_SB_T1_WEST_SB_OUT_B1_valid;
	wire Tile_X02_Y04_SB_T2_EAST_SB_IN_B17_ready;
	wire Tile_X02_Y04_SB_T2_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y04_SB_T2_EAST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y04_SB_T2_EAST_SB_OUT_B17;
	wire Tile_X02_Y04_SB_T2_EAST_SB_OUT_B17_valid;
	wire Tile_X02_Y04_SB_T2_EAST_SB_OUT_B1_valid;
	wire Tile_X02_Y04_SB_T2_NORTH_SB_IN_B17_ready;
	wire Tile_X02_Y04_SB_T2_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B17;
	wire Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B17_valid;
	wire Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B1_valid;
	wire Tile_X02_Y04_SB_T2_SOUTH_SB_IN_B17_ready;
	wire Tile_X02_Y04_SB_T2_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B17;
	wire Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B17_valid;
	wire Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B1_valid;
	wire Tile_X02_Y04_SB_T2_WEST_SB_IN_B17_ready;
	wire Tile_X02_Y04_SB_T2_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y04_SB_T2_WEST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y04_SB_T2_WEST_SB_OUT_B17;
	wire Tile_X02_Y04_SB_T2_WEST_SB_OUT_B17_valid;
	wire Tile_X02_Y04_SB_T2_WEST_SB_OUT_B1_valid;
	wire Tile_X02_Y04_SB_T3_EAST_SB_IN_B17_ready;
	wire Tile_X02_Y04_SB_T3_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y04_SB_T3_EAST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y04_SB_T3_EAST_SB_OUT_B17;
	wire Tile_X02_Y04_SB_T3_EAST_SB_OUT_B17_valid;
	wire Tile_X02_Y04_SB_T3_EAST_SB_OUT_B1_valid;
	wire Tile_X02_Y04_SB_T3_NORTH_SB_IN_B17_ready;
	wire Tile_X02_Y04_SB_T3_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B17;
	wire Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B17_valid;
	wire Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B1_valid;
	wire Tile_X02_Y04_SB_T3_SOUTH_SB_IN_B17_ready;
	wire Tile_X02_Y04_SB_T3_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y04_SB_T3_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y04_SB_T3_SOUTH_SB_OUT_B17;
	wire Tile_X02_Y04_SB_T3_SOUTH_SB_OUT_B17_valid;
	wire Tile_X02_Y04_SB_T3_SOUTH_SB_OUT_B1_valid;
	wire Tile_X02_Y04_SB_T3_WEST_SB_IN_B17_ready;
	wire Tile_X02_Y04_SB_T3_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y04_SB_T3_WEST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y04_SB_T3_WEST_SB_OUT_B17;
	wire Tile_X02_Y04_SB_T3_WEST_SB_OUT_B17_valid;
	wire Tile_X02_Y04_SB_T3_WEST_SB_OUT_B1_valid;
	wire Tile_X02_Y04_SB_T4_EAST_SB_IN_B17_ready;
	wire Tile_X02_Y04_SB_T4_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y04_SB_T4_EAST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y04_SB_T4_EAST_SB_OUT_B17;
	wire Tile_X02_Y04_SB_T4_EAST_SB_OUT_B17_valid;
	wire Tile_X02_Y04_SB_T4_EAST_SB_OUT_B1_valid;
	wire Tile_X02_Y04_SB_T4_NORTH_SB_IN_B17_ready;
	wire Tile_X02_Y04_SB_T4_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B17;
	wire Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B17_valid;
	wire Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B1_valid;
	wire Tile_X02_Y04_SB_T4_SOUTH_SB_IN_B17_ready;
	wire Tile_X02_Y04_SB_T4_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y04_SB_T4_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X02_Y04_SB_T4_SOUTH_SB_OUT_B17;
	wire Tile_X02_Y04_SB_T4_SOUTH_SB_OUT_B17_valid;
	wire Tile_X02_Y04_SB_T4_SOUTH_SB_OUT_B1_valid;
	wire Tile_X02_Y04_SB_T4_WEST_SB_IN_B17_ready;
	wire Tile_X02_Y04_SB_T4_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X02_Y04_SB_T4_WEST_SB_OUT_B1;
	wire [16:0] Tile_X02_Y04_SB_T4_WEST_SB_OUT_B17;
	wire Tile_X02_Y04_SB_T4_WEST_SB_OUT_B17_valid;
	wire Tile_X02_Y04_SB_T4_WEST_SB_OUT_B1_valid;
	wire Tile_X02_Y04_clk_out;
	wire Tile_X02_Y04_clk_pass_through_out_bot;
	wire Tile_X02_Y04_clk_pass_through_out_right;
	wire [31:0] Tile_X02_Y04_config_out_config_addr;
	wire [31:0] Tile_X02_Y04_config_out_config_data;
	wire [0:0] Tile_X02_Y04_config_out_read;
	wire [0:0] Tile_X02_Y04_config_out_write;
	wire [0:0] Tile_X02_Y04_flush_out;
	wire [8:0] Tile_X02_Y04_hi;
	wire [7:0] Tile_X02_Y04_lo;
	wire [31:0] Tile_X02_Y04_read_config_data;
	wire Tile_X02_Y04_reset_out;
	wire [0:0] Tile_X02_Y04_stall_out;
	wire Tile_X03_Y00_clk_out;
	wire [31:0] Tile_X03_Y00_config_out_config_addr;
	wire [31:0] Tile_X03_Y00_config_out_config_data;
	wire [0:0] Tile_X03_Y00_config_out_read;
	wire [0:0] Tile_X03_Y00_config_out_write;
	wire Tile_X03_Y00_f2io_17_ready;
	wire Tile_X03_Y00_f2io_1_ready;
	wire [0:0] Tile_X03_Y00_flush_out;
	wire Tile_X03_Y00_glb2io_17_ready;
	wire Tile_X03_Y00_glb2io_1_ready;
	wire [8:0] Tile_X03_Y00_hi;
	wire [0:0] Tile_X03_Y00_io2f_1;
	wire [16:0] Tile_X03_Y00_io2f_17;
	wire Tile_X03_Y00_io2f_17_valid;
	wire Tile_X03_Y00_io2f_1_valid;
	wire [0:0] Tile_X03_Y00_io2glb_1;
	wire [16:0] Tile_X03_Y00_io2glb_17;
	wire Tile_X03_Y00_io2glb_17_valid;
	wire Tile_X03_Y00_io2glb_1_valid;
	wire [7:0] Tile_X03_Y00_lo;
	wire [31:0] Tile_X03_Y00_read_config_data;
	wire Tile_X03_Y00_reset_out;
	wire [0:0] Tile_X03_Y00_stall_out;
	wire Tile_X03_Y01_SB_T0_EAST_SB_IN_B17_ready;
	wire Tile_X03_Y01_SB_T0_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y01_SB_T0_EAST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y01_SB_T0_EAST_SB_OUT_B17;
	wire Tile_X03_Y01_SB_T0_EAST_SB_OUT_B17_valid;
	wire Tile_X03_Y01_SB_T0_EAST_SB_OUT_B1_valid;
	wire Tile_X03_Y01_SB_T0_NORTH_SB_IN_B17_ready;
	wire Tile_X03_Y01_SB_T0_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B17;
	wire Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B17_valid;
	wire Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B1_valid;
	wire Tile_X03_Y01_SB_T0_SOUTH_SB_IN_B17_ready;
	wire Tile_X03_Y01_SB_T0_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B17;
	wire Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B17_valid;
	wire Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B1_valid;
	wire Tile_X03_Y01_SB_T0_WEST_SB_IN_B17_ready;
	wire Tile_X03_Y01_SB_T0_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y01_SB_T0_WEST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y01_SB_T0_WEST_SB_OUT_B17;
	wire Tile_X03_Y01_SB_T0_WEST_SB_OUT_B17_valid;
	wire Tile_X03_Y01_SB_T0_WEST_SB_OUT_B1_valid;
	wire Tile_X03_Y01_SB_T1_EAST_SB_IN_B17_ready;
	wire Tile_X03_Y01_SB_T1_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y01_SB_T1_EAST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y01_SB_T1_EAST_SB_OUT_B17;
	wire Tile_X03_Y01_SB_T1_EAST_SB_OUT_B17_valid;
	wire Tile_X03_Y01_SB_T1_EAST_SB_OUT_B1_valid;
	wire Tile_X03_Y01_SB_T1_NORTH_SB_IN_B17_ready;
	wire Tile_X03_Y01_SB_T1_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y01_SB_T1_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y01_SB_T1_NORTH_SB_OUT_B17;
	wire Tile_X03_Y01_SB_T1_NORTH_SB_OUT_B17_valid;
	wire Tile_X03_Y01_SB_T1_NORTH_SB_OUT_B1_valid;
	wire Tile_X03_Y01_SB_T1_SOUTH_SB_IN_B17_ready;
	wire Tile_X03_Y01_SB_T1_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B17;
	wire Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B17_valid;
	wire Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B1_valid;
	wire Tile_X03_Y01_SB_T1_WEST_SB_IN_B17_ready;
	wire Tile_X03_Y01_SB_T1_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y01_SB_T1_WEST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y01_SB_T1_WEST_SB_OUT_B17;
	wire Tile_X03_Y01_SB_T1_WEST_SB_OUT_B17_valid;
	wire Tile_X03_Y01_SB_T1_WEST_SB_OUT_B1_valid;
	wire Tile_X03_Y01_SB_T2_EAST_SB_IN_B17_ready;
	wire Tile_X03_Y01_SB_T2_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y01_SB_T2_EAST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y01_SB_T2_EAST_SB_OUT_B17;
	wire Tile_X03_Y01_SB_T2_EAST_SB_OUT_B17_valid;
	wire Tile_X03_Y01_SB_T2_EAST_SB_OUT_B1_valid;
	wire Tile_X03_Y01_SB_T2_NORTH_SB_IN_B17_ready;
	wire Tile_X03_Y01_SB_T2_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y01_SB_T2_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y01_SB_T2_NORTH_SB_OUT_B17;
	wire Tile_X03_Y01_SB_T2_NORTH_SB_OUT_B17_valid;
	wire Tile_X03_Y01_SB_T2_NORTH_SB_OUT_B1_valid;
	wire Tile_X03_Y01_SB_T2_SOUTH_SB_IN_B17_ready;
	wire Tile_X03_Y01_SB_T2_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B17;
	wire Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B17_valid;
	wire Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B1_valid;
	wire Tile_X03_Y01_SB_T2_WEST_SB_IN_B17_ready;
	wire Tile_X03_Y01_SB_T2_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y01_SB_T2_WEST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y01_SB_T2_WEST_SB_OUT_B17;
	wire Tile_X03_Y01_SB_T2_WEST_SB_OUT_B17_valid;
	wire Tile_X03_Y01_SB_T2_WEST_SB_OUT_B1_valid;
	wire Tile_X03_Y01_SB_T3_EAST_SB_IN_B17_ready;
	wire Tile_X03_Y01_SB_T3_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y01_SB_T3_EAST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y01_SB_T3_EAST_SB_OUT_B17;
	wire Tile_X03_Y01_SB_T3_EAST_SB_OUT_B17_valid;
	wire Tile_X03_Y01_SB_T3_EAST_SB_OUT_B1_valid;
	wire Tile_X03_Y01_SB_T3_NORTH_SB_IN_B17_ready;
	wire Tile_X03_Y01_SB_T3_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y01_SB_T3_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y01_SB_T3_NORTH_SB_OUT_B17;
	wire Tile_X03_Y01_SB_T3_NORTH_SB_OUT_B17_valid;
	wire Tile_X03_Y01_SB_T3_NORTH_SB_OUT_B1_valid;
	wire Tile_X03_Y01_SB_T3_SOUTH_SB_IN_B17_ready;
	wire Tile_X03_Y01_SB_T3_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B17;
	wire Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B17_valid;
	wire Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B1_valid;
	wire Tile_X03_Y01_SB_T3_WEST_SB_IN_B17_ready;
	wire Tile_X03_Y01_SB_T3_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y01_SB_T3_WEST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y01_SB_T3_WEST_SB_OUT_B17;
	wire Tile_X03_Y01_SB_T3_WEST_SB_OUT_B17_valid;
	wire Tile_X03_Y01_SB_T3_WEST_SB_OUT_B1_valid;
	wire Tile_X03_Y01_SB_T4_EAST_SB_IN_B17_ready;
	wire Tile_X03_Y01_SB_T4_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y01_SB_T4_EAST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y01_SB_T4_EAST_SB_OUT_B17;
	wire Tile_X03_Y01_SB_T4_EAST_SB_OUT_B17_valid;
	wire Tile_X03_Y01_SB_T4_EAST_SB_OUT_B1_valid;
	wire Tile_X03_Y01_SB_T4_NORTH_SB_IN_B17_ready;
	wire Tile_X03_Y01_SB_T4_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y01_SB_T4_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y01_SB_T4_NORTH_SB_OUT_B17;
	wire Tile_X03_Y01_SB_T4_NORTH_SB_OUT_B17_valid;
	wire Tile_X03_Y01_SB_T4_NORTH_SB_OUT_B1_valid;
	wire Tile_X03_Y01_SB_T4_SOUTH_SB_IN_B17_ready;
	wire Tile_X03_Y01_SB_T4_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B17;
	wire Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B17_valid;
	wire Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B1_valid;
	wire Tile_X03_Y01_SB_T4_WEST_SB_IN_B17_ready;
	wire Tile_X03_Y01_SB_T4_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y01_SB_T4_WEST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y01_SB_T4_WEST_SB_OUT_B17;
	wire Tile_X03_Y01_SB_T4_WEST_SB_OUT_B17_valid;
	wire Tile_X03_Y01_SB_T4_WEST_SB_OUT_B1_valid;
	wire Tile_X03_Y01_clk_out;
	wire [31:0] Tile_X03_Y01_config_out_config_addr;
	wire [31:0] Tile_X03_Y01_config_out_config_data;
	wire [0:0] Tile_X03_Y01_config_out_read;
	wire [0:0] Tile_X03_Y01_config_out_write;
	wire [0:0] Tile_X03_Y01_flush_out;
	wire [8:0] Tile_X03_Y01_hi;
	wire [7:0] Tile_X03_Y01_lo;
	wire [31:0] Tile_X03_Y01_read_config_data;
	wire Tile_X03_Y01_reset_out;
	wire [0:0] Tile_X03_Y01_stall_out;
	wire Tile_X03_Y02_SB_T0_EAST_SB_IN_B17_ready;
	wire Tile_X03_Y02_SB_T0_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y02_SB_T0_EAST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y02_SB_T0_EAST_SB_OUT_B17;
	wire Tile_X03_Y02_SB_T0_EAST_SB_OUT_B17_valid;
	wire Tile_X03_Y02_SB_T0_EAST_SB_OUT_B1_valid;
	wire Tile_X03_Y02_SB_T0_NORTH_SB_IN_B17_ready;
	wire Tile_X03_Y02_SB_T0_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B17;
	wire Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B17_valid;
	wire Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B1_valid;
	wire Tile_X03_Y02_SB_T0_SOUTH_SB_IN_B17_ready;
	wire Tile_X03_Y02_SB_T0_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B17;
	wire Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B17_valid;
	wire Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B1_valid;
	wire Tile_X03_Y02_SB_T0_WEST_SB_IN_B17_ready;
	wire Tile_X03_Y02_SB_T0_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y02_SB_T0_WEST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y02_SB_T0_WEST_SB_OUT_B17;
	wire Tile_X03_Y02_SB_T0_WEST_SB_OUT_B17_valid;
	wire Tile_X03_Y02_SB_T0_WEST_SB_OUT_B1_valid;
	wire Tile_X03_Y02_SB_T1_EAST_SB_IN_B17_ready;
	wire Tile_X03_Y02_SB_T1_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y02_SB_T1_EAST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y02_SB_T1_EAST_SB_OUT_B17;
	wire Tile_X03_Y02_SB_T1_EAST_SB_OUT_B17_valid;
	wire Tile_X03_Y02_SB_T1_EAST_SB_OUT_B1_valid;
	wire Tile_X03_Y02_SB_T1_NORTH_SB_IN_B17_ready;
	wire Tile_X03_Y02_SB_T1_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B17;
	wire Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B17_valid;
	wire Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B1_valid;
	wire Tile_X03_Y02_SB_T1_SOUTH_SB_IN_B17_ready;
	wire Tile_X03_Y02_SB_T1_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B17;
	wire Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B17_valid;
	wire Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B1_valid;
	wire Tile_X03_Y02_SB_T1_WEST_SB_IN_B17_ready;
	wire Tile_X03_Y02_SB_T1_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y02_SB_T1_WEST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y02_SB_T1_WEST_SB_OUT_B17;
	wire Tile_X03_Y02_SB_T1_WEST_SB_OUT_B17_valid;
	wire Tile_X03_Y02_SB_T1_WEST_SB_OUT_B1_valid;
	wire Tile_X03_Y02_SB_T2_EAST_SB_IN_B17_ready;
	wire Tile_X03_Y02_SB_T2_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y02_SB_T2_EAST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y02_SB_T2_EAST_SB_OUT_B17;
	wire Tile_X03_Y02_SB_T2_EAST_SB_OUT_B17_valid;
	wire Tile_X03_Y02_SB_T2_EAST_SB_OUT_B1_valid;
	wire Tile_X03_Y02_SB_T2_NORTH_SB_IN_B17_ready;
	wire Tile_X03_Y02_SB_T2_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B17;
	wire Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B17_valid;
	wire Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B1_valid;
	wire Tile_X03_Y02_SB_T2_SOUTH_SB_IN_B17_ready;
	wire Tile_X03_Y02_SB_T2_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B17;
	wire Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B17_valid;
	wire Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B1_valid;
	wire Tile_X03_Y02_SB_T2_WEST_SB_IN_B17_ready;
	wire Tile_X03_Y02_SB_T2_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y02_SB_T2_WEST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y02_SB_T2_WEST_SB_OUT_B17;
	wire Tile_X03_Y02_SB_T2_WEST_SB_OUT_B17_valid;
	wire Tile_X03_Y02_SB_T2_WEST_SB_OUT_B1_valid;
	wire Tile_X03_Y02_SB_T3_EAST_SB_IN_B17_ready;
	wire Tile_X03_Y02_SB_T3_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y02_SB_T3_EAST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y02_SB_T3_EAST_SB_OUT_B17;
	wire Tile_X03_Y02_SB_T3_EAST_SB_OUT_B17_valid;
	wire Tile_X03_Y02_SB_T3_EAST_SB_OUT_B1_valid;
	wire Tile_X03_Y02_SB_T3_NORTH_SB_IN_B17_ready;
	wire Tile_X03_Y02_SB_T3_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B17;
	wire Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B17_valid;
	wire Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B1_valid;
	wire Tile_X03_Y02_SB_T3_SOUTH_SB_IN_B17_ready;
	wire Tile_X03_Y02_SB_T3_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B17;
	wire Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B17_valid;
	wire Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B1_valid;
	wire Tile_X03_Y02_SB_T3_WEST_SB_IN_B17_ready;
	wire Tile_X03_Y02_SB_T3_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y02_SB_T3_WEST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y02_SB_T3_WEST_SB_OUT_B17;
	wire Tile_X03_Y02_SB_T3_WEST_SB_OUT_B17_valid;
	wire Tile_X03_Y02_SB_T3_WEST_SB_OUT_B1_valid;
	wire Tile_X03_Y02_SB_T4_EAST_SB_IN_B17_ready;
	wire Tile_X03_Y02_SB_T4_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y02_SB_T4_EAST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y02_SB_T4_EAST_SB_OUT_B17;
	wire Tile_X03_Y02_SB_T4_EAST_SB_OUT_B17_valid;
	wire Tile_X03_Y02_SB_T4_EAST_SB_OUT_B1_valid;
	wire Tile_X03_Y02_SB_T4_NORTH_SB_IN_B17_ready;
	wire Tile_X03_Y02_SB_T4_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B17;
	wire Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B17_valid;
	wire Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B1_valid;
	wire Tile_X03_Y02_SB_T4_SOUTH_SB_IN_B17_ready;
	wire Tile_X03_Y02_SB_T4_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B17;
	wire Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B17_valid;
	wire Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B1_valid;
	wire Tile_X03_Y02_SB_T4_WEST_SB_IN_B17_ready;
	wire Tile_X03_Y02_SB_T4_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y02_SB_T4_WEST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y02_SB_T4_WEST_SB_OUT_B17;
	wire Tile_X03_Y02_SB_T4_WEST_SB_OUT_B17_valid;
	wire Tile_X03_Y02_SB_T4_WEST_SB_OUT_B1_valid;
	wire Tile_X03_Y02_clk_out;
	wire [31:0] Tile_X03_Y02_config_out_config_addr;
	wire [31:0] Tile_X03_Y02_config_out_config_data;
	wire [0:0] Tile_X03_Y02_config_out_read;
	wire [0:0] Tile_X03_Y02_config_out_write;
	wire [0:0] Tile_X03_Y02_flush_out;
	wire [8:0] Tile_X03_Y02_hi;
	wire [7:0] Tile_X03_Y02_lo;
	wire [31:0] Tile_X03_Y02_read_config_data;
	wire Tile_X03_Y02_reset_out;
	wire [0:0] Tile_X03_Y02_stall_out;
	wire Tile_X03_Y03_SB_T0_EAST_SB_IN_B17_ready;
	wire Tile_X03_Y03_SB_T0_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y03_SB_T0_EAST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y03_SB_T0_EAST_SB_OUT_B17;
	wire Tile_X03_Y03_SB_T0_EAST_SB_OUT_B17_valid;
	wire Tile_X03_Y03_SB_T0_EAST_SB_OUT_B1_valid;
	wire Tile_X03_Y03_SB_T0_NORTH_SB_IN_B17_ready;
	wire Tile_X03_Y03_SB_T0_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B17;
	wire Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B17_valid;
	wire Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B1_valid;
	wire Tile_X03_Y03_SB_T0_SOUTH_SB_IN_B17_ready;
	wire Tile_X03_Y03_SB_T0_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B17;
	wire Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B17_valid;
	wire Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B1_valid;
	wire Tile_X03_Y03_SB_T0_WEST_SB_IN_B17_ready;
	wire Tile_X03_Y03_SB_T0_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y03_SB_T0_WEST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y03_SB_T0_WEST_SB_OUT_B17;
	wire Tile_X03_Y03_SB_T0_WEST_SB_OUT_B17_valid;
	wire Tile_X03_Y03_SB_T0_WEST_SB_OUT_B1_valid;
	wire Tile_X03_Y03_SB_T1_EAST_SB_IN_B17_ready;
	wire Tile_X03_Y03_SB_T1_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y03_SB_T1_EAST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y03_SB_T1_EAST_SB_OUT_B17;
	wire Tile_X03_Y03_SB_T1_EAST_SB_OUT_B17_valid;
	wire Tile_X03_Y03_SB_T1_EAST_SB_OUT_B1_valid;
	wire Tile_X03_Y03_SB_T1_NORTH_SB_IN_B17_ready;
	wire Tile_X03_Y03_SB_T1_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B17;
	wire Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B17_valid;
	wire Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B1_valid;
	wire Tile_X03_Y03_SB_T1_SOUTH_SB_IN_B17_ready;
	wire Tile_X03_Y03_SB_T1_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B17;
	wire Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B17_valid;
	wire Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B1_valid;
	wire Tile_X03_Y03_SB_T1_WEST_SB_IN_B17_ready;
	wire Tile_X03_Y03_SB_T1_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y03_SB_T1_WEST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y03_SB_T1_WEST_SB_OUT_B17;
	wire Tile_X03_Y03_SB_T1_WEST_SB_OUT_B17_valid;
	wire Tile_X03_Y03_SB_T1_WEST_SB_OUT_B1_valid;
	wire Tile_X03_Y03_SB_T2_EAST_SB_IN_B17_ready;
	wire Tile_X03_Y03_SB_T2_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y03_SB_T2_EAST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y03_SB_T2_EAST_SB_OUT_B17;
	wire Tile_X03_Y03_SB_T2_EAST_SB_OUT_B17_valid;
	wire Tile_X03_Y03_SB_T2_EAST_SB_OUT_B1_valid;
	wire Tile_X03_Y03_SB_T2_NORTH_SB_IN_B17_ready;
	wire Tile_X03_Y03_SB_T2_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B17;
	wire Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B17_valid;
	wire Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B1_valid;
	wire Tile_X03_Y03_SB_T2_SOUTH_SB_IN_B17_ready;
	wire Tile_X03_Y03_SB_T2_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B17;
	wire Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B17_valid;
	wire Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B1_valid;
	wire Tile_X03_Y03_SB_T2_WEST_SB_IN_B17_ready;
	wire Tile_X03_Y03_SB_T2_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y03_SB_T2_WEST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y03_SB_T2_WEST_SB_OUT_B17;
	wire Tile_X03_Y03_SB_T2_WEST_SB_OUT_B17_valid;
	wire Tile_X03_Y03_SB_T2_WEST_SB_OUT_B1_valid;
	wire Tile_X03_Y03_SB_T3_EAST_SB_IN_B17_ready;
	wire Tile_X03_Y03_SB_T3_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y03_SB_T3_EAST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y03_SB_T3_EAST_SB_OUT_B17;
	wire Tile_X03_Y03_SB_T3_EAST_SB_OUT_B17_valid;
	wire Tile_X03_Y03_SB_T3_EAST_SB_OUT_B1_valid;
	wire Tile_X03_Y03_SB_T3_NORTH_SB_IN_B17_ready;
	wire Tile_X03_Y03_SB_T3_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B17;
	wire Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B17_valid;
	wire Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B1_valid;
	wire Tile_X03_Y03_SB_T3_SOUTH_SB_IN_B17_ready;
	wire Tile_X03_Y03_SB_T3_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B17;
	wire Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B17_valid;
	wire Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B1_valid;
	wire Tile_X03_Y03_SB_T3_WEST_SB_IN_B17_ready;
	wire Tile_X03_Y03_SB_T3_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y03_SB_T3_WEST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y03_SB_T3_WEST_SB_OUT_B17;
	wire Tile_X03_Y03_SB_T3_WEST_SB_OUT_B17_valid;
	wire Tile_X03_Y03_SB_T3_WEST_SB_OUT_B1_valid;
	wire Tile_X03_Y03_SB_T4_EAST_SB_IN_B17_ready;
	wire Tile_X03_Y03_SB_T4_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y03_SB_T4_EAST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y03_SB_T4_EAST_SB_OUT_B17;
	wire Tile_X03_Y03_SB_T4_EAST_SB_OUT_B17_valid;
	wire Tile_X03_Y03_SB_T4_EAST_SB_OUT_B1_valid;
	wire Tile_X03_Y03_SB_T4_NORTH_SB_IN_B17_ready;
	wire Tile_X03_Y03_SB_T4_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B17;
	wire Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B17_valid;
	wire Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B1_valid;
	wire Tile_X03_Y03_SB_T4_SOUTH_SB_IN_B17_ready;
	wire Tile_X03_Y03_SB_T4_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B17;
	wire Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B17_valid;
	wire Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B1_valid;
	wire Tile_X03_Y03_SB_T4_WEST_SB_IN_B17_ready;
	wire Tile_X03_Y03_SB_T4_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y03_SB_T4_WEST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y03_SB_T4_WEST_SB_OUT_B17;
	wire Tile_X03_Y03_SB_T4_WEST_SB_OUT_B17_valid;
	wire Tile_X03_Y03_SB_T4_WEST_SB_OUT_B1_valid;
	wire Tile_X03_Y03_clk_out;
	wire [31:0] Tile_X03_Y03_config_out_config_addr;
	wire [31:0] Tile_X03_Y03_config_out_config_data;
	wire [0:0] Tile_X03_Y03_config_out_read;
	wire [0:0] Tile_X03_Y03_config_out_write;
	wire [0:0] Tile_X03_Y03_flush_out;
	wire [8:0] Tile_X03_Y03_hi;
	wire [7:0] Tile_X03_Y03_lo;
	wire [31:0] Tile_X03_Y03_read_config_data;
	wire Tile_X03_Y03_reset_out;
	wire [0:0] Tile_X03_Y03_stall_out;
	wire Tile_X03_Y04_SB_T0_EAST_SB_IN_B17_ready;
	wire Tile_X03_Y04_SB_T0_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y04_SB_T0_EAST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y04_SB_T0_EAST_SB_OUT_B17;
	wire Tile_X03_Y04_SB_T0_EAST_SB_OUT_B17_valid;
	wire Tile_X03_Y04_SB_T0_EAST_SB_OUT_B1_valid;
	wire Tile_X03_Y04_SB_T0_NORTH_SB_IN_B17_ready;
	wire Tile_X03_Y04_SB_T0_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B17;
	wire Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B17_valid;
	wire Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B1_valid;
	wire Tile_X03_Y04_SB_T0_SOUTH_SB_IN_B17_ready;
	wire Tile_X03_Y04_SB_T0_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B17;
	wire Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B17_valid;
	wire Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B1_valid;
	wire Tile_X03_Y04_SB_T0_WEST_SB_IN_B17_ready;
	wire Tile_X03_Y04_SB_T0_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y04_SB_T0_WEST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y04_SB_T0_WEST_SB_OUT_B17;
	wire Tile_X03_Y04_SB_T0_WEST_SB_OUT_B17_valid;
	wire Tile_X03_Y04_SB_T0_WEST_SB_OUT_B1_valid;
	wire Tile_X03_Y04_SB_T1_EAST_SB_IN_B17_ready;
	wire Tile_X03_Y04_SB_T1_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y04_SB_T1_EAST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y04_SB_T1_EAST_SB_OUT_B17;
	wire Tile_X03_Y04_SB_T1_EAST_SB_OUT_B17_valid;
	wire Tile_X03_Y04_SB_T1_EAST_SB_OUT_B1_valid;
	wire Tile_X03_Y04_SB_T1_NORTH_SB_IN_B17_ready;
	wire Tile_X03_Y04_SB_T1_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B17;
	wire Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B17_valid;
	wire Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B1_valid;
	wire Tile_X03_Y04_SB_T1_SOUTH_SB_IN_B17_ready;
	wire Tile_X03_Y04_SB_T1_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B17;
	wire Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B17_valid;
	wire Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B1_valid;
	wire Tile_X03_Y04_SB_T1_WEST_SB_IN_B17_ready;
	wire Tile_X03_Y04_SB_T1_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y04_SB_T1_WEST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y04_SB_T1_WEST_SB_OUT_B17;
	wire Tile_X03_Y04_SB_T1_WEST_SB_OUT_B17_valid;
	wire Tile_X03_Y04_SB_T1_WEST_SB_OUT_B1_valid;
	wire Tile_X03_Y04_SB_T2_EAST_SB_IN_B17_ready;
	wire Tile_X03_Y04_SB_T2_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y04_SB_T2_EAST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y04_SB_T2_EAST_SB_OUT_B17;
	wire Tile_X03_Y04_SB_T2_EAST_SB_OUT_B17_valid;
	wire Tile_X03_Y04_SB_T2_EAST_SB_OUT_B1_valid;
	wire Tile_X03_Y04_SB_T2_NORTH_SB_IN_B17_ready;
	wire Tile_X03_Y04_SB_T2_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B17;
	wire Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B17_valid;
	wire Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B1_valid;
	wire Tile_X03_Y04_SB_T2_SOUTH_SB_IN_B17_ready;
	wire Tile_X03_Y04_SB_T2_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B17;
	wire Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B17_valid;
	wire Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B1_valid;
	wire Tile_X03_Y04_SB_T2_WEST_SB_IN_B17_ready;
	wire Tile_X03_Y04_SB_T2_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y04_SB_T2_WEST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y04_SB_T2_WEST_SB_OUT_B17;
	wire Tile_X03_Y04_SB_T2_WEST_SB_OUT_B17_valid;
	wire Tile_X03_Y04_SB_T2_WEST_SB_OUT_B1_valid;
	wire Tile_X03_Y04_SB_T3_EAST_SB_IN_B17_ready;
	wire Tile_X03_Y04_SB_T3_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y04_SB_T3_EAST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y04_SB_T3_EAST_SB_OUT_B17;
	wire Tile_X03_Y04_SB_T3_EAST_SB_OUT_B17_valid;
	wire Tile_X03_Y04_SB_T3_EAST_SB_OUT_B1_valid;
	wire Tile_X03_Y04_SB_T3_NORTH_SB_IN_B17_ready;
	wire Tile_X03_Y04_SB_T3_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B17;
	wire Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B17_valid;
	wire Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B1_valid;
	wire Tile_X03_Y04_SB_T3_SOUTH_SB_IN_B17_ready;
	wire Tile_X03_Y04_SB_T3_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y04_SB_T3_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y04_SB_T3_SOUTH_SB_OUT_B17;
	wire Tile_X03_Y04_SB_T3_SOUTH_SB_OUT_B17_valid;
	wire Tile_X03_Y04_SB_T3_SOUTH_SB_OUT_B1_valid;
	wire Tile_X03_Y04_SB_T3_WEST_SB_IN_B17_ready;
	wire Tile_X03_Y04_SB_T3_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y04_SB_T3_WEST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y04_SB_T3_WEST_SB_OUT_B17;
	wire Tile_X03_Y04_SB_T3_WEST_SB_OUT_B17_valid;
	wire Tile_X03_Y04_SB_T3_WEST_SB_OUT_B1_valid;
	wire Tile_X03_Y04_SB_T4_EAST_SB_IN_B17_ready;
	wire Tile_X03_Y04_SB_T4_EAST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y04_SB_T4_EAST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y04_SB_T4_EAST_SB_OUT_B17;
	wire Tile_X03_Y04_SB_T4_EAST_SB_OUT_B17_valid;
	wire Tile_X03_Y04_SB_T4_EAST_SB_OUT_B1_valid;
	wire Tile_X03_Y04_SB_T4_NORTH_SB_IN_B17_ready;
	wire Tile_X03_Y04_SB_T4_NORTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B17;
	wire Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B17_valid;
	wire Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B1_valid;
	wire Tile_X03_Y04_SB_T4_SOUTH_SB_IN_B17_ready;
	wire Tile_X03_Y04_SB_T4_SOUTH_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y04_SB_T4_SOUTH_SB_OUT_B1;
	wire [16:0] Tile_X03_Y04_SB_T4_SOUTH_SB_OUT_B17;
	wire Tile_X03_Y04_SB_T4_SOUTH_SB_OUT_B17_valid;
	wire Tile_X03_Y04_SB_T4_SOUTH_SB_OUT_B1_valid;
	wire Tile_X03_Y04_SB_T4_WEST_SB_IN_B17_ready;
	wire Tile_X03_Y04_SB_T4_WEST_SB_IN_B1_ready;
	wire [0:0] Tile_X03_Y04_SB_T4_WEST_SB_OUT_B1;
	wire [16:0] Tile_X03_Y04_SB_T4_WEST_SB_OUT_B17;
	wire Tile_X03_Y04_SB_T4_WEST_SB_OUT_B17_valid;
	wire Tile_X03_Y04_SB_T4_WEST_SB_OUT_B1_valid;
	wire Tile_X03_Y04_clk_out;
	wire [31:0] Tile_X03_Y04_config_out_config_addr;
	wire [31:0] Tile_X03_Y04_config_out_config_data;
	wire [0:0] Tile_X03_Y04_config_out_read;
	wire [0:0] Tile_X03_Y04_config_out_write;
	wire [0:0] Tile_X03_Y04_flush_out;
	wire [8:0] Tile_X03_Y04_hi;
	wire [7:0] Tile_X03_Y04_lo;
	wire [31:0] Tile_X03_Y04_read_config_data;
	wire Tile_X03_Y04_reset_out;
	wire [0:0] Tile_X03_Y04_stall_out;
	wire bit_const_0_None_out;
	wire [0:0] const_0_1_out;
	wire [16:0] const_0_17_out;
	wire [31:0] const_0_32_out;
	wire coreir_wrapInClock_inst0_out;
	wire coreir_wrapInClock_inst1_out;
	wire coreir_wrapInClock_inst2_out;
	wire [31:0] read_config_data_or_final_O;
	wire [3:0] self_stall_out;
	coreir_reg #(
		.clk_posedge(1'b1),
		.init(1'h0),
		.width(1)
	) PipelineRegister_inst0$Register_inst0$reg_P1_inst0(
		.clk(clk),
		.in(flush),
		.out(PipelineRegister_inst0$Register_inst0$reg_P1_inst0_out)
	);
	coreir_reg #(
		.clk_posedge(1'b1),
		.init(1'h0),
		.width(1)
	) PipelineRegister_inst1$Register_inst0$reg_P1_inst0(
		.clk(clk),
		.in(flush),
		.out(PipelineRegister_inst1$Register_inst0$reg_P1_inst0_out)
	);
	coreir_reg #(
		.clk_posedge(1'b1),
		.init(1'h0),
		.width(1)
	) PipelineRegister_inst2$Register_inst0$reg_P1_inst0(
		.clk(clk),
		.in(flush),
		.out(PipelineRegister_inst2$Register_inst0$reg_P1_inst0_out)
	);
	coreir_reg #(
		.clk_posedge(1'b1),
		.init(1'h0),
		.width(1)
	) PipelineRegister_inst3$Register_inst0$reg_P1_inst0(
		.clk(clk),
		.in(flush),
		.out(PipelineRegister_inst3$Register_inst0$reg_P1_inst0_out)
	);
	wire [65:0] PipelineRegister_inst4$Register_inst0$reg_P66_inst0_in;
	assign PipelineRegister_inst4$Register_inst0$reg_P66_inst0_in = {config_0_write[0], config_0_read[0], config_0_config_data, config_0_config_addr};
	coreir_reg #(
		.clk_posedge(1'b1),
		.init(66'h00000000000000000),
		.width(66)
	) PipelineRegister_inst4$Register_inst0$reg_P66_inst0(
		.clk(clk),
		.in(PipelineRegister_inst4$Register_inst0$reg_P66_inst0_in),
		.out(PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out)
	);
	wire [65:0] PipelineRegister_inst5$Register_inst0$reg_P66_inst0_in;
	assign PipelineRegister_inst5$Register_inst0$reg_P66_inst0_in = {config_1_write[0], config_1_read[0], config_1_config_data, config_1_config_addr};
	coreir_reg #(
		.clk_posedge(1'b1),
		.init(66'h00000000000000000),
		.width(66)
	) PipelineRegister_inst5$Register_inst0$reg_P66_inst0(
		.clk(clk),
		.in(PipelineRegister_inst5$Register_inst0$reg_P66_inst0_in),
		.out(PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out)
	);
	wire [65:0] PipelineRegister_inst6$Register_inst0$reg_P66_inst0_in;
	assign PipelineRegister_inst6$Register_inst0$reg_P66_inst0_in = {config_2_write[0], config_2_read[0], config_2_config_data, config_2_config_addr};
	coreir_reg #(
		.clk_posedge(1'b1),
		.init(66'h00000000000000000),
		.width(66)
	) PipelineRegister_inst6$Register_inst0$reg_P66_inst0(
		.clk(clk),
		.in(PipelineRegister_inst6$Register_inst0$reg_P66_inst0_in),
		.out(PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out)
	);
	wire [65:0] PipelineRegister_inst7$Register_inst0$reg_P66_inst0_in;
	assign PipelineRegister_inst7$Register_inst0$reg_P66_inst0_in = {config_3_write[0], config_3_read[0], config_3_config_data, config_3_config_addr};
	coreir_reg #(
		.clk_posedge(1'b1),
		.init(66'h00000000000000000),
		.width(66)
	) PipelineRegister_inst7$Register_inst0$reg_P66_inst0(
		.clk(clk),
		.in(PipelineRegister_inst7$Register_inst0$reg_P66_inst0_in),
		.out(PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out)
	);
	wire [31:0] Tile_X00_Y00_config_config_addr;
	assign Tile_X00_Y00_config_config_addr = {PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[31], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[30], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[29], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[28], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[27], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[26], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[25], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[24], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[23], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[22], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[21], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[20], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[19], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[18], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[17], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[16], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[15], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[14], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[13], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[12], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[11], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[10], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[9], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[8], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[7], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[6], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[5], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[4], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[3], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[2], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[1], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[0]};
	wire [31:0] Tile_X00_Y00_config_config_data;
	assign Tile_X00_Y00_config_config_data = {PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[63], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[62], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[61], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[60], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[59], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[58], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[57], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[56], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[55], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[54], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[53], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[52], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[51], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[50], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[49], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[48], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[47], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[46], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[45], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[44], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[43], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[42], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[41], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[40], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[39], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[38], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[37], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[36], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[35], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[34], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[33], PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[32]};
	wire [4:0] Tile_X00_Y00_io2f_17_ready;
	assign Tile_X00_Y00_io2f_17_ready = {Tile_X00_Y01_SB_T4_NORTH_SB_IN_B17_ready, Tile_X00_Y01_SB_T3_NORTH_SB_IN_B17_ready, Tile_X00_Y01_SB_T2_NORTH_SB_IN_B17_ready, Tile_X00_Y01_SB_T1_NORTH_SB_IN_B17_ready, Tile_X00_Y01_SB_T0_NORTH_SB_IN_B17_ready};
	wire [4:0] Tile_X00_Y00_io2f_1_ready;
	assign Tile_X00_Y00_io2f_1_ready = {Tile_X00_Y01_SB_T4_NORTH_SB_IN_B1_ready, Tile_X00_Y01_SB_T3_NORTH_SB_IN_B1_ready, Tile_X00_Y01_SB_T2_NORTH_SB_IN_B1_ready, Tile_X00_Y01_SB_T1_NORTH_SB_IN_B1_ready, Tile_X00_Y01_SB_T0_NORTH_SB_IN_B1_ready};
	wire [15:0] Tile_X00_Y00_tile_id;
	assign Tile_X00_Y00_tile_id = {Tile_X00_Y00_lo[7], Tile_X00_Y00_lo[7], Tile_X00_Y00_lo[6], Tile_X00_Y00_lo[6], Tile_X00_Y00_lo[5], Tile_X00_Y00_lo[5], Tile_X00_Y00_lo[4], Tile_X00_Y00_lo[4], Tile_X00_Y00_lo[3], Tile_X00_Y00_lo[3], Tile_X00_Y00_lo[2], Tile_X00_Y00_lo[2], Tile_X00_Y00_lo[1], Tile_X00_Y00_lo[1], Tile_X00_Y00_lo[0], Tile_X00_Y00_lo[0]};
	Tile_IOCoreReadyValid Tile_X00_Y00(
		.clk(clk),
		.clk_out(Tile_X00_Y00_clk_out),
		.config_config_addr(Tile_X00_Y00_config_config_addr),
		.config_config_data(Tile_X00_Y00_config_config_data),
		.config_out_config_addr(Tile_X00_Y00_config_out_config_addr),
		.config_out_config_data(Tile_X00_Y00_config_out_config_data),
		.config_out_read(Tile_X00_Y00_config_out_read),
		.config_out_write(Tile_X00_Y00_config_out_write),
		.config_read(PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[64]),
		.config_write(PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[65]),
		.f2io_1(Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B1),
		.f2io_17(Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B17),
		.f2io_17_ready(Tile_X00_Y00_f2io_17_ready),
		.f2io_17_valid(Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B17_valid),
		.f2io_1_ready(Tile_X00_Y00_f2io_1_ready),
		.f2io_1_valid(Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B1_valid),
		.flush(PipelineRegister_inst0$Register_inst0$reg_P1_inst0_out),
		.flush_out(Tile_X00_Y00_flush_out),
		.glb2io_1(glb2io_1_X00_Y00),
		.glb2io_17(glb2io_17_X00_Y00),
		.glb2io_17_ready(Tile_X00_Y00_glb2io_17_ready),
		.glb2io_17_valid(glb2io_17_X00_Y00_valid),
		.glb2io_1_ready(Tile_X00_Y00_glb2io_1_ready),
		.glb2io_1_valid(glb2io_1_X00_Y00_valid),
		.hi(Tile_X00_Y00_hi),
		.io2f_1(Tile_X00_Y00_io2f_1),
		.io2f_17(Tile_X00_Y00_io2f_17),
		.io2f_17_ready(Tile_X00_Y00_io2f_17_ready),
		.io2f_17_valid(Tile_X00_Y00_io2f_17_valid),
		.io2f_1_ready(Tile_X00_Y00_io2f_1_ready),
		.io2f_1_valid(Tile_X00_Y00_io2f_1_valid),
		.io2glb_1(Tile_X00_Y00_io2glb_1),
		.io2glb_17(Tile_X00_Y00_io2glb_17),
		.io2glb_17_ready(io2glb_17_X00_Y00_ready),
		.io2glb_17_valid(Tile_X00_Y00_io2glb_17_valid),
		.io2glb_1_ready(io2glb_1_X00_Y00_ready),
		.io2glb_1_valid(Tile_X00_Y00_io2glb_1_valid),
		.lo(Tile_X00_Y00_lo),
		.read_config_data(Tile_X00_Y00_read_config_data),
		.read_config_data_in(const_0_32_out),
		.reset(reset),
		.reset_out(Tile_X00_Y00_reset_out),
		.stall(self_stall_out[0:0]),
		.stall_out(Tile_X00_Y00_stall_out),
		.tile_id(Tile_X00_Y00_tile_id)
	);
	wire [15:0] Tile_X00_Y01_tile_id;
	assign Tile_X00_Y01_tile_id = {Tile_X00_Y01_lo[7], Tile_X00_Y01_lo[7], Tile_X00_Y01_lo[6], Tile_X00_Y01_lo[6], Tile_X00_Y01_lo[5], Tile_X00_Y01_lo[5], Tile_X00_Y01_lo[4], Tile_X00_Y01_lo[4], Tile_X00_Y01_lo[3], Tile_X00_Y01_lo[3], Tile_X00_Y01_lo[2], Tile_X00_Y01_lo[2], Tile_X00_Y01_lo[1], Tile_X00_Y01_lo[1], Tile_X00_Y01_lo[0], Tile_X00_Y01_hi[0]};
	Tile_PE Tile_X00_Y01(
		.SB_T0_EAST_SB_IN_B1(Tile_X01_Y01_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_EAST_SB_IN_B17(Tile_X01_Y01_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_EAST_SB_IN_B17_ready(Tile_X00_Y01_SB_T0_EAST_SB_IN_B17_ready),
		.SB_T0_EAST_SB_IN_B17_valid(Tile_X01_Y01_SB_T0_WEST_SB_OUT_B17_valid),
		.SB_T0_EAST_SB_IN_B1_ready(Tile_X00_Y01_SB_T0_EAST_SB_IN_B1_ready),
		.SB_T0_EAST_SB_IN_B1_valid(Tile_X01_Y01_SB_T0_WEST_SB_OUT_B1_valid),
		.SB_T0_EAST_SB_OUT_B1(Tile_X00_Y01_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_EAST_SB_OUT_B17(Tile_X00_Y01_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_EAST_SB_OUT_B17_ready(Tile_X01_Y01_SB_T0_WEST_SB_IN_B17_ready),
		.SB_T0_EAST_SB_OUT_B17_valid(Tile_X00_Y01_SB_T0_EAST_SB_OUT_B17_valid),
		.SB_T0_EAST_SB_OUT_B1_ready(Tile_X01_Y01_SB_T0_WEST_SB_IN_B1_ready),
		.SB_T0_EAST_SB_OUT_B1_valid(Tile_X00_Y01_SB_T0_EAST_SB_OUT_B1_valid),
		.SB_T0_NORTH_SB_IN_B1(Tile_X00_Y00_io2f_1),
		.SB_T0_NORTH_SB_IN_B17(Tile_X00_Y00_io2f_17),
		.SB_T0_NORTH_SB_IN_B17_ready(Tile_X00_Y01_SB_T0_NORTH_SB_IN_B17_ready),
		.SB_T0_NORTH_SB_IN_B17_valid(Tile_X00_Y00_io2f_17_valid),
		.SB_T0_NORTH_SB_IN_B1_ready(Tile_X00_Y01_SB_T0_NORTH_SB_IN_B1_ready),
		.SB_T0_NORTH_SB_IN_B1_valid(Tile_X00_Y00_io2f_1_valid),
		.SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_OUT_B17(Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_OUT_B17_ready(Tile_X00_Y00_f2io_17_ready),
		.SB_T0_NORTH_SB_OUT_B17_valid(Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B17_valid),
		.SB_T0_NORTH_SB_OUT_B1_ready(Tile_X00_Y00_f2io_1_ready),
		.SB_T0_NORTH_SB_OUT_B1_valid(Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B1_valid),
		.SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_IN_B17(Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_IN_B17_ready(Tile_X00_Y01_SB_T0_SOUTH_SB_IN_B17_ready),
		.SB_T0_SOUTH_SB_IN_B17_valid(Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B17_valid),
		.SB_T0_SOUTH_SB_IN_B1_ready(Tile_X00_Y01_SB_T0_SOUTH_SB_IN_B1_ready),
		.SB_T0_SOUTH_SB_IN_B1_valid(Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B1_valid),
		.SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_OUT_B17(Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_OUT_B17_ready(Tile_X00_Y02_SB_T0_NORTH_SB_IN_B17_ready),
		.SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B17_valid),
		.SB_T0_SOUTH_SB_OUT_B1_ready(Tile_X00_Y02_SB_T0_NORTH_SB_IN_B1_ready),
		.SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B1_valid),
		.SB_T0_WEST_SB_IN_B1(const_0_1_out),
		.SB_T0_WEST_SB_IN_B17(const_0_17_out),
		.SB_T0_WEST_SB_IN_B17_ready(Tile_X00_Y01_SB_T0_WEST_SB_IN_B17_ready),
		.SB_T0_WEST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T0_WEST_SB_IN_B1_ready(Tile_X00_Y01_SB_T0_WEST_SB_IN_B1_ready),
		.SB_T0_WEST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T0_WEST_SB_OUT_B1(Tile_X00_Y01_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_WEST_SB_OUT_B17(Tile_X00_Y01_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T0_WEST_SB_OUT_B17_valid(Tile_X00_Y01_SB_T0_WEST_SB_OUT_B17_valid),
		.SB_T0_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T0_WEST_SB_OUT_B1_valid(Tile_X00_Y01_SB_T0_WEST_SB_OUT_B1_valid),
		.SB_T1_EAST_SB_IN_B1(Tile_X01_Y01_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_EAST_SB_IN_B17(Tile_X01_Y01_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_EAST_SB_IN_B17_ready(Tile_X00_Y01_SB_T1_EAST_SB_IN_B17_ready),
		.SB_T1_EAST_SB_IN_B17_valid(Tile_X01_Y01_SB_T1_WEST_SB_OUT_B17_valid),
		.SB_T1_EAST_SB_IN_B1_ready(Tile_X00_Y01_SB_T1_EAST_SB_IN_B1_ready),
		.SB_T1_EAST_SB_IN_B1_valid(Tile_X01_Y01_SB_T1_WEST_SB_OUT_B1_valid),
		.SB_T1_EAST_SB_OUT_B1(Tile_X00_Y01_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_EAST_SB_OUT_B17(Tile_X00_Y01_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_EAST_SB_OUT_B17_ready(Tile_X01_Y01_SB_T1_WEST_SB_IN_B17_ready),
		.SB_T1_EAST_SB_OUT_B17_valid(Tile_X00_Y01_SB_T1_EAST_SB_OUT_B17_valid),
		.SB_T1_EAST_SB_OUT_B1_ready(Tile_X01_Y01_SB_T1_WEST_SB_IN_B1_ready),
		.SB_T1_EAST_SB_OUT_B1_valid(Tile_X00_Y01_SB_T1_EAST_SB_OUT_B1_valid),
		.SB_T1_NORTH_SB_IN_B1(Tile_X00_Y00_io2f_1),
		.SB_T1_NORTH_SB_IN_B17(Tile_X00_Y00_io2f_17),
		.SB_T1_NORTH_SB_IN_B17_ready(Tile_X00_Y01_SB_T1_NORTH_SB_IN_B17_ready),
		.SB_T1_NORTH_SB_IN_B17_valid(Tile_X00_Y00_io2f_17_valid),
		.SB_T1_NORTH_SB_IN_B1_ready(Tile_X00_Y01_SB_T1_NORTH_SB_IN_B1_ready),
		.SB_T1_NORTH_SB_IN_B1_valid(Tile_X00_Y00_io2f_1_valid),
		.SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y01_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_OUT_B17(Tile_X00_Y01_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T1_NORTH_SB_OUT_B17_valid(Tile_X00_Y01_SB_T1_NORTH_SB_OUT_B17_valid),
		.SB_T1_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T1_NORTH_SB_OUT_B1_valid(Tile_X00_Y01_SB_T1_NORTH_SB_OUT_B1_valid),
		.SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_IN_B17(Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_IN_B17_ready(Tile_X00_Y01_SB_T1_SOUTH_SB_IN_B17_ready),
		.SB_T1_SOUTH_SB_IN_B17_valid(Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B17_valid),
		.SB_T1_SOUTH_SB_IN_B1_ready(Tile_X00_Y01_SB_T1_SOUTH_SB_IN_B1_ready),
		.SB_T1_SOUTH_SB_IN_B1_valid(Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B1_valid),
		.SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_OUT_B17(Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_OUT_B17_ready(Tile_X00_Y02_SB_T1_NORTH_SB_IN_B17_ready),
		.SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B17_valid),
		.SB_T1_SOUTH_SB_OUT_B1_ready(Tile_X00_Y02_SB_T1_NORTH_SB_IN_B1_ready),
		.SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B1_valid),
		.SB_T1_WEST_SB_IN_B1(const_0_1_out),
		.SB_T1_WEST_SB_IN_B17(const_0_17_out),
		.SB_T1_WEST_SB_IN_B17_ready(Tile_X00_Y01_SB_T1_WEST_SB_IN_B17_ready),
		.SB_T1_WEST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T1_WEST_SB_IN_B1_ready(Tile_X00_Y01_SB_T1_WEST_SB_IN_B1_ready),
		.SB_T1_WEST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T1_WEST_SB_OUT_B1(Tile_X00_Y01_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_WEST_SB_OUT_B17(Tile_X00_Y01_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T1_WEST_SB_OUT_B17_valid(Tile_X00_Y01_SB_T1_WEST_SB_OUT_B17_valid),
		.SB_T1_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T1_WEST_SB_OUT_B1_valid(Tile_X00_Y01_SB_T1_WEST_SB_OUT_B1_valid),
		.SB_T2_EAST_SB_IN_B1(Tile_X01_Y01_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_EAST_SB_IN_B17(Tile_X01_Y01_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_EAST_SB_IN_B17_ready(Tile_X00_Y01_SB_T2_EAST_SB_IN_B17_ready),
		.SB_T2_EAST_SB_IN_B17_valid(Tile_X01_Y01_SB_T2_WEST_SB_OUT_B17_valid),
		.SB_T2_EAST_SB_IN_B1_ready(Tile_X00_Y01_SB_T2_EAST_SB_IN_B1_ready),
		.SB_T2_EAST_SB_IN_B1_valid(Tile_X01_Y01_SB_T2_WEST_SB_OUT_B1_valid),
		.SB_T2_EAST_SB_OUT_B1(Tile_X00_Y01_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_EAST_SB_OUT_B17(Tile_X00_Y01_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_EAST_SB_OUT_B17_ready(Tile_X01_Y01_SB_T2_WEST_SB_IN_B17_ready),
		.SB_T2_EAST_SB_OUT_B17_valid(Tile_X00_Y01_SB_T2_EAST_SB_OUT_B17_valid),
		.SB_T2_EAST_SB_OUT_B1_ready(Tile_X01_Y01_SB_T2_WEST_SB_IN_B1_ready),
		.SB_T2_EAST_SB_OUT_B1_valid(Tile_X00_Y01_SB_T2_EAST_SB_OUT_B1_valid),
		.SB_T2_NORTH_SB_IN_B1(Tile_X00_Y00_io2f_1),
		.SB_T2_NORTH_SB_IN_B17(Tile_X00_Y00_io2f_17),
		.SB_T2_NORTH_SB_IN_B17_ready(Tile_X00_Y01_SB_T2_NORTH_SB_IN_B17_ready),
		.SB_T2_NORTH_SB_IN_B17_valid(Tile_X00_Y00_io2f_17_valid),
		.SB_T2_NORTH_SB_IN_B1_ready(Tile_X00_Y01_SB_T2_NORTH_SB_IN_B1_ready),
		.SB_T2_NORTH_SB_IN_B1_valid(Tile_X00_Y00_io2f_1_valid),
		.SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y01_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_OUT_B17(Tile_X00_Y01_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T2_NORTH_SB_OUT_B17_valid(Tile_X00_Y01_SB_T2_NORTH_SB_OUT_B17_valid),
		.SB_T2_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T2_NORTH_SB_OUT_B1_valid(Tile_X00_Y01_SB_T2_NORTH_SB_OUT_B1_valid),
		.SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_IN_B17(Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_IN_B17_ready(Tile_X00_Y01_SB_T2_SOUTH_SB_IN_B17_ready),
		.SB_T2_SOUTH_SB_IN_B17_valid(Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B17_valid),
		.SB_T2_SOUTH_SB_IN_B1_ready(Tile_X00_Y01_SB_T2_SOUTH_SB_IN_B1_ready),
		.SB_T2_SOUTH_SB_IN_B1_valid(Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B1_valid),
		.SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_OUT_B17(Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_OUT_B17_ready(Tile_X00_Y02_SB_T2_NORTH_SB_IN_B17_ready),
		.SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B17_valid),
		.SB_T2_SOUTH_SB_OUT_B1_ready(Tile_X00_Y02_SB_T2_NORTH_SB_IN_B1_ready),
		.SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B1_valid),
		.SB_T2_WEST_SB_IN_B1(const_0_1_out),
		.SB_T2_WEST_SB_IN_B17(const_0_17_out),
		.SB_T2_WEST_SB_IN_B17_ready(Tile_X00_Y01_SB_T2_WEST_SB_IN_B17_ready),
		.SB_T2_WEST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T2_WEST_SB_IN_B1_ready(Tile_X00_Y01_SB_T2_WEST_SB_IN_B1_ready),
		.SB_T2_WEST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T2_WEST_SB_OUT_B1(Tile_X00_Y01_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_WEST_SB_OUT_B17(Tile_X00_Y01_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T2_WEST_SB_OUT_B17_valid(Tile_X00_Y01_SB_T2_WEST_SB_OUT_B17_valid),
		.SB_T2_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T2_WEST_SB_OUT_B1_valid(Tile_X00_Y01_SB_T2_WEST_SB_OUT_B1_valid),
		.SB_T3_EAST_SB_IN_B1(Tile_X01_Y01_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_EAST_SB_IN_B17(Tile_X01_Y01_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_EAST_SB_IN_B17_ready(Tile_X00_Y01_SB_T3_EAST_SB_IN_B17_ready),
		.SB_T3_EAST_SB_IN_B17_valid(Tile_X01_Y01_SB_T3_WEST_SB_OUT_B17_valid),
		.SB_T3_EAST_SB_IN_B1_ready(Tile_X00_Y01_SB_T3_EAST_SB_IN_B1_ready),
		.SB_T3_EAST_SB_IN_B1_valid(Tile_X01_Y01_SB_T3_WEST_SB_OUT_B1_valid),
		.SB_T3_EAST_SB_OUT_B1(Tile_X00_Y01_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_EAST_SB_OUT_B17(Tile_X00_Y01_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_EAST_SB_OUT_B17_ready(Tile_X01_Y01_SB_T3_WEST_SB_IN_B17_ready),
		.SB_T3_EAST_SB_OUT_B17_valid(Tile_X00_Y01_SB_T3_EAST_SB_OUT_B17_valid),
		.SB_T3_EAST_SB_OUT_B1_ready(Tile_X01_Y01_SB_T3_WEST_SB_IN_B1_ready),
		.SB_T3_EAST_SB_OUT_B1_valid(Tile_X00_Y01_SB_T3_EAST_SB_OUT_B1_valid),
		.SB_T3_NORTH_SB_IN_B1(Tile_X00_Y00_io2f_1),
		.SB_T3_NORTH_SB_IN_B17(Tile_X00_Y00_io2f_17),
		.SB_T3_NORTH_SB_IN_B17_ready(Tile_X00_Y01_SB_T3_NORTH_SB_IN_B17_ready),
		.SB_T3_NORTH_SB_IN_B17_valid(Tile_X00_Y00_io2f_17_valid),
		.SB_T3_NORTH_SB_IN_B1_ready(Tile_X00_Y01_SB_T3_NORTH_SB_IN_B1_ready),
		.SB_T3_NORTH_SB_IN_B1_valid(Tile_X00_Y00_io2f_1_valid),
		.SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y01_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_OUT_B17(Tile_X00_Y01_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T3_NORTH_SB_OUT_B17_valid(Tile_X00_Y01_SB_T3_NORTH_SB_OUT_B17_valid),
		.SB_T3_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T3_NORTH_SB_OUT_B1_valid(Tile_X00_Y01_SB_T3_NORTH_SB_OUT_B1_valid),
		.SB_T3_SOUTH_SB_IN_B1(Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_IN_B17(Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_IN_B17_ready(Tile_X00_Y01_SB_T3_SOUTH_SB_IN_B17_ready),
		.SB_T3_SOUTH_SB_IN_B17_valid(Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B17_valid),
		.SB_T3_SOUTH_SB_IN_B1_ready(Tile_X00_Y01_SB_T3_SOUTH_SB_IN_B1_ready),
		.SB_T3_SOUTH_SB_IN_B1_valid(Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B1_valid),
		.SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_OUT_B17(Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_OUT_B17_ready(Tile_X00_Y02_SB_T3_NORTH_SB_IN_B17_ready),
		.SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B17_valid),
		.SB_T3_SOUTH_SB_OUT_B1_ready(Tile_X00_Y02_SB_T3_NORTH_SB_IN_B1_ready),
		.SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B1_valid),
		.SB_T3_WEST_SB_IN_B1(const_0_1_out),
		.SB_T3_WEST_SB_IN_B17(const_0_17_out),
		.SB_T3_WEST_SB_IN_B17_ready(Tile_X00_Y01_SB_T3_WEST_SB_IN_B17_ready),
		.SB_T3_WEST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T3_WEST_SB_IN_B1_ready(Tile_X00_Y01_SB_T3_WEST_SB_IN_B1_ready),
		.SB_T3_WEST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T3_WEST_SB_OUT_B1(Tile_X00_Y01_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_WEST_SB_OUT_B17(Tile_X00_Y01_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T3_WEST_SB_OUT_B17_valid(Tile_X00_Y01_SB_T3_WEST_SB_OUT_B17_valid),
		.SB_T3_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T3_WEST_SB_OUT_B1_valid(Tile_X00_Y01_SB_T3_WEST_SB_OUT_B1_valid),
		.SB_T4_EAST_SB_IN_B1(Tile_X01_Y01_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_EAST_SB_IN_B17(Tile_X01_Y01_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_EAST_SB_IN_B17_ready(Tile_X00_Y01_SB_T4_EAST_SB_IN_B17_ready),
		.SB_T4_EAST_SB_IN_B17_valid(Tile_X01_Y01_SB_T4_WEST_SB_OUT_B17_valid),
		.SB_T4_EAST_SB_IN_B1_ready(Tile_X00_Y01_SB_T4_EAST_SB_IN_B1_ready),
		.SB_T4_EAST_SB_IN_B1_valid(Tile_X01_Y01_SB_T4_WEST_SB_OUT_B1_valid),
		.SB_T4_EAST_SB_OUT_B1(Tile_X00_Y01_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_EAST_SB_OUT_B17(Tile_X00_Y01_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_EAST_SB_OUT_B17_ready(Tile_X01_Y01_SB_T4_WEST_SB_IN_B17_ready),
		.SB_T4_EAST_SB_OUT_B17_valid(Tile_X00_Y01_SB_T4_EAST_SB_OUT_B17_valid),
		.SB_T4_EAST_SB_OUT_B1_ready(Tile_X01_Y01_SB_T4_WEST_SB_IN_B1_ready),
		.SB_T4_EAST_SB_OUT_B1_valid(Tile_X00_Y01_SB_T4_EAST_SB_OUT_B1_valid),
		.SB_T4_NORTH_SB_IN_B1(Tile_X00_Y00_io2f_1),
		.SB_T4_NORTH_SB_IN_B17(Tile_X00_Y00_io2f_17),
		.SB_T4_NORTH_SB_IN_B17_ready(Tile_X00_Y01_SB_T4_NORTH_SB_IN_B17_ready),
		.SB_T4_NORTH_SB_IN_B17_valid(Tile_X00_Y00_io2f_17_valid),
		.SB_T4_NORTH_SB_IN_B1_ready(Tile_X00_Y01_SB_T4_NORTH_SB_IN_B1_ready),
		.SB_T4_NORTH_SB_IN_B1_valid(Tile_X00_Y00_io2f_1_valid),
		.SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y01_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_OUT_B17(Tile_X00_Y01_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T4_NORTH_SB_OUT_B17_valid(Tile_X00_Y01_SB_T4_NORTH_SB_OUT_B17_valid),
		.SB_T4_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T4_NORTH_SB_OUT_B1_valid(Tile_X00_Y01_SB_T4_NORTH_SB_OUT_B1_valid),
		.SB_T4_SOUTH_SB_IN_B1(Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_IN_B17(Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_IN_B17_ready(Tile_X00_Y01_SB_T4_SOUTH_SB_IN_B17_ready),
		.SB_T4_SOUTH_SB_IN_B17_valid(Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B17_valid),
		.SB_T4_SOUTH_SB_IN_B1_ready(Tile_X00_Y01_SB_T4_SOUTH_SB_IN_B1_ready),
		.SB_T4_SOUTH_SB_IN_B1_valid(Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B1_valid),
		.SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_OUT_B17(Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_OUT_B17_ready(Tile_X00_Y02_SB_T4_NORTH_SB_IN_B17_ready),
		.SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B17_valid),
		.SB_T4_SOUTH_SB_OUT_B1_ready(Tile_X00_Y02_SB_T4_NORTH_SB_IN_B1_ready),
		.SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B1_valid),
		.SB_T4_WEST_SB_IN_B1(const_0_1_out),
		.SB_T4_WEST_SB_IN_B17(const_0_17_out),
		.SB_T4_WEST_SB_IN_B17_ready(Tile_X00_Y01_SB_T4_WEST_SB_IN_B17_ready),
		.SB_T4_WEST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T4_WEST_SB_IN_B1_ready(Tile_X00_Y01_SB_T4_WEST_SB_IN_B1_ready),
		.SB_T4_WEST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T4_WEST_SB_OUT_B1(Tile_X00_Y01_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_WEST_SB_OUT_B17(Tile_X00_Y01_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T4_WEST_SB_OUT_B17_valid(Tile_X00_Y01_SB_T4_WEST_SB_OUT_B17_valid),
		.SB_T4_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T4_WEST_SB_OUT_B1_valid(Tile_X00_Y01_SB_T4_WEST_SB_OUT_B1_valid),
		.clk(Tile_X00_Y00_clk_out),
		.clk_out(Tile_X00_Y01_clk_out),
		.clk_pass_through(coreir_wrapInClock_inst0_out),
		.clk_pass_through_out_bot(Tile_X00_Y01_clk_pass_through_out_bot),
		.clk_pass_through_out_right(Tile_X00_Y01_clk_pass_through_out_right),
		.config_config_addr(Tile_X00_Y00_config_out_config_addr),
		.config_config_data(Tile_X00_Y00_config_out_config_data),
		.config_out_config_addr(Tile_X00_Y01_config_out_config_addr),
		.config_out_config_data(Tile_X00_Y01_config_out_config_data),
		.config_out_read(Tile_X00_Y01_config_out_read),
		.config_out_write(Tile_X00_Y01_config_out_write),
		.config_read(Tile_X00_Y00_config_out_read),
		.config_write(Tile_X00_Y00_config_out_write),
		.flush(Tile_X00_Y00_flush_out),
		.flush_out(Tile_X00_Y01_flush_out),
		.hi(Tile_X00_Y01_hi),
		.lo(Tile_X00_Y01_lo),
		.read_config_data(Tile_X00_Y01_read_config_data),
		.read_config_data_in(Tile_X00_Y00_read_config_data),
		.reset(Tile_X00_Y00_reset_out),
		.reset_out(Tile_X00_Y01_reset_out),
		.stall(Tile_X00_Y00_stall_out),
		.stall_out(Tile_X00_Y01_stall_out),
		.tile_id(Tile_X00_Y01_tile_id)
	);
	wire [15:0] Tile_X00_Y02_tile_id;
	assign Tile_X00_Y02_tile_id = {Tile_X00_Y02_lo[7], Tile_X00_Y02_lo[7], Tile_X00_Y02_lo[6], Tile_X00_Y02_lo[6], Tile_X00_Y02_lo[5], Tile_X00_Y02_lo[5], Tile_X00_Y02_lo[4], Tile_X00_Y02_lo[4], Tile_X00_Y02_lo[3], Tile_X00_Y02_lo[3], Tile_X00_Y02_lo[2], Tile_X00_Y02_lo[2], Tile_X00_Y02_lo[1], Tile_X00_Y02_lo[1], Tile_X00_Y02_hi[1], Tile_X00_Y02_lo[0]};
	Tile_PE Tile_X00_Y02(
		.SB_T0_EAST_SB_IN_B1(Tile_X01_Y02_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_EAST_SB_IN_B17(Tile_X01_Y02_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_EAST_SB_IN_B17_ready(Tile_X00_Y02_SB_T0_EAST_SB_IN_B17_ready),
		.SB_T0_EAST_SB_IN_B17_valid(Tile_X01_Y02_SB_T0_WEST_SB_OUT_B17_valid),
		.SB_T0_EAST_SB_IN_B1_ready(Tile_X00_Y02_SB_T0_EAST_SB_IN_B1_ready),
		.SB_T0_EAST_SB_IN_B1_valid(Tile_X01_Y02_SB_T0_WEST_SB_OUT_B1_valid),
		.SB_T0_EAST_SB_OUT_B1(Tile_X00_Y02_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_EAST_SB_OUT_B17(Tile_X00_Y02_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_EAST_SB_OUT_B17_ready(Tile_X01_Y02_SB_T0_WEST_SB_IN_B17_ready),
		.SB_T0_EAST_SB_OUT_B17_valid(Tile_X00_Y02_SB_T0_EAST_SB_OUT_B17_valid),
		.SB_T0_EAST_SB_OUT_B1_ready(Tile_X01_Y02_SB_T0_WEST_SB_IN_B1_ready),
		.SB_T0_EAST_SB_OUT_B1_valid(Tile_X00_Y02_SB_T0_EAST_SB_OUT_B1_valid),
		.SB_T0_NORTH_SB_IN_B1(Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_IN_B17(Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_IN_B17_ready(Tile_X00_Y02_SB_T0_NORTH_SB_IN_B17_ready),
		.SB_T0_NORTH_SB_IN_B17_valid(Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B17_valid),
		.SB_T0_NORTH_SB_IN_B1_ready(Tile_X00_Y02_SB_T0_NORTH_SB_IN_B1_ready),
		.SB_T0_NORTH_SB_IN_B1_valid(Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B1_valid),
		.SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_OUT_B17(Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_OUT_B17_ready(Tile_X00_Y01_SB_T0_SOUTH_SB_IN_B17_ready),
		.SB_T0_NORTH_SB_OUT_B17_valid(Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B17_valid),
		.SB_T0_NORTH_SB_OUT_B1_ready(Tile_X00_Y01_SB_T0_SOUTH_SB_IN_B1_ready),
		.SB_T0_NORTH_SB_OUT_B1_valid(Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B1_valid),
		.SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_IN_B17(Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_IN_B17_ready(Tile_X00_Y02_SB_T0_SOUTH_SB_IN_B17_ready),
		.SB_T0_SOUTH_SB_IN_B17_valid(Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B17_valid),
		.SB_T0_SOUTH_SB_IN_B1_ready(Tile_X00_Y02_SB_T0_SOUTH_SB_IN_B1_ready),
		.SB_T0_SOUTH_SB_IN_B1_valid(Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B1_valid),
		.SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_OUT_B17(Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_OUT_B17_ready(Tile_X00_Y03_SB_T0_NORTH_SB_IN_B17_ready),
		.SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B17_valid),
		.SB_T0_SOUTH_SB_OUT_B1_ready(Tile_X00_Y03_SB_T0_NORTH_SB_IN_B1_ready),
		.SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B1_valid),
		.SB_T0_WEST_SB_IN_B1(const_0_1_out),
		.SB_T0_WEST_SB_IN_B17(const_0_17_out),
		.SB_T0_WEST_SB_IN_B17_ready(Tile_X00_Y02_SB_T0_WEST_SB_IN_B17_ready),
		.SB_T0_WEST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T0_WEST_SB_IN_B1_ready(Tile_X00_Y02_SB_T0_WEST_SB_IN_B1_ready),
		.SB_T0_WEST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T0_WEST_SB_OUT_B1(Tile_X00_Y02_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_WEST_SB_OUT_B17(Tile_X00_Y02_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T0_WEST_SB_OUT_B17_valid(Tile_X00_Y02_SB_T0_WEST_SB_OUT_B17_valid),
		.SB_T0_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T0_WEST_SB_OUT_B1_valid(Tile_X00_Y02_SB_T0_WEST_SB_OUT_B1_valid),
		.SB_T1_EAST_SB_IN_B1(Tile_X01_Y02_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_EAST_SB_IN_B17(Tile_X01_Y02_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_EAST_SB_IN_B17_ready(Tile_X00_Y02_SB_T1_EAST_SB_IN_B17_ready),
		.SB_T1_EAST_SB_IN_B17_valid(Tile_X01_Y02_SB_T1_WEST_SB_OUT_B17_valid),
		.SB_T1_EAST_SB_IN_B1_ready(Tile_X00_Y02_SB_T1_EAST_SB_IN_B1_ready),
		.SB_T1_EAST_SB_IN_B1_valid(Tile_X01_Y02_SB_T1_WEST_SB_OUT_B1_valid),
		.SB_T1_EAST_SB_OUT_B1(Tile_X00_Y02_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_EAST_SB_OUT_B17(Tile_X00_Y02_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_EAST_SB_OUT_B17_ready(Tile_X01_Y02_SB_T1_WEST_SB_IN_B17_ready),
		.SB_T1_EAST_SB_OUT_B17_valid(Tile_X00_Y02_SB_T1_EAST_SB_OUT_B17_valid),
		.SB_T1_EAST_SB_OUT_B1_ready(Tile_X01_Y02_SB_T1_WEST_SB_IN_B1_ready),
		.SB_T1_EAST_SB_OUT_B1_valid(Tile_X00_Y02_SB_T1_EAST_SB_OUT_B1_valid),
		.SB_T1_NORTH_SB_IN_B1(Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_IN_B17(Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_IN_B17_ready(Tile_X00_Y02_SB_T1_NORTH_SB_IN_B17_ready),
		.SB_T1_NORTH_SB_IN_B17_valid(Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B17_valid),
		.SB_T1_NORTH_SB_IN_B1_ready(Tile_X00_Y02_SB_T1_NORTH_SB_IN_B1_ready),
		.SB_T1_NORTH_SB_IN_B1_valid(Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B1_valid),
		.SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_OUT_B17(Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_OUT_B17_ready(Tile_X00_Y01_SB_T1_SOUTH_SB_IN_B17_ready),
		.SB_T1_NORTH_SB_OUT_B17_valid(Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B17_valid),
		.SB_T1_NORTH_SB_OUT_B1_ready(Tile_X00_Y01_SB_T1_SOUTH_SB_IN_B1_ready),
		.SB_T1_NORTH_SB_OUT_B1_valid(Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B1_valid),
		.SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_IN_B17(Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_IN_B17_ready(Tile_X00_Y02_SB_T1_SOUTH_SB_IN_B17_ready),
		.SB_T1_SOUTH_SB_IN_B17_valid(Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B17_valid),
		.SB_T1_SOUTH_SB_IN_B1_ready(Tile_X00_Y02_SB_T1_SOUTH_SB_IN_B1_ready),
		.SB_T1_SOUTH_SB_IN_B1_valid(Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B1_valid),
		.SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_OUT_B17(Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_OUT_B17_ready(Tile_X00_Y03_SB_T1_NORTH_SB_IN_B17_ready),
		.SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B17_valid),
		.SB_T1_SOUTH_SB_OUT_B1_ready(Tile_X00_Y03_SB_T1_NORTH_SB_IN_B1_ready),
		.SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B1_valid),
		.SB_T1_WEST_SB_IN_B1(const_0_1_out),
		.SB_T1_WEST_SB_IN_B17(const_0_17_out),
		.SB_T1_WEST_SB_IN_B17_ready(Tile_X00_Y02_SB_T1_WEST_SB_IN_B17_ready),
		.SB_T1_WEST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T1_WEST_SB_IN_B1_ready(Tile_X00_Y02_SB_T1_WEST_SB_IN_B1_ready),
		.SB_T1_WEST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T1_WEST_SB_OUT_B1(Tile_X00_Y02_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_WEST_SB_OUT_B17(Tile_X00_Y02_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T1_WEST_SB_OUT_B17_valid(Tile_X00_Y02_SB_T1_WEST_SB_OUT_B17_valid),
		.SB_T1_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T1_WEST_SB_OUT_B1_valid(Tile_X00_Y02_SB_T1_WEST_SB_OUT_B1_valid),
		.SB_T2_EAST_SB_IN_B1(Tile_X01_Y02_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_EAST_SB_IN_B17(Tile_X01_Y02_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_EAST_SB_IN_B17_ready(Tile_X00_Y02_SB_T2_EAST_SB_IN_B17_ready),
		.SB_T2_EAST_SB_IN_B17_valid(Tile_X01_Y02_SB_T2_WEST_SB_OUT_B17_valid),
		.SB_T2_EAST_SB_IN_B1_ready(Tile_X00_Y02_SB_T2_EAST_SB_IN_B1_ready),
		.SB_T2_EAST_SB_IN_B1_valid(Tile_X01_Y02_SB_T2_WEST_SB_OUT_B1_valid),
		.SB_T2_EAST_SB_OUT_B1(Tile_X00_Y02_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_EAST_SB_OUT_B17(Tile_X00_Y02_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_EAST_SB_OUT_B17_ready(Tile_X01_Y02_SB_T2_WEST_SB_IN_B17_ready),
		.SB_T2_EAST_SB_OUT_B17_valid(Tile_X00_Y02_SB_T2_EAST_SB_OUT_B17_valid),
		.SB_T2_EAST_SB_OUT_B1_ready(Tile_X01_Y02_SB_T2_WEST_SB_IN_B1_ready),
		.SB_T2_EAST_SB_OUT_B1_valid(Tile_X00_Y02_SB_T2_EAST_SB_OUT_B1_valid),
		.SB_T2_NORTH_SB_IN_B1(Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_IN_B17(Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_IN_B17_ready(Tile_X00_Y02_SB_T2_NORTH_SB_IN_B17_ready),
		.SB_T2_NORTH_SB_IN_B17_valid(Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B17_valid),
		.SB_T2_NORTH_SB_IN_B1_ready(Tile_X00_Y02_SB_T2_NORTH_SB_IN_B1_ready),
		.SB_T2_NORTH_SB_IN_B1_valid(Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B1_valid),
		.SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_OUT_B17(Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_OUT_B17_ready(Tile_X00_Y01_SB_T2_SOUTH_SB_IN_B17_ready),
		.SB_T2_NORTH_SB_OUT_B17_valid(Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B17_valid),
		.SB_T2_NORTH_SB_OUT_B1_ready(Tile_X00_Y01_SB_T2_SOUTH_SB_IN_B1_ready),
		.SB_T2_NORTH_SB_OUT_B1_valid(Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B1_valid),
		.SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_IN_B17(Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_IN_B17_ready(Tile_X00_Y02_SB_T2_SOUTH_SB_IN_B17_ready),
		.SB_T2_SOUTH_SB_IN_B17_valid(Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B17_valid),
		.SB_T2_SOUTH_SB_IN_B1_ready(Tile_X00_Y02_SB_T2_SOUTH_SB_IN_B1_ready),
		.SB_T2_SOUTH_SB_IN_B1_valid(Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B1_valid),
		.SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_OUT_B17(Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_OUT_B17_ready(Tile_X00_Y03_SB_T2_NORTH_SB_IN_B17_ready),
		.SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B17_valid),
		.SB_T2_SOUTH_SB_OUT_B1_ready(Tile_X00_Y03_SB_T2_NORTH_SB_IN_B1_ready),
		.SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B1_valid),
		.SB_T2_WEST_SB_IN_B1(const_0_1_out),
		.SB_T2_WEST_SB_IN_B17(const_0_17_out),
		.SB_T2_WEST_SB_IN_B17_ready(Tile_X00_Y02_SB_T2_WEST_SB_IN_B17_ready),
		.SB_T2_WEST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T2_WEST_SB_IN_B1_ready(Tile_X00_Y02_SB_T2_WEST_SB_IN_B1_ready),
		.SB_T2_WEST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T2_WEST_SB_OUT_B1(Tile_X00_Y02_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_WEST_SB_OUT_B17(Tile_X00_Y02_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T2_WEST_SB_OUT_B17_valid(Tile_X00_Y02_SB_T2_WEST_SB_OUT_B17_valid),
		.SB_T2_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T2_WEST_SB_OUT_B1_valid(Tile_X00_Y02_SB_T2_WEST_SB_OUT_B1_valid),
		.SB_T3_EAST_SB_IN_B1(Tile_X01_Y02_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_EAST_SB_IN_B17(Tile_X01_Y02_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_EAST_SB_IN_B17_ready(Tile_X00_Y02_SB_T3_EAST_SB_IN_B17_ready),
		.SB_T3_EAST_SB_IN_B17_valid(Tile_X01_Y02_SB_T3_WEST_SB_OUT_B17_valid),
		.SB_T3_EAST_SB_IN_B1_ready(Tile_X00_Y02_SB_T3_EAST_SB_IN_B1_ready),
		.SB_T3_EAST_SB_IN_B1_valid(Tile_X01_Y02_SB_T3_WEST_SB_OUT_B1_valid),
		.SB_T3_EAST_SB_OUT_B1(Tile_X00_Y02_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_EAST_SB_OUT_B17(Tile_X00_Y02_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_EAST_SB_OUT_B17_ready(Tile_X01_Y02_SB_T3_WEST_SB_IN_B17_ready),
		.SB_T3_EAST_SB_OUT_B17_valid(Tile_X00_Y02_SB_T3_EAST_SB_OUT_B17_valid),
		.SB_T3_EAST_SB_OUT_B1_ready(Tile_X01_Y02_SB_T3_WEST_SB_IN_B1_ready),
		.SB_T3_EAST_SB_OUT_B1_valid(Tile_X00_Y02_SB_T3_EAST_SB_OUT_B1_valid),
		.SB_T3_NORTH_SB_IN_B1(Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_IN_B17(Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_IN_B17_ready(Tile_X00_Y02_SB_T3_NORTH_SB_IN_B17_ready),
		.SB_T3_NORTH_SB_IN_B17_valid(Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B17_valid),
		.SB_T3_NORTH_SB_IN_B1_ready(Tile_X00_Y02_SB_T3_NORTH_SB_IN_B1_ready),
		.SB_T3_NORTH_SB_IN_B1_valid(Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B1_valid),
		.SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_OUT_B17(Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_OUT_B17_ready(Tile_X00_Y01_SB_T3_SOUTH_SB_IN_B17_ready),
		.SB_T3_NORTH_SB_OUT_B17_valid(Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B17_valid),
		.SB_T3_NORTH_SB_OUT_B1_ready(Tile_X00_Y01_SB_T3_SOUTH_SB_IN_B1_ready),
		.SB_T3_NORTH_SB_OUT_B1_valid(Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B1_valid),
		.SB_T3_SOUTH_SB_IN_B1(Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_IN_B17(Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_IN_B17_ready(Tile_X00_Y02_SB_T3_SOUTH_SB_IN_B17_ready),
		.SB_T3_SOUTH_SB_IN_B17_valid(Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B17_valid),
		.SB_T3_SOUTH_SB_IN_B1_ready(Tile_X00_Y02_SB_T3_SOUTH_SB_IN_B1_ready),
		.SB_T3_SOUTH_SB_IN_B1_valid(Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B1_valid),
		.SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_OUT_B17(Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_OUT_B17_ready(Tile_X00_Y03_SB_T3_NORTH_SB_IN_B17_ready),
		.SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B17_valid),
		.SB_T3_SOUTH_SB_OUT_B1_ready(Tile_X00_Y03_SB_T3_NORTH_SB_IN_B1_ready),
		.SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B1_valid),
		.SB_T3_WEST_SB_IN_B1(const_0_1_out),
		.SB_T3_WEST_SB_IN_B17(const_0_17_out),
		.SB_T3_WEST_SB_IN_B17_ready(Tile_X00_Y02_SB_T3_WEST_SB_IN_B17_ready),
		.SB_T3_WEST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T3_WEST_SB_IN_B1_ready(Tile_X00_Y02_SB_T3_WEST_SB_IN_B1_ready),
		.SB_T3_WEST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T3_WEST_SB_OUT_B1(Tile_X00_Y02_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_WEST_SB_OUT_B17(Tile_X00_Y02_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T3_WEST_SB_OUT_B17_valid(Tile_X00_Y02_SB_T3_WEST_SB_OUT_B17_valid),
		.SB_T3_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T3_WEST_SB_OUT_B1_valid(Tile_X00_Y02_SB_T3_WEST_SB_OUT_B1_valid),
		.SB_T4_EAST_SB_IN_B1(Tile_X01_Y02_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_EAST_SB_IN_B17(Tile_X01_Y02_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_EAST_SB_IN_B17_ready(Tile_X00_Y02_SB_T4_EAST_SB_IN_B17_ready),
		.SB_T4_EAST_SB_IN_B17_valid(Tile_X01_Y02_SB_T4_WEST_SB_OUT_B17_valid),
		.SB_T4_EAST_SB_IN_B1_ready(Tile_X00_Y02_SB_T4_EAST_SB_IN_B1_ready),
		.SB_T4_EAST_SB_IN_B1_valid(Tile_X01_Y02_SB_T4_WEST_SB_OUT_B1_valid),
		.SB_T4_EAST_SB_OUT_B1(Tile_X00_Y02_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_EAST_SB_OUT_B17(Tile_X00_Y02_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_EAST_SB_OUT_B17_ready(Tile_X01_Y02_SB_T4_WEST_SB_IN_B17_ready),
		.SB_T4_EAST_SB_OUT_B17_valid(Tile_X00_Y02_SB_T4_EAST_SB_OUT_B17_valid),
		.SB_T4_EAST_SB_OUT_B1_ready(Tile_X01_Y02_SB_T4_WEST_SB_IN_B1_ready),
		.SB_T4_EAST_SB_OUT_B1_valid(Tile_X00_Y02_SB_T4_EAST_SB_OUT_B1_valid),
		.SB_T4_NORTH_SB_IN_B1(Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_IN_B17(Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_IN_B17_ready(Tile_X00_Y02_SB_T4_NORTH_SB_IN_B17_ready),
		.SB_T4_NORTH_SB_IN_B17_valid(Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B17_valid),
		.SB_T4_NORTH_SB_IN_B1_ready(Tile_X00_Y02_SB_T4_NORTH_SB_IN_B1_ready),
		.SB_T4_NORTH_SB_IN_B1_valid(Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B1_valid),
		.SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_OUT_B17(Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_OUT_B17_ready(Tile_X00_Y01_SB_T4_SOUTH_SB_IN_B17_ready),
		.SB_T4_NORTH_SB_OUT_B17_valid(Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B17_valid),
		.SB_T4_NORTH_SB_OUT_B1_ready(Tile_X00_Y01_SB_T4_SOUTH_SB_IN_B1_ready),
		.SB_T4_NORTH_SB_OUT_B1_valid(Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B1_valid),
		.SB_T4_SOUTH_SB_IN_B1(Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_IN_B17(Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_IN_B17_ready(Tile_X00_Y02_SB_T4_SOUTH_SB_IN_B17_ready),
		.SB_T4_SOUTH_SB_IN_B17_valid(Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B17_valid),
		.SB_T4_SOUTH_SB_IN_B1_ready(Tile_X00_Y02_SB_T4_SOUTH_SB_IN_B1_ready),
		.SB_T4_SOUTH_SB_IN_B1_valid(Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B1_valid),
		.SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_OUT_B17(Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_OUT_B17_ready(Tile_X00_Y03_SB_T4_NORTH_SB_IN_B17_ready),
		.SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B17_valid),
		.SB_T4_SOUTH_SB_OUT_B1_ready(Tile_X00_Y03_SB_T4_NORTH_SB_IN_B1_ready),
		.SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B1_valid),
		.SB_T4_WEST_SB_IN_B1(const_0_1_out),
		.SB_T4_WEST_SB_IN_B17(const_0_17_out),
		.SB_T4_WEST_SB_IN_B17_ready(Tile_X00_Y02_SB_T4_WEST_SB_IN_B17_ready),
		.SB_T4_WEST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T4_WEST_SB_IN_B1_ready(Tile_X00_Y02_SB_T4_WEST_SB_IN_B1_ready),
		.SB_T4_WEST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T4_WEST_SB_OUT_B1(Tile_X00_Y02_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_WEST_SB_OUT_B17(Tile_X00_Y02_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T4_WEST_SB_OUT_B17_valid(Tile_X00_Y02_SB_T4_WEST_SB_OUT_B17_valid),
		.SB_T4_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T4_WEST_SB_OUT_B1_valid(Tile_X00_Y02_SB_T4_WEST_SB_OUT_B1_valid),
		.clk(Tile_X00_Y01_clk_out),
		.clk_out(Tile_X00_Y02_clk_out),
		.clk_pass_through(Tile_X00_Y01_clk_pass_through_out_bot),
		.clk_pass_through_out_bot(Tile_X00_Y02_clk_pass_through_out_bot),
		.clk_pass_through_out_right(Tile_X00_Y02_clk_pass_through_out_right),
		.config_config_addr(Tile_X00_Y01_config_out_config_addr),
		.config_config_data(Tile_X00_Y01_config_out_config_data),
		.config_out_config_addr(Tile_X00_Y02_config_out_config_addr),
		.config_out_config_data(Tile_X00_Y02_config_out_config_data),
		.config_out_read(Tile_X00_Y02_config_out_read),
		.config_out_write(Tile_X00_Y02_config_out_write),
		.config_read(Tile_X00_Y01_config_out_read),
		.config_write(Tile_X00_Y01_config_out_write),
		.flush(Tile_X00_Y01_flush_out),
		.flush_out(Tile_X00_Y02_flush_out),
		.hi(Tile_X00_Y02_hi),
		.lo(Tile_X00_Y02_lo),
		.read_config_data(Tile_X00_Y02_read_config_data),
		.read_config_data_in(Tile_X00_Y01_read_config_data),
		.reset(Tile_X00_Y01_reset_out),
		.reset_out(Tile_X00_Y02_reset_out),
		.stall(Tile_X00_Y01_stall_out),
		.stall_out(Tile_X00_Y02_stall_out),
		.tile_id(Tile_X00_Y02_tile_id)
	);
	wire [15:0] Tile_X00_Y03_tile_id;
	assign Tile_X00_Y03_tile_id = {Tile_X00_Y03_lo[7], Tile_X00_Y03_lo[7], Tile_X00_Y03_lo[6], Tile_X00_Y03_lo[6], Tile_X00_Y03_lo[5], Tile_X00_Y03_lo[5], Tile_X00_Y03_lo[4], Tile_X00_Y03_lo[4], Tile_X00_Y03_lo[3], Tile_X00_Y03_lo[3], Tile_X00_Y03_lo[2], Tile_X00_Y03_lo[2], Tile_X00_Y03_lo[1], Tile_X00_Y03_lo[1], Tile_X00_Y03_hi[1], Tile_X00_Y03_hi[0]};
	Tile_PE Tile_X00_Y03(
		.SB_T0_EAST_SB_IN_B1(Tile_X01_Y03_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_EAST_SB_IN_B17(Tile_X01_Y03_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_EAST_SB_IN_B17_ready(Tile_X00_Y03_SB_T0_EAST_SB_IN_B17_ready),
		.SB_T0_EAST_SB_IN_B17_valid(Tile_X01_Y03_SB_T0_WEST_SB_OUT_B17_valid),
		.SB_T0_EAST_SB_IN_B1_ready(Tile_X00_Y03_SB_T0_EAST_SB_IN_B1_ready),
		.SB_T0_EAST_SB_IN_B1_valid(Tile_X01_Y03_SB_T0_WEST_SB_OUT_B1_valid),
		.SB_T0_EAST_SB_OUT_B1(Tile_X00_Y03_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_EAST_SB_OUT_B17(Tile_X00_Y03_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_EAST_SB_OUT_B17_ready(Tile_X01_Y03_SB_T0_WEST_SB_IN_B17_ready),
		.SB_T0_EAST_SB_OUT_B17_valid(Tile_X00_Y03_SB_T0_EAST_SB_OUT_B17_valid),
		.SB_T0_EAST_SB_OUT_B1_ready(Tile_X01_Y03_SB_T0_WEST_SB_IN_B1_ready),
		.SB_T0_EAST_SB_OUT_B1_valid(Tile_X00_Y03_SB_T0_EAST_SB_OUT_B1_valid),
		.SB_T0_NORTH_SB_IN_B1(Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_IN_B17(Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_IN_B17_ready(Tile_X00_Y03_SB_T0_NORTH_SB_IN_B17_ready),
		.SB_T0_NORTH_SB_IN_B17_valid(Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B17_valid),
		.SB_T0_NORTH_SB_IN_B1_ready(Tile_X00_Y03_SB_T0_NORTH_SB_IN_B1_ready),
		.SB_T0_NORTH_SB_IN_B1_valid(Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B1_valid),
		.SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_OUT_B17(Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_OUT_B17_ready(Tile_X00_Y02_SB_T0_SOUTH_SB_IN_B17_ready),
		.SB_T0_NORTH_SB_OUT_B17_valid(Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B17_valid),
		.SB_T0_NORTH_SB_OUT_B1_ready(Tile_X00_Y02_SB_T0_SOUTH_SB_IN_B1_ready),
		.SB_T0_NORTH_SB_OUT_B1_valid(Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B1_valid),
		.SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_IN_B17(Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_IN_B17_ready(Tile_X00_Y03_SB_T0_SOUTH_SB_IN_B17_ready),
		.SB_T0_SOUTH_SB_IN_B17_valid(Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B17_valid),
		.SB_T0_SOUTH_SB_IN_B1_ready(Tile_X00_Y03_SB_T0_SOUTH_SB_IN_B1_ready),
		.SB_T0_SOUTH_SB_IN_B1_valid(Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B1_valid),
		.SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_OUT_B17(Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_OUT_B17_ready(Tile_X00_Y04_SB_T0_NORTH_SB_IN_B17_ready),
		.SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B17_valid),
		.SB_T0_SOUTH_SB_OUT_B1_ready(Tile_X00_Y04_SB_T0_NORTH_SB_IN_B1_ready),
		.SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B1_valid),
		.SB_T0_WEST_SB_IN_B1(const_0_1_out),
		.SB_T0_WEST_SB_IN_B17(const_0_17_out),
		.SB_T0_WEST_SB_IN_B17_ready(Tile_X00_Y03_SB_T0_WEST_SB_IN_B17_ready),
		.SB_T0_WEST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T0_WEST_SB_IN_B1_ready(Tile_X00_Y03_SB_T0_WEST_SB_IN_B1_ready),
		.SB_T0_WEST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T0_WEST_SB_OUT_B1(Tile_X00_Y03_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_WEST_SB_OUT_B17(Tile_X00_Y03_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T0_WEST_SB_OUT_B17_valid(Tile_X00_Y03_SB_T0_WEST_SB_OUT_B17_valid),
		.SB_T0_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T0_WEST_SB_OUT_B1_valid(Tile_X00_Y03_SB_T0_WEST_SB_OUT_B1_valid),
		.SB_T1_EAST_SB_IN_B1(Tile_X01_Y03_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_EAST_SB_IN_B17(Tile_X01_Y03_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_EAST_SB_IN_B17_ready(Tile_X00_Y03_SB_T1_EAST_SB_IN_B17_ready),
		.SB_T1_EAST_SB_IN_B17_valid(Tile_X01_Y03_SB_T1_WEST_SB_OUT_B17_valid),
		.SB_T1_EAST_SB_IN_B1_ready(Tile_X00_Y03_SB_T1_EAST_SB_IN_B1_ready),
		.SB_T1_EAST_SB_IN_B1_valid(Tile_X01_Y03_SB_T1_WEST_SB_OUT_B1_valid),
		.SB_T1_EAST_SB_OUT_B1(Tile_X00_Y03_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_EAST_SB_OUT_B17(Tile_X00_Y03_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_EAST_SB_OUT_B17_ready(Tile_X01_Y03_SB_T1_WEST_SB_IN_B17_ready),
		.SB_T1_EAST_SB_OUT_B17_valid(Tile_X00_Y03_SB_T1_EAST_SB_OUT_B17_valid),
		.SB_T1_EAST_SB_OUT_B1_ready(Tile_X01_Y03_SB_T1_WEST_SB_IN_B1_ready),
		.SB_T1_EAST_SB_OUT_B1_valid(Tile_X00_Y03_SB_T1_EAST_SB_OUT_B1_valid),
		.SB_T1_NORTH_SB_IN_B1(Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_IN_B17(Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_IN_B17_ready(Tile_X00_Y03_SB_T1_NORTH_SB_IN_B17_ready),
		.SB_T1_NORTH_SB_IN_B17_valid(Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B17_valid),
		.SB_T1_NORTH_SB_IN_B1_ready(Tile_X00_Y03_SB_T1_NORTH_SB_IN_B1_ready),
		.SB_T1_NORTH_SB_IN_B1_valid(Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B1_valid),
		.SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_OUT_B17(Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_OUT_B17_ready(Tile_X00_Y02_SB_T1_SOUTH_SB_IN_B17_ready),
		.SB_T1_NORTH_SB_OUT_B17_valid(Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B17_valid),
		.SB_T1_NORTH_SB_OUT_B1_ready(Tile_X00_Y02_SB_T1_SOUTH_SB_IN_B1_ready),
		.SB_T1_NORTH_SB_OUT_B1_valid(Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B1_valid),
		.SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_IN_B17(Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_IN_B17_ready(Tile_X00_Y03_SB_T1_SOUTH_SB_IN_B17_ready),
		.SB_T1_SOUTH_SB_IN_B17_valid(Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B17_valid),
		.SB_T1_SOUTH_SB_IN_B1_ready(Tile_X00_Y03_SB_T1_SOUTH_SB_IN_B1_ready),
		.SB_T1_SOUTH_SB_IN_B1_valid(Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B1_valid),
		.SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_OUT_B17(Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_OUT_B17_ready(Tile_X00_Y04_SB_T1_NORTH_SB_IN_B17_ready),
		.SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B17_valid),
		.SB_T1_SOUTH_SB_OUT_B1_ready(Tile_X00_Y04_SB_T1_NORTH_SB_IN_B1_ready),
		.SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B1_valid),
		.SB_T1_WEST_SB_IN_B1(const_0_1_out),
		.SB_T1_WEST_SB_IN_B17(const_0_17_out),
		.SB_T1_WEST_SB_IN_B17_ready(Tile_X00_Y03_SB_T1_WEST_SB_IN_B17_ready),
		.SB_T1_WEST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T1_WEST_SB_IN_B1_ready(Tile_X00_Y03_SB_T1_WEST_SB_IN_B1_ready),
		.SB_T1_WEST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T1_WEST_SB_OUT_B1(Tile_X00_Y03_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_WEST_SB_OUT_B17(Tile_X00_Y03_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T1_WEST_SB_OUT_B17_valid(Tile_X00_Y03_SB_T1_WEST_SB_OUT_B17_valid),
		.SB_T1_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T1_WEST_SB_OUT_B1_valid(Tile_X00_Y03_SB_T1_WEST_SB_OUT_B1_valid),
		.SB_T2_EAST_SB_IN_B1(Tile_X01_Y03_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_EAST_SB_IN_B17(Tile_X01_Y03_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_EAST_SB_IN_B17_ready(Tile_X00_Y03_SB_T2_EAST_SB_IN_B17_ready),
		.SB_T2_EAST_SB_IN_B17_valid(Tile_X01_Y03_SB_T2_WEST_SB_OUT_B17_valid),
		.SB_T2_EAST_SB_IN_B1_ready(Tile_X00_Y03_SB_T2_EAST_SB_IN_B1_ready),
		.SB_T2_EAST_SB_IN_B1_valid(Tile_X01_Y03_SB_T2_WEST_SB_OUT_B1_valid),
		.SB_T2_EAST_SB_OUT_B1(Tile_X00_Y03_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_EAST_SB_OUT_B17(Tile_X00_Y03_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_EAST_SB_OUT_B17_ready(Tile_X01_Y03_SB_T2_WEST_SB_IN_B17_ready),
		.SB_T2_EAST_SB_OUT_B17_valid(Tile_X00_Y03_SB_T2_EAST_SB_OUT_B17_valid),
		.SB_T2_EAST_SB_OUT_B1_ready(Tile_X01_Y03_SB_T2_WEST_SB_IN_B1_ready),
		.SB_T2_EAST_SB_OUT_B1_valid(Tile_X00_Y03_SB_T2_EAST_SB_OUT_B1_valid),
		.SB_T2_NORTH_SB_IN_B1(Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_IN_B17(Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_IN_B17_ready(Tile_X00_Y03_SB_T2_NORTH_SB_IN_B17_ready),
		.SB_T2_NORTH_SB_IN_B17_valid(Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B17_valid),
		.SB_T2_NORTH_SB_IN_B1_ready(Tile_X00_Y03_SB_T2_NORTH_SB_IN_B1_ready),
		.SB_T2_NORTH_SB_IN_B1_valid(Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B1_valid),
		.SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_OUT_B17(Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_OUT_B17_ready(Tile_X00_Y02_SB_T2_SOUTH_SB_IN_B17_ready),
		.SB_T2_NORTH_SB_OUT_B17_valid(Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B17_valid),
		.SB_T2_NORTH_SB_OUT_B1_ready(Tile_X00_Y02_SB_T2_SOUTH_SB_IN_B1_ready),
		.SB_T2_NORTH_SB_OUT_B1_valid(Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B1_valid),
		.SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_IN_B17(Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_IN_B17_ready(Tile_X00_Y03_SB_T2_SOUTH_SB_IN_B17_ready),
		.SB_T2_SOUTH_SB_IN_B17_valid(Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B17_valid),
		.SB_T2_SOUTH_SB_IN_B1_ready(Tile_X00_Y03_SB_T2_SOUTH_SB_IN_B1_ready),
		.SB_T2_SOUTH_SB_IN_B1_valid(Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B1_valid),
		.SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_OUT_B17(Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_OUT_B17_ready(Tile_X00_Y04_SB_T2_NORTH_SB_IN_B17_ready),
		.SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B17_valid),
		.SB_T2_SOUTH_SB_OUT_B1_ready(Tile_X00_Y04_SB_T2_NORTH_SB_IN_B1_ready),
		.SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B1_valid),
		.SB_T2_WEST_SB_IN_B1(const_0_1_out),
		.SB_T2_WEST_SB_IN_B17(const_0_17_out),
		.SB_T2_WEST_SB_IN_B17_ready(Tile_X00_Y03_SB_T2_WEST_SB_IN_B17_ready),
		.SB_T2_WEST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T2_WEST_SB_IN_B1_ready(Tile_X00_Y03_SB_T2_WEST_SB_IN_B1_ready),
		.SB_T2_WEST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T2_WEST_SB_OUT_B1(Tile_X00_Y03_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_WEST_SB_OUT_B17(Tile_X00_Y03_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T2_WEST_SB_OUT_B17_valid(Tile_X00_Y03_SB_T2_WEST_SB_OUT_B17_valid),
		.SB_T2_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T2_WEST_SB_OUT_B1_valid(Tile_X00_Y03_SB_T2_WEST_SB_OUT_B1_valid),
		.SB_T3_EAST_SB_IN_B1(Tile_X01_Y03_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_EAST_SB_IN_B17(Tile_X01_Y03_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_EAST_SB_IN_B17_ready(Tile_X00_Y03_SB_T3_EAST_SB_IN_B17_ready),
		.SB_T3_EAST_SB_IN_B17_valid(Tile_X01_Y03_SB_T3_WEST_SB_OUT_B17_valid),
		.SB_T3_EAST_SB_IN_B1_ready(Tile_X00_Y03_SB_T3_EAST_SB_IN_B1_ready),
		.SB_T3_EAST_SB_IN_B1_valid(Tile_X01_Y03_SB_T3_WEST_SB_OUT_B1_valid),
		.SB_T3_EAST_SB_OUT_B1(Tile_X00_Y03_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_EAST_SB_OUT_B17(Tile_X00_Y03_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_EAST_SB_OUT_B17_ready(Tile_X01_Y03_SB_T3_WEST_SB_IN_B17_ready),
		.SB_T3_EAST_SB_OUT_B17_valid(Tile_X00_Y03_SB_T3_EAST_SB_OUT_B17_valid),
		.SB_T3_EAST_SB_OUT_B1_ready(Tile_X01_Y03_SB_T3_WEST_SB_IN_B1_ready),
		.SB_T3_EAST_SB_OUT_B1_valid(Tile_X00_Y03_SB_T3_EAST_SB_OUT_B1_valid),
		.SB_T3_NORTH_SB_IN_B1(Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_IN_B17(Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_IN_B17_ready(Tile_X00_Y03_SB_T3_NORTH_SB_IN_B17_ready),
		.SB_T3_NORTH_SB_IN_B17_valid(Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B17_valid),
		.SB_T3_NORTH_SB_IN_B1_ready(Tile_X00_Y03_SB_T3_NORTH_SB_IN_B1_ready),
		.SB_T3_NORTH_SB_IN_B1_valid(Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B1_valid),
		.SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_OUT_B17(Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_OUT_B17_ready(Tile_X00_Y02_SB_T3_SOUTH_SB_IN_B17_ready),
		.SB_T3_NORTH_SB_OUT_B17_valid(Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B17_valid),
		.SB_T3_NORTH_SB_OUT_B1_ready(Tile_X00_Y02_SB_T3_SOUTH_SB_IN_B1_ready),
		.SB_T3_NORTH_SB_OUT_B1_valid(Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B1_valid),
		.SB_T3_SOUTH_SB_IN_B1(Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_IN_B17(Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_IN_B17_ready(Tile_X00_Y03_SB_T3_SOUTH_SB_IN_B17_ready),
		.SB_T3_SOUTH_SB_IN_B17_valid(Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B17_valid),
		.SB_T3_SOUTH_SB_IN_B1_ready(Tile_X00_Y03_SB_T3_SOUTH_SB_IN_B1_ready),
		.SB_T3_SOUTH_SB_IN_B1_valid(Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B1_valid),
		.SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_OUT_B17(Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_OUT_B17_ready(Tile_X00_Y04_SB_T3_NORTH_SB_IN_B17_ready),
		.SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B17_valid),
		.SB_T3_SOUTH_SB_OUT_B1_ready(Tile_X00_Y04_SB_T3_NORTH_SB_IN_B1_ready),
		.SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B1_valid),
		.SB_T3_WEST_SB_IN_B1(const_0_1_out),
		.SB_T3_WEST_SB_IN_B17(const_0_17_out),
		.SB_T3_WEST_SB_IN_B17_ready(Tile_X00_Y03_SB_T3_WEST_SB_IN_B17_ready),
		.SB_T3_WEST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T3_WEST_SB_IN_B1_ready(Tile_X00_Y03_SB_T3_WEST_SB_IN_B1_ready),
		.SB_T3_WEST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T3_WEST_SB_OUT_B1(Tile_X00_Y03_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_WEST_SB_OUT_B17(Tile_X00_Y03_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T3_WEST_SB_OUT_B17_valid(Tile_X00_Y03_SB_T3_WEST_SB_OUT_B17_valid),
		.SB_T3_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T3_WEST_SB_OUT_B1_valid(Tile_X00_Y03_SB_T3_WEST_SB_OUT_B1_valid),
		.SB_T4_EAST_SB_IN_B1(Tile_X01_Y03_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_EAST_SB_IN_B17(Tile_X01_Y03_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_EAST_SB_IN_B17_ready(Tile_X00_Y03_SB_T4_EAST_SB_IN_B17_ready),
		.SB_T4_EAST_SB_IN_B17_valid(Tile_X01_Y03_SB_T4_WEST_SB_OUT_B17_valid),
		.SB_T4_EAST_SB_IN_B1_ready(Tile_X00_Y03_SB_T4_EAST_SB_IN_B1_ready),
		.SB_T4_EAST_SB_IN_B1_valid(Tile_X01_Y03_SB_T4_WEST_SB_OUT_B1_valid),
		.SB_T4_EAST_SB_OUT_B1(Tile_X00_Y03_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_EAST_SB_OUT_B17(Tile_X00_Y03_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_EAST_SB_OUT_B17_ready(Tile_X01_Y03_SB_T4_WEST_SB_IN_B17_ready),
		.SB_T4_EAST_SB_OUT_B17_valid(Tile_X00_Y03_SB_T4_EAST_SB_OUT_B17_valid),
		.SB_T4_EAST_SB_OUT_B1_ready(Tile_X01_Y03_SB_T4_WEST_SB_IN_B1_ready),
		.SB_T4_EAST_SB_OUT_B1_valid(Tile_X00_Y03_SB_T4_EAST_SB_OUT_B1_valid),
		.SB_T4_NORTH_SB_IN_B1(Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_IN_B17(Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_IN_B17_ready(Tile_X00_Y03_SB_T4_NORTH_SB_IN_B17_ready),
		.SB_T4_NORTH_SB_IN_B17_valid(Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B17_valid),
		.SB_T4_NORTH_SB_IN_B1_ready(Tile_X00_Y03_SB_T4_NORTH_SB_IN_B1_ready),
		.SB_T4_NORTH_SB_IN_B1_valid(Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B1_valid),
		.SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_OUT_B17(Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_OUT_B17_ready(Tile_X00_Y02_SB_T4_SOUTH_SB_IN_B17_ready),
		.SB_T4_NORTH_SB_OUT_B17_valid(Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B17_valid),
		.SB_T4_NORTH_SB_OUT_B1_ready(Tile_X00_Y02_SB_T4_SOUTH_SB_IN_B1_ready),
		.SB_T4_NORTH_SB_OUT_B1_valid(Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B1_valid),
		.SB_T4_SOUTH_SB_IN_B1(Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_IN_B17(Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_IN_B17_ready(Tile_X00_Y03_SB_T4_SOUTH_SB_IN_B17_ready),
		.SB_T4_SOUTH_SB_IN_B17_valid(Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B17_valid),
		.SB_T4_SOUTH_SB_IN_B1_ready(Tile_X00_Y03_SB_T4_SOUTH_SB_IN_B1_ready),
		.SB_T4_SOUTH_SB_IN_B1_valid(Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B1_valid),
		.SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_OUT_B17(Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_OUT_B17_ready(Tile_X00_Y04_SB_T4_NORTH_SB_IN_B17_ready),
		.SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B17_valid),
		.SB_T4_SOUTH_SB_OUT_B1_ready(Tile_X00_Y04_SB_T4_NORTH_SB_IN_B1_ready),
		.SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B1_valid),
		.SB_T4_WEST_SB_IN_B1(const_0_1_out),
		.SB_T4_WEST_SB_IN_B17(const_0_17_out),
		.SB_T4_WEST_SB_IN_B17_ready(Tile_X00_Y03_SB_T4_WEST_SB_IN_B17_ready),
		.SB_T4_WEST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T4_WEST_SB_IN_B1_ready(Tile_X00_Y03_SB_T4_WEST_SB_IN_B1_ready),
		.SB_T4_WEST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T4_WEST_SB_OUT_B1(Tile_X00_Y03_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_WEST_SB_OUT_B17(Tile_X00_Y03_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T4_WEST_SB_OUT_B17_valid(Tile_X00_Y03_SB_T4_WEST_SB_OUT_B17_valid),
		.SB_T4_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T4_WEST_SB_OUT_B1_valid(Tile_X00_Y03_SB_T4_WEST_SB_OUT_B1_valid),
		.clk(Tile_X00_Y02_clk_out),
		.clk_out(Tile_X00_Y03_clk_out),
		.clk_pass_through(Tile_X00_Y02_clk_pass_through_out_bot),
		.clk_pass_through_out_bot(Tile_X00_Y03_clk_pass_through_out_bot),
		.clk_pass_through_out_right(Tile_X00_Y03_clk_pass_through_out_right),
		.config_config_addr(Tile_X00_Y02_config_out_config_addr),
		.config_config_data(Tile_X00_Y02_config_out_config_data),
		.config_out_config_addr(Tile_X00_Y03_config_out_config_addr),
		.config_out_config_data(Tile_X00_Y03_config_out_config_data),
		.config_out_read(Tile_X00_Y03_config_out_read),
		.config_out_write(Tile_X00_Y03_config_out_write),
		.config_read(Tile_X00_Y02_config_out_read),
		.config_write(Tile_X00_Y02_config_out_write),
		.flush(Tile_X00_Y02_flush_out),
		.flush_out(Tile_X00_Y03_flush_out),
		.hi(Tile_X00_Y03_hi),
		.lo(Tile_X00_Y03_lo),
		.read_config_data(Tile_X00_Y03_read_config_data),
		.read_config_data_in(Tile_X00_Y02_read_config_data),
		.reset(Tile_X00_Y02_reset_out),
		.reset_out(Tile_X00_Y03_reset_out),
		.stall(Tile_X00_Y02_stall_out),
		.stall_out(Tile_X00_Y03_stall_out),
		.tile_id(Tile_X00_Y03_tile_id)
	);
	wire [15:0] Tile_X00_Y04_tile_id;
	assign Tile_X00_Y04_tile_id = {Tile_X00_Y04_lo[7], Tile_X00_Y04_lo[7], Tile_X00_Y04_lo[6], Tile_X00_Y04_lo[6], Tile_X00_Y04_lo[5], Tile_X00_Y04_lo[5], Tile_X00_Y04_lo[4], Tile_X00_Y04_lo[4], Tile_X00_Y04_lo[3], Tile_X00_Y04_lo[3], Tile_X00_Y04_lo[2], Tile_X00_Y04_lo[2], Tile_X00_Y04_lo[1], Tile_X00_Y04_hi[1], Tile_X00_Y04_lo[0], Tile_X00_Y04_lo[0]};
	Tile_PE Tile_X00_Y04(
		.SB_T0_EAST_SB_IN_B1(Tile_X01_Y04_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_EAST_SB_IN_B17(Tile_X01_Y04_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_EAST_SB_IN_B17_ready(Tile_X00_Y04_SB_T0_EAST_SB_IN_B17_ready),
		.SB_T0_EAST_SB_IN_B17_valid(Tile_X01_Y04_SB_T0_WEST_SB_OUT_B17_valid),
		.SB_T0_EAST_SB_IN_B1_ready(Tile_X00_Y04_SB_T0_EAST_SB_IN_B1_ready),
		.SB_T0_EAST_SB_IN_B1_valid(Tile_X01_Y04_SB_T0_WEST_SB_OUT_B1_valid),
		.SB_T0_EAST_SB_OUT_B1(Tile_X00_Y04_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_EAST_SB_OUT_B17(Tile_X00_Y04_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_EAST_SB_OUT_B17_ready(Tile_X01_Y04_SB_T0_WEST_SB_IN_B17_ready),
		.SB_T0_EAST_SB_OUT_B17_valid(Tile_X00_Y04_SB_T0_EAST_SB_OUT_B17_valid),
		.SB_T0_EAST_SB_OUT_B1_ready(Tile_X01_Y04_SB_T0_WEST_SB_IN_B1_ready),
		.SB_T0_EAST_SB_OUT_B1_valid(Tile_X00_Y04_SB_T0_EAST_SB_OUT_B1_valid),
		.SB_T0_NORTH_SB_IN_B1(Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_IN_B17(Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_IN_B17_ready(Tile_X00_Y04_SB_T0_NORTH_SB_IN_B17_ready),
		.SB_T0_NORTH_SB_IN_B17_valid(Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B17_valid),
		.SB_T0_NORTH_SB_IN_B1_ready(Tile_X00_Y04_SB_T0_NORTH_SB_IN_B1_ready),
		.SB_T0_NORTH_SB_IN_B1_valid(Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B1_valid),
		.SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_OUT_B17(Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_OUT_B17_ready(Tile_X00_Y03_SB_T0_SOUTH_SB_IN_B17_ready),
		.SB_T0_NORTH_SB_OUT_B17_valid(Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B17_valid),
		.SB_T0_NORTH_SB_OUT_B1_ready(Tile_X00_Y03_SB_T0_SOUTH_SB_IN_B1_ready),
		.SB_T0_NORTH_SB_OUT_B1_valid(Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B1_valid),
		.SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
		.SB_T0_SOUTH_SB_IN_B17(const_0_17_out),
		.SB_T0_SOUTH_SB_IN_B17_ready(Tile_X00_Y04_SB_T0_SOUTH_SB_IN_B17_ready),
		.SB_T0_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T0_SOUTH_SB_IN_B1_ready(Tile_X00_Y04_SB_T0_SOUTH_SB_IN_B1_ready),
		.SB_T0_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_OUT_B17(Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B17_valid),
		.SB_T0_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B1_valid),
		.SB_T0_WEST_SB_IN_B1(const_0_1_out),
		.SB_T0_WEST_SB_IN_B17(const_0_17_out),
		.SB_T0_WEST_SB_IN_B17_ready(Tile_X00_Y04_SB_T0_WEST_SB_IN_B17_ready),
		.SB_T0_WEST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T0_WEST_SB_IN_B1_ready(Tile_X00_Y04_SB_T0_WEST_SB_IN_B1_ready),
		.SB_T0_WEST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T0_WEST_SB_OUT_B1(Tile_X00_Y04_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_WEST_SB_OUT_B17(Tile_X00_Y04_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T0_WEST_SB_OUT_B17_valid(Tile_X00_Y04_SB_T0_WEST_SB_OUT_B17_valid),
		.SB_T0_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T0_WEST_SB_OUT_B1_valid(Tile_X00_Y04_SB_T0_WEST_SB_OUT_B1_valid),
		.SB_T1_EAST_SB_IN_B1(Tile_X01_Y04_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_EAST_SB_IN_B17(Tile_X01_Y04_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_EAST_SB_IN_B17_ready(Tile_X00_Y04_SB_T1_EAST_SB_IN_B17_ready),
		.SB_T1_EAST_SB_IN_B17_valid(Tile_X01_Y04_SB_T1_WEST_SB_OUT_B17_valid),
		.SB_T1_EAST_SB_IN_B1_ready(Tile_X00_Y04_SB_T1_EAST_SB_IN_B1_ready),
		.SB_T1_EAST_SB_IN_B1_valid(Tile_X01_Y04_SB_T1_WEST_SB_OUT_B1_valid),
		.SB_T1_EAST_SB_OUT_B1(Tile_X00_Y04_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_EAST_SB_OUT_B17(Tile_X00_Y04_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_EAST_SB_OUT_B17_ready(Tile_X01_Y04_SB_T1_WEST_SB_IN_B17_ready),
		.SB_T1_EAST_SB_OUT_B17_valid(Tile_X00_Y04_SB_T1_EAST_SB_OUT_B17_valid),
		.SB_T1_EAST_SB_OUT_B1_ready(Tile_X01_Y04_SB_T1_WEST_SB_IN_B1_ready),
		.SB_T1_EAST_SB_OUT_B1_valid(Tile_X00_Y04_SB_T1_EAST_SB_OUT_B1_valid),
		.SB_T1_NORTH_SB_IN_B1(Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_IN_B17(Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_IN_B17_ready(Tile_X00_Y04_SB_T1_NORTH_SB_IN_B17_ready),
		.SB_T1_NORTH_SB_IN_B17_valid(Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B17_valid),
		.SB_T1_NORTH_SB_IN_B1_ready(Tile_X00_Y04_SB_T1_NORTH_SB_IN_B1_ready),
		.SB_T1_NORTH_SB_IN_B1_valid(Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B1_valid),
		.SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_OUT_B17(Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_OUT_B17_ready(Tile_X00_Y03_SB_T1_SOUTH_SB_IN_B17_ready),
		.SB_T1_NORTH_SB_OUT_B17_valid(Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B17_valid),
		.SB_T1_NORTH_SB_OUT_B1_ready(Tile_X00_Y03_SB_T1_SOUTH_SB_IN_B1_ready),
		.SB_T1_NORTH_SB_OUT_B1_valid(Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B1_valid),
		.SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
		.SB_T1_SOUTH_SB_IN_B17(const_0_17_out),
		.SB_T1_SOUTH_SB_IN_B17_ready(Tile_X00_Y04_SB_T1_SOUTH_SB_IN_B17_ready),
		.SB_T1_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T1_SOUTH_SB_IN_B1_ready(Tile_X00_Y04_SB_T1_SOUTH_SB_IN_B1_ready),
		.SB_T1_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_OUT_B17(Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B17_valid),
		.SB_T1_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B1_valid),
		.SB_T1_WEST_SB_IN_B1(const_0_1_out),
		.SB_T1_WEST_SB_IN_B17(const_0_17_out),
		.SB_T1_WEST_SB_IN_B17_ready(Tile_X00_Y04_SB_T1_WEST_SB_IN_B17_ready),
		.SB_T1_WEST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T1_WEST_SB_IN_B1_ready(Tile_X00_Y04_SB_T1_WEST_SB_IN_B1_ready),
		.SB_T1_WEST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T1_WEST_SB_OUT_B1(Tile_X00_Y04_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_WEST_SB_OUT_B17(Tile_X00_Y04_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T1_WEST_SB_OUT_B17_valid(Tile_X00_Y04_SB_T1_WEST_SB_OUT_B17_valid),
		.SB_T1_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T1_WEST_SB_OUT_B1_valid(Tile_X00_Y04_SB_T1_WEST_SB_OUT_B1_valid),
		.SB_T2_EAST_SB_IN_B1(Tile_X01_Y04_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_EAST_SB_IN_B17(Tile_X01_Y04_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_EAST_SB_IN_B17_ready(Tile_X00_Y04_SB_T2_EAST_SB_IN_B17_ready),
		.SB_T2_EAST_SB_IN_B17_valid(Tile_X01_Y04_SB_T2_WEST_SB_OUT_B17_valid),
		.SB_T2_EAST_SB_IN_B1_ready(Tile_X00_Y04_SB_T2_EAST_SB_IN_B1_ready),
		.SB_T2_EAST_SB_IN_B1_valid(Tile_X01_Y04_SB_T2_WEST_SB_OUT_B1_valid),
		.SB_T2_EAST_SB_OUT_B1(Tile_X00_Y04_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_EAST_SB_OUT_B17(Tile_X00_Y04_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_EAST_SB_OUT_B17_ready(Tile_X01_Y04_SB_T2_WEST_SB_IN_B17_ready),
		.SB_T2_EAST_SB_OUT_B17_valid(Tile_X00_Y04_SB_T2_EAST_SB_OUT_B17_valid),
		.SB_T2_EAST_SB_OUT_B1_ready(Tile_X01_Y04_SB_T2_WEST_SB_IN_B1_ready),
		.SB_T2_EAST_SB_OUT_B1_valid(Tile_X00_Y04_SB_T2_EAST_SB_OUT_B1_valid),
		.SB_T2_NORTH_SB_IN_B1(Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_IN_B17(Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_IN_B17_ready(Tile_X00_Y04_SB_T2_NORTH_SB_IN_B17_ready),
		.SB_T2_NORTH_SB_IN_B17_valid(Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B17_valid),
		.SB_T2_NORTH_SB_IN_B1_ready(Tile_X00_Y04_SB_T2_NORTH_SB_IN_B1_ready),
		.SB_T2_NORTH_SB_IN_B1_valid(Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B1_valid),
		.SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_OUT_B17(Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_OUT_B17_ready(Tile_X00_Y03_SB_T2_SOUTH_SB_IN_B17_ready),
		.SB_T2_NORTH_SB_OUT_B17_valid(Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B17_valid),
		.SB_T2_NORTH_SB_OUT_B1_ready(Tile_X00_Y03_SB_T2_SOUTH_SB_IN_B1_ready),
		.SB_T2_NORTH_SB_OUT_B1_valid(Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B1_valid),
		.SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
		.SB_T2_SOUTH_SB_IN_B17(const_0_17_out),
		.SB_T2_SOUTH_SB_IN_B17_ready(Tile_X00_Y04_SB_T2_SOUTH_SB_IN_B17_ready),
		.SB_T2_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T2_SOUTH_SB_IN_B1_ready(Tile_X00_Y04_SB_T2_SOUTH_SB_IN_B1_ready),
		.SB_T2_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_OUT_B17(Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B17_valid),
		.SB_T2_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B1_valid),
		.SB_T2_WEST_SB_IN_B1(const_0_1_out),
		.SB_T2_WEST_SB_IN_B17(const_0_17_out),
		.SB_T2_WEST_SB_IN_B17_ready(Tile_X00_Y04_SB_T2_WEST_SB_IN_B17_ready),
		.SB_T2_WEST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T2_WEST_SB_IN_B1_ready(Tile_X00_Y04_SB_T2_WEST_SB_IN_B1_ready),
		.SB_T2_WEST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T2_WEST_SB_OUT_B1(Tile_X00_Y04_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_WEST_SB_OUT_B17(Tile_X00_Y04_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T2_WEST_SB_OUT_B17_valid(Tile_X00_Y04_SB_T2_WEST_SB_OUT_B17_valid),
		.SB_T2_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T2_WEST_SB_OUT_B1_valid(Tile_X00_Y04_SB_T2_WEST_SB_OUT_B1_valid),
		.SB_T3_EAST_SB_IN_B1(Tile_X01_Y04_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_EAST_SB_IN_B17(Tile_X01_Y04_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_EAST_SB_IN_B17_ready(Tile_X00_Y04_SB_T3_EAST_SB_IN_B17_ready),
		.SB_T3_EAST_SB_IN_B17_valid(Tile_X01_Y04_SB_T3_WEST_SB_OUT_B17_valid),
		.SB_T3_EAST_SB_IN_B1_ready(Tile_X00_Y04_SB_T3_EAST_SB_IN_B1_ready),
		.SB_T3_EAST_SB_IN_B1_valid(Tile_X01_Y04_SB_T3_WEST_SB_OUT_B1_valid),
		.SB_T3_EAST_SB_OUT_B1(Tile_X00_Y04_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_EAST_SB_OUT_B17(Tile_X00_Y04_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_EAST_SB_OUT_B17_ready(Tile_X01_Y04_SB_T3_WEST_SB_IN_B17_ready),
		.SB_T3_EAST_SB_OUT_B17_valid(Tile_X00_Y04_SB_T3_EAST_SB_OUT_B17_valid),
		.SB_T3_EAST_SB_OUT_B1_ready(Tile_X01_Y04_SB_T3_WEST_SB_IN_B1_ready),
		.SB_T3_EAST_SB_OUT_B1_valid(Tile_X00_Y04_SB_T3_EAST_SB_OUT_B1_valid),
		.SB_T3_NORTH_SB_IN_B1(Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_IN_B17(Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_IN_B17_ready(Tile_X00_Y04_SB_T3_NORTH_SB_IN_B17_ready),
		.SB_T3_NORTH_SB_IN_B17_valid(Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B17_valid),
		.SB_T3_NORTH_SB_IN_B1_ready(Tile_X00_Y04_SB_T3_NORTH_SB_IN_B1_ready),
		.SB_T3_NORTH_SB_IN_B1_valid(Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B1_valid),
		.SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_OUT_B17(Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_OUT_B17_ready(Tile_X00_Y03_SB_T3_SOUTH_SB_IN_B17_ready),
		.SB_T3_NORTH_SB_OUT_B17_valid(Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B17_valid),
		.SB_T3_NORTH_SB_OUT_B1_ready(Tile_X00_Y03_SB_T3_SOUTH_SB_IN_B1_ready),
		.SB_T3_NORTH_SB_OUT_B1_valid(Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B1_valid),
		.SB_T3_SOUTH_SB_IN_B1(const_0_1_out),
		.SB_T3_SOUTH_SB_IN_B17(const_0_17_out),
		.SB_T3_SOUTH_SB_IN_B17_ready(Tile_X00_Y04_SB_T3_SOUTH_SB_IN_B17_ready),
		.SB_T3_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T3_SOUTH_SB_IN_B1_ready(Tile_X00_Y04_SB_T3_SOUTH_SB_IN_B1_ready),
		.SB_T3_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y04_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_OUT_B17(Tile_X00_Y04_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X00_Y04_SB_T3_SOUTH_SB_OUT_B17_valid),
		.SB_T3_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X00_Y04_SB_T3_SOUTH_SB_OUT_B1_valid),
		.SB_T3_WEST_SB_IN_B1(const_0_1_out),
		.SB_T3_WEST_SB_IN_B17(const_0_17_out),
		.SB_T3_WEST_SB_IN_B17_ready(Tile_X00_Y04_SB_T3_WEST_SB_IN_B17_ready),
		.SB_T3_WEST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T3_WEST_SB_IN_B1_ready(Tile_X00_Y04_SB_T3_WEST_SB_IN_B1_ready),
		.SB_T3_WEST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T3_WEST_SB_OUT_B1(Tile_X00_Y04_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_WEST_SB_OUT_B17(Tile_X00_Y04_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T3_WEST_SB_OUT_B17_valid(Tile_X00_Y04_SB_T3_WEST_SB_OUT_B17_valid),
		.SB_T3_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T3_WEST_SB_OUT_B1_valid(Tile_X00_Y04_SB_T3_WEST_SB_OUT_B1_valid),
		.SB_T4_EAST_SB_IN_B1(Tile_X01_Y04_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_EAST_SB_IN_B17(Tile_X01_Y04_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_EAST_SB_IN_B17_ready(Tile_X00_Y04_SB_T4_EAST_SB_IN_B17_ready),
		.SB_T4_EAST_SB_IN_B17_valid(Tile_X01_Y04_SB_T4_WEST_SB_OUT_B17_valid),
		.SB_T4_EAST_SB_IN_B1_ready(Tile_X00_Y04_SB_T4_EAST_SB_IN_B1_ready),
		.SB_T4_EAST_SB_IN_B1_valid(Tile_X01_Y04_SB_T4_WEST_SB_OUT_B1_valid),
		.SB_T4_EAST_SB_OUT_B1(Tile_X00_Y04_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_EAST_SB_OUT_B17(Tile_X00_Y04_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_EAST_SB_OUT_B17_ready(Tile_X01_Y04_SB_T4_WEST_SB_IN_B17_ready),
		.SB_T4_EAST_SB_OUT_B17_valid(Tile_X00_Y04_SB_T4_EAST_SB_OUT_B17_valid),
		.SB_T4_EAST_SB_OUT_B1_ready(Tile_X01_Y04_SB_T4_WEST_SB_IN_B1_ready),
		.SB_T4_EAST_SB_OUT_B1_valid(Tile_X00_Y04_SB_T4_EAST_SB_OUT_B1_valid),
		.SB_T4_NORTH_SB_IN_B1(Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_IN_B17(Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_IN_B17_ready(Tile_X00_Y04_SB_T4_NORTH_SB_IN_B17_ready),
		.SB_T4_NORTH_SB_IN_B17_valid(Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B17_valid),
		.SB_T4_NORTH_SB_IN_B1_ready(Tile_X00_Y04_SB_T4_NORTH_SB_IN_B1_ready),
		.SB_T4_NORTH_SB_IN_B1_valid(Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B1_valid),
		.SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_OUT_B17(Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_OUT_B17_ready(Tile_X00_Y03_SB_T4_SOUTH_SB_IN_B17_ready),
		.SB_T4_NORTH_SB_OUT_B17_valid(Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B17_valid),
		.SB_T4_NORTH_SB_OUT_B1_ready(Tile_X00_Y03_SB_T4_SOUTH_SB_IN_B1_ready),
		.SB_T4_NORTH_SB_OUT_B1_valid(Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B1_valid),
		.SB_T4_SOUTH_SB_IN_B1(const_0_1_out),
		.SB_T4_SOUTH_SB_IN_B17(const_0_17_out),
		.SB_T4_SOUTH_SB_IN_B17_ready(Tile_X00_Y04_SB_T4_SOUTH_SB_IN_B17_ready),
		.SB_T4_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T4_SOUTH_SB_IN_B1_ready(Tile_X00_Y04_SB_T4_SOUTH_SB_IN_B1_ready),
		.SB_T4_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y04_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_OUT_B17(Tile_X00_Y04_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X00_Y04_SB_T4_SOUTH_SB_OUT_B17_valid),
		.SB_T4_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X00_Y04_SB_T4_SOUTH_SB_OUT_B1_valid),
		.SB_T4_WEST_SB_IN_B1(const_0_1_out),
		.SB_T4_WEST_SB_IN_B17(const_0_17_out),
		.SB_T4_WEST_SB_IN_B17_ready(Tile_X00_Y04_SB_T4_WEST_SB_IN_B17_ready),
		.SB_T4_WEST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T4_WEST_SB_IN_B1_ready(Tile_X00_Y04_SB_T4_WEST_SB_IN_B1_ready),
		.SB_T4_WEST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T4_WEST_SB_OUT_B1(Tile_X00_Y04_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_WEST_SB_OUT_B17(Tile_X00_Y04_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T4_WEST_SB_OUT_B17_valid(Tile_X00_Y04_SB_T4_WEST_SB_OUT_B17_valid),
		.SB_T4_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T4_WEST_SB_OUT_B1_valid(Tile_X00_Y04_SB_T4_WEST_SB_OUT_B1_valid),
		.clk(Tile_X00_Y03_clk_out),
		.clk_out(Tile_X00_Y04_clk_out),
		.clk_pass_through(Tile_X00_Y03_clk_pass_through_out_bot),
		.clk_pass_through_out_bot(Tile_X00_Y04_clk_pass_through_out_bot),
		.clk_pass_through_out_right(Tile_X00_Y04_clk_pass_through_out_right),
		.config_config_addr(Tile_X00_Y03_config_out_config_addr),
		.config_config_data(Tile_X00_Y03_config_out_config_data),
		.config_out_config_addr(Tile_X00_Y04_config_out_config_addr),
		.config_out_config_data(Tile_X00_Y04_config_out_config_data),
		.config_out_read(Tile_X00_Y04_config_out_read),
		.config_out_write(Tile_X00_Y04_config_out_write),
		.config_read(Tile_X00_Y03_config_out_read),
		.config_write(Tile_X00_Y03_config_out_write),
		.flush(Tile_X00_Y03_flush_out),
		.flush_out(Tile_X00_Y04_flush_out),
		.hi(Tile_X00_Y04_hi),
		.lo(Tile_X00_Y04_lo),
		.read_config_data(Tile_X00_Y04_read_config_data),
		.read_config_data_in(Tile_X00_Y03_read_config_data),
		.reset(Tile_X00_Y03_reset_out),
		.reset_out(Tile_X00_Y04_reset_out),
		.stall(Tile_X00_Y03_stall_out),
		.stall_out(Tile_X00_Y04_stall_out),
		.tile_id(Tile_X00_Y04_tile_id)
	);
	wire [31:0] Tile_X01_Y00_config_config_addr;
	assign Tile_X01_Y00_config_config_addr = {PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[31], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[30], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[29], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[28], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[27], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[26], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[25], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[24], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[23], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[22], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[21], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[20], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[19], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[18], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[17], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[16], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[15], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[14], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[13], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[12], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[11], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[10], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[9], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[8], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[7], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[6], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[5], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[4], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[3], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[2], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[1], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[0]};
	wire [31:0] Tile_X01_Y00_config_config_data;
	assign Tile_X01_Y00_config_config_data = {PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[63], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[62], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[61], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[60], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[59], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[58], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[57], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[56], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[55], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[54], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[53], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[52], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[51], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[50], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[49], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[48], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[47], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[46], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[45], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[44], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[43], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[42], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[41], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[40], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[39], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[38], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[37], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[36], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[35], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[34], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[33], PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[32]};
	wire [4:0] Tile_X01_Y00_io2f_17_ready;
	assign Tile_X01_Y00_io2f_17_ready = {Tile_X01_Y01_SB_T4_NORTH_SB_IN_B17_ready, Tile_X01_Y01_SB_T3_NORTH_SB_IN_B17_ready, Tile_X01_Y01_SB_T2_NORTH_SB_IN_B17_ready, Tile_X01_Y01_SB_T1_NORTH_SB_IN_B17_ready, Tile_X01_Y01_SB_T0_NORTH_SB_IN_B17_ready};
	wire [4:0] Tile_X01_Y00_io2f_1_ready;
	assign Tile_X01_Y00_io2f_1_ready = {Tile_X01_Y01_SB_T4_NORTH_SB_IN_B1_ready, Tile_X01_Y01_SB_T3_NORTH_SB_IN_B1_ready, Tile_X01_Y01_SB_T2_NORTH_SB_IN_B1_ready, Tile_X01_Y01_SB_T1_NORTH_SB_IN_B1_ready, Tile_X01_Y01_SB_T0_NORTH_SB_IN_B1_ready};
	wire [15:0] Tile_X01_Y00_tile_id;
	assign Tile_X01_Y00_tile_id = {Tile_X01_Y00_lo[7], Tile_X01_Y00_lo[7], Tile_X01_Y00_lo[6], Tile_X01_Y00_lo[6], Tile_X01_Y00_lo[5], Tile_X01_Y00_lo[5], Tile_X01_Y00_lo[4], Tile_X01_Y00_hi[4], Tile_X01_Y00_lo[3], Tile_X01_Y00_lo[3], Tile_X01_Y00_lo[2], Tile_X01_Y00_lo[2], Tile_X01_Y00_lo[1], Tile_X01_Y00_lo[1], Tile_X01_Y00_lo[0], Tile_X01_Y00_lo[0]};
	Tile_IOCoreReadyValid Tile_X01_Y00(
		.clk(clk),
		.clk_out(Tile_X01_Y00_clk_out),
		.config_config_addr(Tile_X01_Y00_config_config_addr),
		.config_config_data(Tile_X01_Y00_config_config_data),
		.config_out_config_addr(Tile_X01_Y00_config_out_config_addr),
		.config_out_config_data(Tile_X01_Y00_config_out_config_data),
		.config_out_read(Tile_X01_Y00_config_out_read),
		.config_out_write(Tile_X01_Y00_config_out_write),
		.config_read(PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[64]),
		.config_write(PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[65]),
		.f2io_1(Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B1),
		.f2io_17(Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B17),
		.f2io_17_ready(Tile_X01_Y00_f2io_17_ready),
		.f2io_17_valid(Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B17_valid),
		.f2io_1_ready(Tile_X01_Y00_f2io_1_ready),
		.f2io_1_valid(Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B1_valid),
		.flush(PipelineRegister_inst1$Register_inst0$reg_P1_inst0_out),
		.flush_out(Tile_X01_Y00_flush_out),
		.glb2io_1(glb2io_1_X01_Y00),
		.glb2io_17(glb2io_17_X01_Y00),
		.glb2io_17_ready(Tile_X01_Y00_glb2io_17_ready),
		.glb2io_17_valid(glb2io_17_X01_Y00_valid),
		.glb2io_1_ready(Tile_X01_Y00_glb2io_1_ready),
		.glb2io_1_valid(glb2io_1_X01_Y00_valid),
		.hi(Tile_X01_Y00_hi),
		.io2f_1(Tile_X01_Y00_io2f_1),
		.io2f_17(Tile_X01_Y00_io2f_17),
		.io2f_17_ready(Tile_X01_Y00_io2f_17_ready),
		.io2f_17_valid(Tile_X01_Y00_io2f_17_valid),
		.io2f_1_ready(Tile_X01_Y00_io2f_1_ready),
		.io2f_1_valid(Tile_X01_Y00_io2f_1_valid),
		.io2glb_1(Tile_X01_Y00_io2glb_1),
		.io2glb_17(Tile_X01_Y00_io2glb_17),
		.io2glb_17_ready(io2glb_17_X01_Y00_ready),
		.io2glb_17_valid(Tile_X01_Y00_io2glb_17_valid),
		.io2glb_1_ready(io2glb_1_X01_Y00_ready),
		.io2glb_1_valid(Tile_X01_Y00_io2glb_1_valid),
		.lo(Tile_X01_Y00_lo),
		.read_config_data(Tile_X01_Y00_read_config_data),
		.read_config_data_in(const_0_32_out),
		.reset(reset),
		.reset_out(Tile_X01_Y00_reset_out),
		.stall(self_stall_out[1:1]),
		.stall_out(Tile_X01_Y00_stall_out),
		.tile_id(Tile_X01_Y00_tile_id)
	);
	wire [15:0] Tile_X01_Y01_tile_id;
	assign Tile_X01_Y01_tile_id = {Tile_X01_Y01_lo[7], Tile_X01_Y01_lo[7], Tile_X01_Y01_lo[6], Tile_X01_Y01_lo[6], Tile_X01_Y01_lo[5], Tile_X01_Y01_lo[5], Tile_X01_Y01_lo[4], Tile_X01_Y01_hi[4], Tile_X01_Y01_lo[3], Tile_X01_Y01_lo[3], Tile_X01_Y01_lo[2], Tile_X01_Y01_lo[2], Tile_X01_Y01_lo[1], Tile_X01_Y01_lo[1], Tile_X01_Y01_lo[0], Tile_X01_Y01_hi[0]};
	Tile_PE Tile_X01_Y01(
		.SB_T0_EAST_SB_IN_B1(Tile_X02_Y01_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_EAST_SB_IN_B17(Tile_X02_Y01_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_EAST_SB_IN_B17_ready(Tile_X01_Y01_SB_T0_EAST_SB_IN_B17_ready),
		.SB_T0_EAST_SB_IN_B17_valid(Tile_X02_Y01_SB_T0_WEST_SB_OUT_B17_valid),
		.SB_T0_EAST_SB_IN_B1_ready(Tile_X01_Y01_SB_T0_EAST_SB_IN_B1_ready),
		.SB_T0_EAST_SB_IN_B1_valid(Tile_X02_Y01_SB_T0_WEST_SB_OUT_B1_valid),
		.SB_T0_EAST_SB_OUT_B1(Tile_X01_Y01_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_EAST_SB_OUT_B17(Tile_X01_Y01_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_EAST_SB_OUT_B17_ready(Tile_X02_Y01_SB_T0_WEST_SB_IN_B17_ready),
		.SB_T0_EAST_SB_OUT_B17_valid(Tile_X01_Y01_SB_T0_EAST_SB_OUT_B17_valid),
		.SB_T0_EAST_SB_OUT_B1_ready(Tile_X02_Y01_SB_T0_WEST_SB_IN_B1_ready),
		.SB_T0_EAST_SB_OUT_B1_valid(Tile_X01_Y01_SB_T0_EAST_SB_OUT_B1_valid),
		.SB_T0_NORTH_SB_IN_B1(Tile_X01_Y00_io2f_1),
		.SB_T0_NORTH_SB_IN_B17(Tile_X01_Y00_io2f_17),
		.SB_T0_NORTH_SB_IN_B17_ready(Tile_X01_Y01_SB_T0_NORTH_SB_IN_B17_ready),
		.SB_T0_NORTH_SB_IN_B17_valid(Tile_X01_Y00_io2f_17_valid),
		.SB_T0_NORTH_SB_IN_B1_ready(Tile_X01_Y01_SB_T0_NORTH_SB_IN_B1_ready),
		.SB_T0_NORTH_SB_IN_B1_valid(Tile_X01_Y00_io2f_1_valid),
		.SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_OUT_B17(Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_OUT_B17_ready(Tile_X01_Y00_f2io_17_ready),
		.SB_T0_NORTH_SB_OUT_B17_valid(Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B17_valid),
		.SB_T0_NORTH_SB_OUT_B1_ready(Tile_X01_Y00_f2io_1_ready),
		.SB_T0_NORTH_SB_OUT_B1_valid(Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B1_valid),
		.SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_IN_B17(Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_IN_B17_ready(Tile_X01_Y01_SB_T0_SOUTH_SB_IN_B17_ready),
		.SB_T0_SOUTH_SB_IN_B17_valid(Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B17_valid),
		.SB_T0_SOUTH_SB_IN_B1_ready(Tile_X01_Y01_SB_T0_SOUTH_SB_IN_B1_ready),
		.SB_T0_SOUTH_SB_IN_B1_valid(Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B1_valid),
		.SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_OUT_B17(Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_OUT_B17_ready(Tile_X01_Y02_SB_T0_NORTH_SB_IN_B17_ready),
		.SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B17_valid),
		.SB_T0_SOUTH_SB_OUT_B1_ready(Tile_X01_Y02_SB_T0_NORTH_SB_IN_B1_ready),
		.SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B1_valid),
		.SB_T0_WEST_SB_IN_B1(Tile_X00_Y01_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_WEST_SB_IN_B17(Tile_X00_Y01_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_WEST_SB_IN_B17_ready(Tile_X01_Y01_SB_T0_WEST_SB_IN_B17_ready),
		.SB_T0_WEST_SB_IN_B17_valid(Tile_X00_Y01_SB_T0_EAST_SB_OUT_B17_valid),
		.SB_T0_WEST_SB_IN_B1_ready(Tile_X01_Y01_SB_T0_WEST_SB_IN_B1_ready),
		.SB_T0_WEST_SB_IN_B1_valid(Tile_X00_Y01_SB_T0_EAST_SB_OUT_B1_valid),
		.SB_T0_WEST_SB_OUT_B1(Tile_X01_Y01_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_WEST_SB_OUT_B17(Tile_X01_Y01_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_WEST_SB_OUT_B17_ready(Tile_X00_Y01_SB_T0_EAST_SB_IN_B17_ready),
		.SB_T0_WEST_SB_OUT_B17_valid(Tile_X01_Y01_SB_T0_WEST_SB_OUT_B17_valid),
		.SB_T0_WEST_SB_OUT_B1_ready(Tile_X00_Y01_SB_T0_EAST_SB_IN_B1_ready),
		.SB_T0_WEST_SB_OUT_B1_valid(Tile_X01_Y01_SB_T0_WEST_SB_OUT_B1_valid),
		.SB_T1_EAST_SB_IN_B1(Tile_X02_Y01_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_EAST_SB_IN_B17(Tile_X02_Y01_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_EAST_SB_IN_B17_ready(Tile_X01_Y01_SB_T1_EAST_SB_IN_B17_ready),
		.SB_T1_EAST_SB_IN_B17_valid(Tile_X02_Y01_SB_T1_WEST_SB_OUT_B17_valid),
		.SB_T1_EAST_SB_IN_B1_ready(Tile_X01_Y01_SB_T1_EAST_SB_IN_B1_ready),
		.SB_T1_EAST_SB_IN_B1_valid(Tile_X02_Y01_SB_T1_WEST_SB_OUT_B1_valid),
		.SB_T1_EAST_SB_OUT_B1(Tile_X01_Y01_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_EAST_SB_OUT_B17(Tile_X01_Y01_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_EAST_SB_OUT_B17_ready(Tile_X02_Y01_SB_T1_WEST_SB_IN_B17_ready),
		.SB_T1_EAST_SB_OUT_B17_valid(Tile_X01_Y01_SB_T1_EAST_SB_OUT_B17_valid),
		.SB_T1_EAST_SB_OUT_B1_ready(Tile_X02_Y01_SB_T1_WEST_SB_IN_B1_ready),
		.SB_T1_EAST_SB_OUT_B1_valid(Tile_X01_Y01_SB_T1_EAST_SB_OUT_B1_valid),
		.SB_T1_NORTH_SB_IN_B1(Tile_X01_Y00_io2f_1),
		.SB_T1_NORTH_SB_IN_B17(Tile_X01_Y00_io2f_17),
		.SB_T1_NORTH_SB_IN_B17_ready(Tile_X01_Y01_SB_T1_NORTH_SB_IN_B17_ready),
		.SB_T1_NORTH_SB_IN_B17_valid(Tile_X01_Y00_io2f_17_valid),
		.SB_T1_NORTH_SB_IN_B1_ready(Tile_X01_Y01_SB_T1_NORTH_SB_IN_B1_ready),
		.SB_T1_NORTH_SB_IN_B1_valid(Tile_X01_Y00_io2f_1_valid),
		.SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y01_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_OUT_B17(Tile_X01_Y01_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T1_NORTH_SB_OUT_B17_valid(Tile_X01_Y01_SB_T1_NORTH_SB_OUT_B17_valid),
		.SB_T1_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T1_NORTH_SB_OUT_B1_valid(Tile_X01_Y01_SB_T1_NORTH_SB_OUT_B1_valid),
		.SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_IN_B17(Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_IN_B17_ready(Tile_X01_Y01_SB_T1_SOUTH_SB_IN_B17_ready),
		.SB_T1_SOUTH_SB_IN_B17_valid(Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B17_valid),
		.SB_T1_SOUTH_SB_IN_B1_ready(Tile_X01_Y01_SB_T1_SOUTH_SB_IN_B1_ready),
		.SB_T1_SOUTH_SB_IN_B1_valid(Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B1_valid),
		.SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_OUT_B17(Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_OUT_B17_ready(Tile_X01_Y02_SB_T1_NORTH_SB_IN_B17_ready),
		.SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B17_valid),
		.SB_T1_SOUTH_SB_OUT_B1_ready(Tile_X01_Y02_SB_T1_NORTH_SB_IN_B1_ready),
		.SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B1_valid),
		.SB_T1_WEST_SB_IN_B1(Tile_X00_Y01_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_WEST_SB_IN_B17(Tile_X00_Y01_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_WEST_SB_IN_B17_ready(Tile_X01_Y01_SB_T1_WEST_SB_IN_B17_ready),
		.SB_T1_WEST_SB_IN_B17_valid(Tile_X00_Y01_SB_T1_EAST_SB_OUT_B17_valid),
		.SB_T1_WEST_SB_IN_B1_ready(Tile_X01_Y01_SB_T1_WEST_SB_IN_B1_ready),
		.SB_T1_WEST_SB_IN_B1_valid(Tile_X00_Y01_SB_T1_EAST_SB_OUT_B1_valid),
		.SB_T1_WEST_SB_OUT_B1(Tile_X01_Y01_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_WEST_SB_OUT_B17(Tile_X01_Y01_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_WEST_SB_OUT_B17_ready(Tile_X00_Y01_SB_T1_EAST_SB_IN_B17_ready),
		.SB_T1_WEST_SB_OUT_B17_valid(Tile_X01_Y01_SB_T1_WEST_SB_OUT_B17_valid),
		.SB_T1_WEST_SB_OUT_B1_ready(Tile_X00_Y01_SB_T1_EAST_SB_IN_B1_ready),
		.SB_T1_WEST_SB_OUT_B1_valid(Tile_X01_Y01_SB_T1_WEST_SB_OUT_B1_valid),
		.SB_T2_EAST_SB_IN_B1(Tile_X02_Y01_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_EAST_SB_IN_B17(Tile_X02_Y01_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_EAST_SB_IN_B17_ready(Tile_X01_Y01_SB_T2_EAST_SB_IN_B17_ready),
		.SB_T2_EAST_SB_IN_B17_valid(Tile_X02_Y01_SB_T2_WEST_SB_OUT_B17_valid),
		.SB_T2_EAST_SB_IN_B1_ready(Tile_X01_Y01_SB_T2_EAST_SB_IN_B1_ready),
		.SB_T2_EAST_SB_IN_B1_valid(Tile_X02_Y01_SB_T2_WEST_SB_OUT_B1_valid),
		.SB_T2_EAST_SB_OUT_B1(Tile_X01_Y01_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_EAST_SB_OUT_B17(Tile_X01_Y01_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_EAST_SB_OUT_B17_ready(Tile_X02_Y01_SB_T2_WEST_SB_IN_B17_ready),
		.SB_T2_EAST_SB_OUT_B17_valid(Tile_X01_Y01_SB_T2_EAST_SB_OUT_B17_valid),
		.SB_T2_EAST_SB_OUT_B1_ready(Tile_X02_Y01_SB_T2_WEST_SB_IN_B1_ready),
		.SB_T2_EAST_SB_OUT_B1_valid(Tile_X01_Y01_SB_T2_EAST_SB_OUT_B1_valid),
		.SB_T2_NORTH_SB_IN_B1(Tile_X01_Y00_io2f_1),
		.SB_T2_NORTH_SB_IN_B17(Tile_X01_Y00_io2f_17),
		.SB_T2_NORTH_SB_IN_B17_ready(Tile_X01_Y01_SB_T2_NORTH_SB_IN_B17_ready),
		.SB_T2_NORTH_SB_IN_B17_valid(Tile_X01_Y00_io2f_17_valid),
		.SB_T2_NORTH_SB_IN_B1_ready(Tile_X01_Y01_SB_T2_NORTH_SB_IN_B1_ready),
		.SB_T2_NORTH_SB_IN_B1_valid(Tile_X01_Y00_io2f_1_valid),
		.SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y01_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_OUT_B17(Tile_X01_Y01_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T2_NORTH_SB_OUT_B17_valid(Tile_X01_Y01_SB_T2_NORTH_SB_OUT_B17_valid),
		.SB_T2_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T2_NORTH_SB_OUT_B1_valid(Tile_X01_Y01_SB_T2_NORTH_SB_OUT_B1_valid),
		.SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_IN_B17(Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_IN_B17_ready(Tile_X01_Y01_SB_T2_SOUTH_SB_IN_B17_ready),
		.SB_T2_SOUTH_SB_IN_B17_valid(Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B17_valid),
		.SB_T2_SOUTH_SB_IN_B1_ready(Tile_X01_Y01_SB_T2_SOUTH_SB_IN_B1_ready),
		.SB_T2_SOUTH_SB_IN_B1_valid(Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B1_valid),
		.SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_OUT_B17(Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_OUT_B17_ready(Tile_X01_Y02_SB_T2_NORTH_SB_IN_B17_ready),
		.SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B17_valid),
		.SB_T2_SOUTH_SB_OUT_B1_ready(Tile_X01_Y02_SB_T2_NORTH_SB_IN_B1_ready),
		.SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B1_valid),
		.SB_T2_WEST_SB_IN_B1(Tile_X00_Y01_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_WEST_SB_IN_B17(Tile_X00_Y01_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_WEST_SB_IN_B17_ready(Tile_X01_Y01_SB_T2_WEST_SB_IN_B17_ready),
		.SB_T2_WEST_SB_IN_B17_valid(Tile_X00_Y01_SB_T2_EAST_SB_OUT_B17_valid),
		.SB_T2_WEST_SB_IN_B1_ready(Tile_X01_Y01_SB_T2_WEST_SB_IN_B1_ready),
		.SB_T2_WEST_SB_IN_B1_valid(Tile_X00_Y01_SB_T2_EAST_SB_OUT_B1_valid),
		.SB_T2_WEST_SB_OUT_B1(Tile_X01_Y01_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_WEST_SB_OUT_B17(Tile_X01_Y01_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_WEST_SB_OUT_B17_ready(Tile_X00_Y01_SB_T2_EAST_SB_IN_B17_ready),
		.SB_T2_WEST_SB_OUT_B17_valid(Tile_X01_Y01_SB_T2_WEST_SB_OUT_B17_valid),
		.SB_T2_WEST_SB_OUT_B1_ready(Tile_X00_Y01_SB_T2_EAST_SB_IN_B1_ready),
		.SB_T2_WEST_SB_OUT_B1_valid(Tile_X01_Y01_SB_T2_WEST_SB_OUT_B1_valid),
		.SB_T3_EAST_SB_IN_B1(Tile_X02_Y01_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_EAST_SB_IN_B17(Tile_X02_Y01_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_EAST_SB_IN_B17_ready(Tile_X01_Y01_SB_T3_EAST_SB_IN_B17_ready),
		.SB_T3_EAST_SB_IN_B17_valid(Tile_X02_Y01_SB_T3_WEST_SB_OUT_B17_valid),
		.SB_T3_EAST_SB_IN_B1_ready(Tile_X01_Y01_SB_T3_EAST_SB_IN_B1_ready),
		.SB_T3_EAST_SB_IN_B1_valid(Tile_X02_Y01_SB_T3_WEST_SB_OUT_B1_valid),
		.SB_T3_EAST_SB_OUT_B1(Tile_X01_Y01_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_EAST_SB_OUT_B17(Tile_X01_Y01_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_EAST_SB_OUT_B17_ready(Tile_X02_Y01_SB_T3_WEST_SB_IN_B17_ready),
		.SB_T3_EAST_SB_OUT_B17_valid(Tile_X01_Y01_SB_T3_EAST_SB_OUT_B17_valid),
		.SB_T3_EAST_SB_OUT_B1_ready(Tile_X02_Y01_SB_T3_WEST_SB_IN_B1_ready),
		.SB_T3_EAST_SB_OUT_B1_valid(Tile_X01_Y01_SB_T3_EAST_SB_OUT_B1_valid),
		.SB_T3_NORTH_SB_IN_B1(Tile_X01_Y00_io2f_1),
		.SB_T3_NORTH_SB_IN_B17(Tile_X01_Y00_io2f_17),
		.SB_T3_NORTH_SB_IN_B17_ready(Tile_X01_Y01_SB_T3_NORTH_SB_IN_B17_ready),
		.SB_T3_NORTH_SB_IN_B17_valid(Tile_X01_Y00_io2f_17_valid),
		.SB_T3_NORTH_SB_IN_B1_ready(Tile_X01_Y01_SB_T3_NORTH_SB_IN_B1_ready),
		.SB_T3_NORTH_SB_IN_B1_valid(Tile_X01_Y00_io2f_1_valid),
		.SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y01_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_OUT_B17(Tile_X01_Y01_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T3_NORTH_SB_OUT_B17_valid(Tile_X01_Y01_SB_T3_NORTH_SB_OUT_B17_valid),
		.SB_T3_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T3_NORTH_SB_OUT_B1_valid(Tile_X01_Y01_SB_T3_NORTH_SB_OUT_B1_valid),
		.SB_T3_SOUTH_SB_IN_B1(Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_IN_B17(Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_IN_B17_ready(Tile_X01_Y01_SB_T3_SOUTH_SB_IN_B17_ready),
		.SB_T3_SOUTH_SB_IN_B17_valid(Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B17_valid),
		.SB_T3_SOUTH_SB_IN_B1_ready(Tile_X01_Y01_SB_T3_SOUTH_SB_IN_B1_ready),
		.SB_T3_SOUTH_SB_IN_B1_valid(Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B1_valid),
		.SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_OUT_B17(Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_OUT_B17_ready(Tile_X01_Y02_SB_T3_NORTH_SB_IN_B17_ready),
		.SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B17_valid),
		.SB_T3_SOUTH_SB_OUT_B1_ready(Tile_X01_Y02_SB_T3_NORTH_SB_IN_B1_ready),
		.SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B1_valid),
		.SB_T3_WEST_SB_IN_B1(Tile_X00_Y01_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_WEST_SB_IN_B17(Tile_X00_Y01_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_WEST_SB_IN_B17_ready(Tile_X01_Y01_SB_T3_WEST_SB_IN_B17_ready),
		.SB_T3_WEST_SB_IN_B17_valid(Tile_X00_Y01_SB_T3_EAST_SB_OUT_B17_valid),
		.SB_T3_WEST_SB_IN_B1_ready(Tile_X01_Y01_SB_T3_WEST_SB_IN_B1_ready),
		.SB_T3_WEST_SB_IN_B1_valid(Tile_X00_Y01_SB_T3_EAST_SB_OUT_B1_valid),
		.SB_T3_WEST_SB_OUT_B1(Tile_X01_Y01_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_WEST_SB_OUT_B17(Tile_X01_Y01_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_WEST_SB_OUT_B17_ready(Tile_X00_Y01_SB_T3_EAST_SB_IN_B17_ready),
		.SB_T3_WEST_SB_OUT_B17_valid(Tile_X01_Y01_SB_T3_WEST_SB_OUT_B17_valid),
		.SB_T3_WEST_SB_OUT_B1_ready(Tile_X00_Y01_SB_T3_EAST_SB_IN_B1_ready),
		.SB_T3_WEST_SB_OUT_B1_valid(Tile_X01_Y01_SB_T3_WEST_SB_OUT_B1_valid),
		.SB_T4_EAST_SB_IN_B1(Tile_X02_Y01_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_EAST_SB_IN_B17(Tile_X02_Y01_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_EAST_SB_IN_B17_ready(Tile_X01_Y01_SB_T4_EAST_SB_IN_B17_ready),
		.SB_T4_EAST_SB_IN_B17_valid(Tile_X02_Y01_SB_T4_WEST_SB_OUT_B17_valid),
		.SB_T4_EAST_SB_IN_B1_ready(Tile_X01_Y01_SB_T4_EAST_SB_IN_B1_ready),
		.SB_T4_EAST_SB_IN_B1_valid(Tile_X02_Y01_SB_T4_WEST_SB_OUT_B1_valid),
		.SB_T4_EAST_SB_OUT_B1(Tile_X01_Y01_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_EAST_SB_OUT_B17(Tile_X01_Y01_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_EAST_SB_OUT_B17_ready(Tile_X02_Y01_SB_T4_WEST_SB_IN_B17_ready),
		.SB_T4_EAST_SB_OUT_B17_valid(Tile_X01_Y01_SB_T4_EAST_SB_OUT_B17_valid),
		.SB_T4_EAST_SB_OUT_B1_ready(Tile_X02_Y01_SB_T4_WEST_SB_IN_B1_ready),
		.SB_T4_EAST_SB_OUT_B1_valid(Tile_X01_Y01_SB_T4_EAST_SB_OUT_B1_valid),
		.SB_T4_NORTH_SB_IN_B1(Tile_X01_Y00_io2f_1),
		.SB_T4_NORTH_SB_IN_B17(Tile_X01_Y00_io2f_17),
		.SB_T4_NORTH_SB_IN_B17_ready(Tile_X01_Y01_SB_T4_NORTH_SB_IN_B17_ready),
		.SB_T4_NORTH_SB_IN_B17_valid(Tile_X01_Y00_io2f_17_valid),
		.SB_T4_NORTH_SB_IN_B1_ready(Tile_X01_Y01_SB_T4_NORTH_SB_IN_B1_ready),
		.SB_T4_NORTH_SB_IN_B1_valid(Tile_X01_Y00_io2f_1_valid),
		.SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y01_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_OUT_B17(Tile_X01_Y01_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T4_NORTH_SB_OUT_B17_valid(Tile_X01_Y01_SB_T4_NORTH_SB_OUT_B17_valid),
		.SB_T4_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T4_NORTH_SB_OUT_B1_valid(Tile_X01_Y01_SB_T4_NORTH_SB_OUT_B1_valid),
		.SB_T4_SOUTH_SB_IN_B1(Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_IN_B17(Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_IN_B17_ready(Tile_X01_Y01_SB_T4_SOUTH_SB_IN_B17_ready),
		.SB_T4_SOUTH_SB_IN_B17_valid(Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B17_valid),
		.SB_T4_SOUTH_SB_IN_B1_ready(Tile_X01_Y01_SB_T4_SOUTH_SB_IN_B1_ready),
		.SB_T4_SOUTH_SB_IN_B1_valid(Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B1_valid),
		.SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_OUT_B17(Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_OUT_B17_ready(Tile_X01_Y02_SB_T4_NORTH_SB_IN_B17_ready),
		.SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B17_valid),
		.SB_T4_SOUTH_SB_OUT_B1_ready(Tile_X01_Y02_SB_T4_NORTH_SB_IN_B1_ready),
		.SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B1_valid),
		.SB_T4_WEST_SB_IN_B1(Tile_X00_Y01_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_WEST_SB_IN_B17(Tile_X00_Y01_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_WEST_SB_IN_B17_ready(Tile_X01_Y01_SB_T4_WEST_SB_IN_B17_ready),
		.SB_T4_WEST_SB_IN_B17_valid(Tile_X00_Y01_SB_T4_EAST_SB_OUT_B17_valid),
		.SB_T4_WEST_SB_IN_B1_ready(Tile_X01_Y01_SB_T4_WEST_SB_IN_B1_ready),
		.SB_T4_WEST_SB_IN_B1_valid(Tile_X00_Y01_SB_T4_EAST_SB_OUT_B1_valid),
		.SB_T4_WEST_SB_OUT_B1(Tile_X01_Y01_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_WEST_SB_OUT_B17(Tile_X01_Y01_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_WEST_SB_OUT_B17_ready(Tile_X00_Y01_SB_T4_EAST_SB_IN_B17_ready),
		.SB_T4_WEST_SB_OUT_B17_valid(Tile_X01_Y01_SB_T4_WEST_SB_OUT_B17_valid),
		.SB_T4_WEST_SB_OUT_B1_ready(Tile_X00_Y01_SB_T4_EAST_SB_IN_B1_ready),
		.SB_T4_WEST_SB_OUT_B1_valid(Tile_X01_Y01_SB_T4_WEST_SB_OUT_B1_valid),
		.clk(Tile_X01_Y00_clk_out),
		.clk_out(Tile_X01_Y01_clk_out),
		.clk_pass_through(coreir_wrapInClock_inst1_out),
		.clk_pass_through_out_bot(Tile_X01_Y01_clk_pass_through_out_bot),
		.clk_pass_through_out_right(Tile_X01_Y01_clk_pass_through_out_right),
		.config_config_addr(Tile_X01_Y00_config_out_config_addr),
		.config_config_data(Tile_X01_Y00_config_out_config_data),
		.config_out_config_addr(Tile_X01_Y01_config_out_config_addr),
		.config_out_config_data(Tile_X01_Y01_config_out_config_data),
		.config_out_read(Tile_X01_Y01_config_out_read),
		.config_out_write(Tile_X01_Y01_config_out_write),
		.config_read(Tile_X01_Y00_config_out_read),
		.config_write(Tile_X01_Y00_config_out_write),
		.flush(Tile_X01_Y00_flush_out),
		.flush_out(Tile_X01_Y01_flush_out),
		.hi(Tile_X01_Y01_hi),
		.lo(Tile_X01_Y01_lo),
		.read_config_data(Tile_X01_Y01_read_config_data),
		.read_config_data_in(Tile_X01_Y00_read_config_data),
		.reset(Tile_X01_Y00_reset_out),
		.reset_out(Tile_X01_Y01_reset_out),
		.stall(Tile_X01_Y00_stall_out),
		.stall_out(Tile_X01_Y01_stall_out),
		.tile_id(Tile_X01_Y01_tile_id)
	);
	wire [15:0] Tile_X01_Y02_tile_id;
	assign Tile_X01_Y02_tile_id = {Tile_X01_Y02_lo[7], Tile_X01_Y02_lo[7], Tile_X01_Y02_lo[6], Tile_X01_Y02_lo[6], Tile_X01_Y02_lo[5], Tile_X01_Y02_lo[5], Tile_X01_Y02_lo[4], Tile_X01_Y02_hi[4], Tile_X01_Y02_lo[3], Tile_X01_Y02_lo[3], Tile_X01_Y02_lo[2], Tile_X01_Y02_lo[2], Tile_X01_Y02_lo[1], Tile_X01_Y02_lo[1], Tile_X01_Y02_hi[1], Tile_X01_Y02_lo[0]};
	Tile_PE Tile_X01_Y02(
		.SB_T0_EAST_SB_IN_B1(Tile_X02_Y02_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_EAST_SB_IN_B17(Tile_X02_Y02_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_EAST_SB_IN_B17_ready(Tile_X01_Y02_SB_T0_EAST_SB_IN_B17_ready),
		.SB_T0_EAST_SB_IN_B17_valid(Tile_X02_Y02_SB_T0_WEST_SB_OUT_B17_valid),
		.SB_T0_EAST_SB_IN_B1_ready(Tile_X01_Y02_SB_T0_EAST_SB_IN_B1_ready),
		.SB_T0_EAST_SB_IN_B1_valid(Tile_X02_Y02_SB_T0_WEST_SB_OUT_B1_valid),
		.SB_T0_EAST_SB_OUT_B1(Tile_X01_Y02_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_EAST_SB_OUT_B17(Tile_X01_Y02_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_EAST_SB_OUT_B17_ready(Tile_X02_Y02_SB_T0_WEST_SB_IN_B17_ready),
		.SB_T0_EAST_SB_OUT_B17_valid(Tile_X01_Y02_SB_T0_EAST_SB_OUT_B17_valid),
		.SB_T0_EAST_SB_OUT_B1_ready(Tile_X02_Y02_SB_T0_WEST_SB_IN_B1_ready),
		.SB_T0_EAST_SB_OUT_B1_valid(Tile_X01_Y02_SB_T0_EAST_SB_OUT_B1_valid),
		.SB_T0_NORTH_SB_IN_B1(Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_IN_B17(Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_IN_B17_ready(Tile_X01_Y02_SB_T0_NORTH_SB_IN_B17_ready),
		.SB_T0_NORTH_SB_IN_B17_valid(Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B17_valid),
		.SB_T0_NORTH_SB_IN_B1_ready(Tile_X01_Y02_SB_T0_NORTH_SB_IN_B1_ready),
		.SB_T0_NORTH_SB_IN_B1_valid(Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B1_valid),
		.SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_OUT_B17(Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_OUT_B17_ready(Tile_X01_Y01_SB_T0_SOUTH_SB_IN_B17_ready),
		.SB_T0_NORTH_SB_OUT_B17_valid(Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B17_valid),
		.SB_T0_NORTH_SB_OUT_B1_ready(Tile_X01_Y01_SB_T0_SOUTH_SB_IN_B1_ready),
		.SB_T0_NORTH_SB_OUT_B1_valid(Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B1_valid),
		.SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_IN_B17(Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_IN_B17_ready(Tile_X01_Y02_SB_T0_SOUTH_SB_IN_B17_ready),
		.SB_T0_SOUTH_SB_IN_B17_valid(Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B17_valid),
		.SB_T0_SOUTH_SB_IN_B1_ready(Tile_X01_Y02_SB_T0_SOUTH_SB_IN_B1_ready),
		.SB_T0_SOUTH_SB_IN_B1_valid(Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B1_valid),
		.SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_OUT_B17(Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_OUT_B17_ready(Tile_X01_Y03_SB_T0_NORTH_SB_IN_B17_ready),
		.SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B17_valid),
		.SB_T0_SOUTH_SB_OUT_B1_ready(Tile_X01_Y03_SB_T0_NORTH_SB_IN_B1_ready),
		.SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B1_valid),
		.SB_T0_WEST_SB_IN_B1(Tile_X00_Y02_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_WEST_SB_IN_B17(Tile_X00_Y02_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_WEST_SB_IN_B17_ready(Tile_X01_Y02_SB_T0_WEST_SB_IN_B17_ready),
		.SB_T0_WEST_SB_IN_B17_valid(Tile_X00_Y02_SB_T0_EAST_SB_OUT_B17_valid),
		.SB_T0_WEST_SB_IN_B1_ready(Tile_X01_Y02_SB_T0_WEST_SB_IN_B1_ready),
		.SB_T0_WEST_SB_IN_B1_valid(Tile_X00_Y02_SB_T0_EAST_SB_OUT_B1_valid),
		.SB_T0_WEST_SB_OUT_B1(Tile_X01_Y02_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_WEST_SB_OUT_B17(Tile_X01_Y02_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_WEST_SB_OUT_B17_ready(Tile_X00_Y02_SB_T0_EAST_SB_IN_B17_ready),
		.SB_T0_WEST_SB_OUT_B17_valid(Tile_X01_Y02_SB_T0_WEST_SB_OUT_B17_valid),
		.SB_T0_WEST_SB_OUT_B1_ready(Tile_X00_Y02_SB_T0_EAST_SB_IN_B1_ready),
		.SB_T0_WEST_SB_OUT_B1_valid(Tile_X01_Y02_SB_T0_WEST_SB_OUT_B1_valid),
		.SB_T1_EAST_SB_IN_B1(Tile_X02_Y02_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_EAST_SB_IN_B17(Tile_X02_Y02_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_EAST_SB_IN_B17_ready(Tile_X01_Y02_SB_T1_EAST_SB_IN_B17_ready),
		.SB_T1_EAST_SB_IN_B17_valid(Tile_X02_Y02_SB_T1_WEST_SB_OUT_B17_valid),
		.SB_T1_EAST_SB_IN_B1_ready(Tile_X01_Y02_SB_T1_EAST_SB_IN_B1_ready),
		.SB_T1_EAST_SB_IN_B1_valid(Tile_X02_Y02_SB_T1_WEST_SB_OUT_B1_valid),
		.SB_T1_EAST_SB_OUT_B1(Tile_X01_Y02_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_EAST_SB_OUT_B17(Tile_X01_Y02_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_EAST_SB_OUT_B17_ready(Tile_X02_Y02_SB_T1_WEST_SB_IN_B17_ready),
		.SB_T1_EAST_SB_OUT_B17_valid(Tile_X01_Y02_SB_T1_EAST_SB_OUT_B17_valid),
		.SB_T1_EAST_SB_OUT_B1_ready(Tile_X02_Y02_SB_T1_WEST_SB_IN_B1_ready),
		.SB_T1_EAST_SB_OUT_B1_valid(Tile_X01_Y02_SB_T1_EAST_SB_OUT_B1_valid),
		.SB_T1_NORTH_SB_IN_B1(Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_IN_B17(Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_IN_B17_ready(Tile_X01_Y02_SB_T1_NORTH_SB_IN_B17_ready),
		.SB_T1_NORTH_SB_IN_B17_valid(Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B17_valid),
		.SB_T1_NORTH_SB_IN_B1_ready(Tile_X01_Y02_SB_T1_NORTH_SB_IN_B1_ready),
		.SB_T1_NORTH_SB_IN_B1_valid(Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B1_valid),
		.SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_OUT_B17(Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_OUT_B17_ready(Tile_X01_Y01_SB_T1_SOUTH_SB_IN_B17_ready),
		.SB_T1_NORTH_SB_OUT_B17_valid(Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B17_valid),
		.SB_T1_NORTH_SB_OUT_B1_ready(Tile_X01_Y01_SB_T1_SOUTH_SB_IN_B1_ready),
		.SB_T1_NORTH_SB_OUT_B1_valid(Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B1_valid),
		.SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_IN_B17(Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_IN_B17_ready(Tile_X01_Y02_SB_T1_SOUTH_SB_IN_B17_ready),
		.SB_T1_SOUTH_SB_IN_B17_valid(Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B17_valid),
		.SB_T1_SOUTH_SB_IN_B1_ready(Tile_X01_Y02_SB_T1_SOUTH_SB_IN_B1_ready),
		.SB_T1_SOUTH_SB_IN_B1_valid(Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B1_valid),
		.SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_OUT_B17(Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_OUT_B17_ready(Tile_X01_Y03_SB_T1_NORTH_SB_IN_B17_ready),
		.SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B17_valid),
		.SB_T1_SOUTH_SB_OUT_B1_ready(Tile_X01_Y03_SB_T1_NORTH_SB_IN_B1_ready),
		.SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B1_valid),
		.SB_T1_WEST_SB_IN_B1(Tile_X00_Y02_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_WEST_SB_IN_B17(Tile_X00_Y02_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_WEST_SB_IN_B17_ready(Tile_X01_Y02_SB_T1_WEST_SB_IN_B17_ready),
		.SB_T1_WEST_SB_IN_B17_valid(Tile_X00_Y02_SB_T1_EAST_SB_OUT_B17_valid),
		.SB_T1_WEST_SB_IN_B1_ready(Tile_X01_Y02_SB_T1_WEST_SB_IN_B1_ready),
		.SB_T1_WEST_SB_IN_B1_valid(Tile_X00_Y02_SB_T1_EAST_SB_OUT_B1_valid),
		.SB_T1_WEST_SB_OUT_B1(Tile_X01_Y02_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_WEST_SB_OUT_B17(Tile_X01_Y02_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_WEST_SB_OUT_B17_ready(Tile_X00_Y02_SB_T1_EAST_SB_IN_B17_ready),
		.SB_T1_WEST_SB_OUT_B17_valid(Tile_X01_Y02_SB_T1_WEST_SB_OUT_B17_valid),
		.SB_T1_WEST_SB_OUT_B1_ready(Tile_X00_Y02_SB_T1_EAST_SB_IN_B1_ready),
		.SB_T1_WEST_SB_OUT_B1_valid(Tile_X01_Y02_SB_T1_WEST_SB_OUT_B1_valid),
		.SB_T2_EAST_SB_IN_B1(Tile_X02_Y02_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_EAST_SB_IN_B17(Tile_X02_Y02_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_EAST_SB_IN_B17_ready(Tile_X01_Y02_SB_T2_EAST_SB_IN_B17_ready),
		.SB_T2_EAST_SB_IN_B17_valid(Tile_X02_Y02_SB_T2_WEST_SB_OUT_B17_valid),
		.SB_T2_EAST_SB_IN_B1_ready(Tile_X01_Y02_SB_T2_EAST_SB_IN_B1_ready),
		.SB_T2_EAST_SB_IN_B1_valid(Tile_X02_Y02_SB_T2_WEST_SB_OUT_B1_valid),
		.SB_T2_EAST_SB_OUT_B1(Tile_X01_Y02_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_EAST_SB_OUT_B17(Tile_X01_Y02_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_EAST_SB_OUT_B17_ready(Tile_X02_Y02_SB_T2_WEST_SB_IN_B17_ready),
		.SB_T2_EAST_SB_OUT_B17_valid(Tile_X01_Y02_SB_T2_EAST_SB_OUT_B17_valid),
		.SB_T2_EAST_SB_OUT_B1_ready(Tile_X02_Y02_SB_T2_WEST_SB_IN_B1_ready),
		.SB_T2_EAST_SB_OUT_B1_valid(Tile_X01_Y02_SB_T2_EAST_SB_OUT_B1_valid),
		.SB_T2_NORTH_SB_IN_B1(Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_IN_B17(Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_IN_B17_ready(Tile_X01_Y02_SB_T2_NORTH_SB_IN_B17_ready),
		.SB_T2_NORTH_SB_IN_B17_valid(Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B17_valid),
		.SB_T2_NORTH_SB_IN_B1_ready(Tile_X01_Y02_SB_T2_NORTH_SB_IN_B1_ready),
		.SB_T2_NORTH_SB_IN_B1_valid(Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B1_valid),
		.SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_OUT_B17(Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_OUT_B17_ready(Tile_X01_Y01_SB_T2_SOUTH_SB_IN_B17_ready),
		.SB_T2_NORTH_SB_OUT_B17_valid(Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B17_valid),
		.SB_T2_NORTH_SB_OUT_B1_ready(Tile_X01_Y01_SB_T2_SOUTH_SB_IN_B1_ready),
		.SB_T2_NORTH_SB_OUT_B1_valid(Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B1_valid),
		.SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_IN_B17(Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_IN_B17_ready(Tile_X01_Y02_SB_T2_SOUTH_SB_IN_B17_ready),
		.SB_T2_SOUTH_SB_IN_B17_valid(Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B17_valid),
		.SB_T2_SOUTH_SB_IN_B1_ready(Tile_X01_Y02_SB_T2_SOUTH_SB_IN_B1_ready),
		.SB_T2_SOUTH_SB_IN_B1_valid(Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B1_valid),
		.SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_OUT_B17(Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_OUT_B17_ready(Tile_X01_Y03_SB_T2_NORTH_SB_IN_B17_ready),
		.SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B17_valid),
		.SB_T2_SOUTH_SB_OUT_B1_ready(Tile_X01_Y03_SB_T2_NORTH_SB_IN_B1_ready),
		.SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B1_valid),
		.SB_T2_WEST_SB_IN_B1(Tile_X00_Y02_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_WEST_SB_IN_B17(Tile_X00_Y02_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_WEST_SB_IN_B17_ready(Tile_X01_Y02_SB_T2_WEST_SB_IN_B17_ready),
		.SB_T2_WEST_SB_IN_B17_valid(Tile_X00_Y02_SB_T2_EAST_SB_OUT_B17_valid),
		.SB_T2_WEST_SB_IN_B1_ready(Tile_X01_Y02_SB_T2_WEST_SB_IN_B1_ready),
		.SB_T2_WEST_SB_IN_B1_valid(Tile_X00_Y02_SB_T2_EAST_SB_OUT_B1_valid),
		.SB_T2_WEST_SB_OUT_B1(Tile_X01_Y02_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_WEST_SB_OUT_B17(Tile_X01_Y02_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_WEST_SB_OUT_B17_ready(Tile_X00_Y02_SB_T2_EAST_SB_IN_B17_ready),
		.SB_T2_WEST_SB_OUT_B17_valid(Tile_X01_Y02_SB_T2_WEST_SB_OUT_B17_valid),
		.SB_T2_WEST_SB_OUT_B1_ready(Tile_X00_Y02_SB_T2_EAST_SB_IN_B1_ready),
		.SB_T2_WEST_SB_OUT_B1_valid(Tile_X01_Y02_SB_T2_WEST_SB_OUT_B1_valid),
		.SB_T3_EAST_SB_IN_B1(Tile_X02_Y02_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_EAST_SB_IN_B17(Tile_X02_Y02_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_EAST_SB_IN_B17_ready(Tile_X01_Y02_SB_T3_EAST_SB_IN_B17_ready),
		.SB_T3_EAST_SB_IN_B17_valid(Tile_X02_Y02_SB_T3_WEST_SB_OUT_B17_valid),
		.SB_T3_EAST_SB_IN_B1_ready(Tile_X01_Y02_SB_T3_EAST_SB_IN_B1_ready),
		.SB_T3_EAST_SB_IN_B1_valid(Tile_X02_Y02_SB_T3_WEST_SB_OUT_B1_valid),
		.SB_T3_EAST_SB_OUT_B1(Tile_X01_Y02_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_EAST_SB_OUT_B17(Tile_X01_Y02_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_EAST_SB_OUT_B17_ready(Tile_X02_Y02_SB_T3_WEST_SB_IN_B17_ready),
		.SB_T3_EAST_SB_OUT_B17_valid(Tile_X01_Y02_SB_T3_EAST_SB_OUT_B17_valid),
		.SB_T3_EAST_SB_OUT_B1_ready(Tile_X02_Y02_SB_T3_WEST_SB_IN_B1_ready),
		.SB_T3_EAST_SB_OUT_B1_valid(Tile_X01_Y02_SB_T3_EAST_SB_OUT_B1_valid),
		.SB_T3_NORTH_SB_IN_B1(Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_IN_B17(Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_IN_B17_ready(Tile_X01_Y02_SB_T3_NORTH_SB_IN_B17_ready),
		.SB_T3_NORTH_SB_IN_B17_valid(Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B17_valid),
		.SB_T3_NORTH_SB_IN_B1_ready(Tile_X01_Y02_SB_T3_NORTH_SB_IN_B1_ready),
		.SB_T3_NORTH_SB_IN_B1_valid(Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B1_valid),
		.SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_OUT_B17(Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_OUT_B17_ready(Tile_X01_Y01_SB_T3_SOUTH_SB_IN_B17_ready),
		.SB_T3_NORTH_SB_OUT_B17_valid(Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B17_valid),
		.SB_T3_NORTH_SB_OUT_B1_ready(Tile_X01_Y01_SB_T3_SOUTH_SB_IN_B1_ready),
		.SB_T3_NORTH_SB_OUT_B1_valid(Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B1_valid),
		.SB_T3_SOUTH_SB_IN_B1(Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_IN_B17(Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_IN_B17_ready(Tile_X01_Y02_SB_T3_SOUTH_SB_IN_B17_ready),
		.SB_T3_SOUTH_SB_IN_B17_valid(Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B17_valid),
		.SB_T3_SOUTH_SB_IN_B1_ready(Tile_X01_Y02_SB_T3_SOUTH_SB_IN_B1_ready),
		.SB_T3_SOUTH_SB_IN_B1_valid(Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B1_valid),
		.SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_OUT_B17(Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_OUT_B17_ready(Tile_X01_Y03_SB_T3_NORTH_SB_IN_B17_ready),
		.SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B17_valid),
		.SB_T3_SOUTH_SB_OUT_B1_ready(Tile_X01_Y03_SB_T3_NORTH_SB_IN_B1_ready),
		.SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B1_valid),
		.SB_T3_WEST_SB_IN_B1(Tile_X00_Y02_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_WEST_SB_IN_B17(Tile_X00_Y02_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_WEST_SB_IN_B17_ready(Tile_X01_Y02_SB_T3_WEST_SB_IN_B17_ready),
		.SB_T3_WEST_SB_IN_B17_valid(Tile_X00_Y02_SB_T3_EAST_SB_OUT_B17_valid),
		.SB_T3_WEST_SB_IN_B1_ready(Tile_X01_Y02_SB_T3_WEST_SB_IN_B1_ready),
		.SB_T3_WEST_SB_IN_B1_valid(Tile_X00_Y02_SB_T3_EAST_SB_OUT_B1_valid),
		.SB_T3_WEST_SB_OUT_B1(Tile_X01_Y02_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_WEST_SB_OUT_B17(Tile_X01_Y02_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_WEST_SB_OUT_B17_ready(Tile_X00_Y02_SB_T3_EAST_SB_IN_B17_ready),
		.SB_T3_WEST_SB_OUT_B17_valid(Tile_X01_Y02_SB_T3_WEST_SB_OUT_B17_valid),
		.SB_T3_WEST_SB_OUT_B1_ready(Tile_X00_Y02_SB_T3_EAST_SB_IN_B1_ready),
		.SB_T3_WEST_SB_OUT_B1_valid(Tile_X01_Y02_SB_T3_WEST_SB_OUT_B1_valid),
		.SB_T4_EAST_SB_IN_B1(Tile_X02_Y02_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_EAST_SB_IN_B17(Tile_X02_Y02_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_EAST_SB_IN_B17_ready(Tile_X01_Y02_SB_T4_EAST_SB_IN_B17_ready),
		.SB_T4_EAST_SB_IN_B17_valid(Tile_X02_Y02_SB_T4_WEST_SB_OUT_B17_valid),
		.SB_T4_EAST_SB_IN_B1_ready(Tile_X01_Y02_SB_T4_EAST_SB_IN_B1_ready),
		.SB_T4_EAST_SB_IN_B1_valid(Tile_X02_Y02_SB_T4_WEST_SB_OUT_B1_valid),
		.SB_T4_EAST_SB_OUT_B1(Tile_X01_Y02_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_EAST_SB_OUT_B17(Tile_X01_Y02_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_EAST_SB_OUT_B17_ready(Tile_X02_Y02_SB_T4_WEST_SB_IN_B17_ready),
		.SB_T4_EAST_SB_OUT_B17_valid(Tile_X01_Y02_SB_T4_EAST_SB_OUT_B17_valid),
		.SB_T4_EAST_SB_OUT_B1_ready(Tile_X02_Y02_SB_T4_WEST_SB_IN_B1_ready),
		.SB_T4_EAST_SB_OUT_B1_valid(Tile_X01_Y02_SB_T4_EAST_SB_OUT_B1_valid),
		.SB_T4_NORTH_SB_IN_B1(Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_IN_B17(Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_IN_B17_ready(Tile_X01_Y02_SB_T4_NORTH_SB_IN_B17_ready),
		.SB_T4_NORTH_SB_IN_B17_valid(Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B17_valid),
		.SB_T4_NORTH_SB_IN_B1_ready(Tile_X01_Y02_SB_T4_NORTH_SB_IN_B1_ready),
		.SB_T4_NORTH_SB_IN_B1_valid(Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B1_valid),
		.SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_OUT_B17(Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_OUT_B17_ready(Tile_X01_Y01_SB_T4_SOUTH_SB_IN_B17_ready),
		.SB_T4_NORTH_SB_OUT_B17_valid(Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B17_valid),
		.SB_T4_NORTH_SB_OUT_B1_ready(Tile_X01_Y01_SB_T4_SOUTH_SB_IN_B1_ready),
		.SB_T4_NORTH_SB_OUT_B1_valid(Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B1_valid),
		.SB_T4_SOUTH_SB_IN_B1(Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_IN_B17(Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_IN_B17_ready(Tile_X01_Y02_SB_T4_SOUTH_SB_IN_B17_ready),
		.SB_T4_SOUTH_SB_IN_B17_valid(Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B17_valid),
		.SB_T4_SOUTH_SB_IN_B1_ready(Tile_X01_Y02_SB_T4_SOUTH_SB_IN_B1_ready),
		.SB_T4_SOUTH_SB_IN_B1_valid(Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B1_valid),
		.SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_OUT_B17(Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_OUT_B17_ready(Tile_X01_Y03_SB_T4_NORTH_SB_IN_B17_ready),
		.SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B17_valid),
		.SB_T4_SOUTH_SB_OUT_B1_ready(Tile_X01_Y03_SB_T4_NORTH_SB_IN_B1_ready),
		.SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B1_valid),
		.SB_T4_WEST_SB_IN_B1(Tile_X00_Y02_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_WEST_SB_IN_B17(Tile_X00_Y02_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_WEST_SB_IN_B17_ready(Tile_X01_Y02_SB_T4_WEST_SB_IN_B17_ready),
		.SB_T4_WEST_SB_IN_B17_valid(Tile_X00_Y02_SB_T4_EAST_SB_OUT_B17_valid),
		.SB_T4_WEST_SB_IN_B1_ready(Tile_X01_Y02_SB_T4_WEST_SB_IN_B1_ready),
		.SB_T4_WEST_SB_IN_B1_valid(Tile_X00_Y02_SB_T4_EAST_SB_OUT_B1_valid),
		.SB_T4_WEST_SB_OUT_B1(Tile_X01_Y02_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_WEST_SB_OUT_B17(Tile_X01_Y02_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_WEST_SB_OUT_B17_ready(Tile_X00_Y02_SB_T4_EAST_SB_IN_B17_ready),
		.SB_T4_WEST_SB_OUT_B17_valid(Tile_X01_Y02_SB_T4_WEST_SB_OUT_B17_valid),
		.SB_T4_WEST_SB_OUT_B1_ready(Tile_X00_Y02_SB_T4_EAST_SB_IN_B1_ready),
		.SB_T4_WEST_SB_OUT_B1_valid(Tile_X01_Y02_SB_T4_WEST_SB_OUT_B1_valid),
		.clk(Tile_X01_Y01_clk_out),
		.clk_out(Tile_X01_Y02_clk_out),
		.clk_pass_through(Tile_X01_Y01_clk_pass_through_out_bot),
		.clk_pass_through_out_bot(Tile_X01_Y02_clk_pass_through_out_bot),
		.clk_pass_through_out_right(Tile_X01_Y02_clk_pass_through_out_right),
		.config_config_addr(Tile_X01_Y01_config_out_config_addr),
		.config_config_data(Tile_X01_Y01_config_out_config_data),
		.config_out_config_addr(Tile_X01_Y02_config_out_config_addr),
		.config_out_config_data(Tile_X01_Y02_config_out_config_data),
		.config_out_read(Tile_X01_Y02_config_out_read),
		.config_out_write(Tile_X01_Y02_config_out_write),
		.config_read(Tile_X01_Y01_config_out_read),
		.config_write(Tile_X01_Y01_config_out_write),
		.flush(Tile_X01_Y01_flush_out),
		.flush_out(Tile_X01_Y02_flush_out),
		.hi(Tile_X01_Y02_hi),
		.lo(Tile_X01_Y02_lo),
		.read_config_data(Tile_X01_Y02_read_config_data),
		.read_config_data_in(Tile_X01_Y01_read_config_data),
		.reset(Tile_X01_Y01_reset_out),
		.reset_out(Tile_X01_Y02_reset_out),
		.stall(Tile_X01_Y01_stall_out),
		.stall_out(Tile_X01_Y02_stall_out),
		.tile_id(Tile_X01_Y02_tile_id)
	);
	wire [15:0] Tile_X01_Y03_tile_id;
	assign Tile_X01_Y03_tile_id = {Tile_X01_Y03_lo[7], Tile_X01_Y03_lo[7], Tile_X01_Y03_lo[6], Tile_X01_Y03_lo[6], Tile_X01_Y03_lo[5], Tile_X01_Y03_lo[5], Tile_X01_Y03_lo[4], Tile_X01_Y03_hi[4], Tile_X01_Y03_lo[3], Tile_X01_Y03_lo[3], Tile_X01_Y03_lo[2], Tile_X01_Y03_lo[2], Tile_X01_Y03_lo[1], Tile_X01_Y03_lo[1], Tile_X01_Y03_hi[1], Tile_X01_Y03_hi[0]};
	Tile_PE Tile_X01_Y03(
		.SB_T0_EAST_SB_IN_B1(Tile_X02_Y03_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_EAST_SB_IN_B17(Tile_X02_Y03_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_EAST_SB_IN_B17_ready(Tile_X01_Y03_SB_T0_EAST_SB_IN_B17_ready),
		.SB_T0_EAST_SB_IN_B17_valid(Tile_X02_Y03_SB_T0_WEST_SB_OUT_B17_valid),
		.SB_T0_EAST_SB_IN_B1_ready(Tile_X01_Y03_SB_T0_EAST_SB_IN_B1_ready),
		.SB_T0_EAST_SB_IN_B1_valid(Tile_X02_Y03_SB_T0_WEST_SB_OUT_B1_valid),
		.SB_T0_EAST_SB_OUT_B1(Tile_X01_Y03_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_EAST_SB_OUT_B17(Tile_X01_Y03_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_EAST_SB_OUT_B17_ready(Tile_X02_Y03_SB_T0_WEST_SB_IN_B17_ready),
		.SB_T0_EAST_SB_OUT_B17_valid(Tile_X01_Y03_SB_T0_EAST_SB_OUT_B17_valid),
		.SB_T0_EAST_SB_OUT_B1_ready(Tile_X02_Y03_SB_T0_WEST_SB_IN_B1_ready),
		.SB_T0_EAST_SB_OUT_B1_valid(Tile_X01_Y03_SB_T0_EAST_SB_OUT_B1_valid),
		.SB_T0_NORTH_SB_IN_B1(Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_IN_B17(Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_IN_B17_ready(Tile_X01_Y03_SB_T0_NORTH_SB_IN_B17_ready),
		.SB_T0_NORTH_SB_IN_B17_valid(Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B17_valid),
		.SB_T0_NORTH_SB_IN_B1_ready(Tile_X01_Y03_SB_T0_NORTH_SB_IN_B1_ready),
		.SB_T0_NORTH_SB_IN_B1_valid(Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B1_valid),
		.SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_OUT_B17(Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_OUT_B17_ready(Tile_X01_Y02_SB_T0_SOUTH_SB_IN_B17_ready),
		.SB_T0_NORTH_SB_OUT_B17_valid(Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B17_valid),
		.SB_T0_NORTH_SB_OUT_B1_ready(Tile_X01_Y02_SB_T0_SOUTH_SB_IN_B1_ready),
		.SB_T0_NORTH_SB_OUT_B1_valid(Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B1_valid),
		.SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_IN_B17(Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_IN_B17_ready(Tile_X01_Y03_SB_T0_SOUTH_SB_IN_B17_ready),
		.SB_T0_SOUTH_SB_IN_B17_valid(Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B17_valid),
		.SB_T0_SOUTH_SB_IN_B1_ready(Tile_X01_Y03_SB_T0_SOUTH_SB_IN_B1_ready),
		.SB_T0_SOUTH_SB_IN_B1_valid(Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B1_valid),
		.SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_OUT_B17(Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_OUT_B17_ready(Tile_X01_Y04_SB_T0_NORTH_SB_IN_B17_ready),
		.SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B17_valid),
		.SB_T0_SOUTH_SB_OUT_B1_ready(Tile_X01_Y04_SB_T0_NORTH_SB_IN_B1_ready),
		.SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B1_valid),
		.SB_T0_WEST_SB_IN_B1(Tile_X00_Y03_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_WEST_SB_IN_B17(Tile_X00_Y03_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_WEST_SB_IN_B17_ready(Tile_X01_Y03_SB_T0_WEST_SB_IN_B17_ready),
		.SB_T0_WEST_SB_IN_B17_valid(Tile_X00_Y03_SB_T0_EAST_SB_OUT_B17_valid),
		.SB_T0_WEST_SB_IN_B1_ready(Tile_X01_Y03_SB_T0_WEST_SB_IN_B1_ready),
		.SB_T0_WEST_SB_IN_B1_valid(Tile_X00_Y03_SB_T0_EAST_SB_OUT_B1_valid),
		.SB_T0_WEST_SB_OUT_B1(Tile_X01_Y03_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_WEST_SB_OUT_B17(Tile_X01_Y03_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_WEST_SB_OUT_B17_ready(Tile_X00_Y03_SB_T0_EAST_SB_IN_B17_ready),
		.SB_T0_WEST_SB_OUT_B17_valid(Tile_X01_Y03_SB_T0_WEST_SB_OUT_B17_valid),
		.SB_T0_WEST_SB_OUT_B1_ready(Tile_X00_Y03_SB_T0_EAST_SB_IN_B1_ready),
		.SB_T0_WEST_SB_OUT_B1_valid(Tile_X01_Y03_SB_T0_WEST_SB_OUT_B1_valid),
		.SB_T1_EAST_SB_IN_B1(Tile_X02_Y03_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_EAST_SB_IN_B17(Tile_X02_Y03_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_EAST_SB_IN_B17_ready(Tile_X01_Y03_SB_T1_EAST_SB_IN_B17_ready),
		.SB_T1_EAST_SB_IN_B17_valid(Tile_X02_Y03_SB_T1_WEST_SB_OUT_B17_valid),
		.SB_T1_EAST_SB_IN_B1_ready(Tile_X01_Y03_SB_T1_EAST_SB_IN_B1_ready),
		.SB_T1_EAST_SB_IN_B1_valid(Tile_X02_Y03_SB_T1_WEST_SB_OUT_B1_valid),
		.SB_T1_EAST_SB_OUT_B1(Tile_X01_Y03_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_EAST_SB_OUT_B17(Tile_X01_Y03_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_EAST_SB_OUT_B17_ready(Tile_X02_Y03_SB_T1_WEST_SB_IN_B17_ready),
		.SB_T1_EAST_SB_OUT_B17_valid(Tile_X01_Y03_SB_T1_EAST_SB_OUT_B17_valid),
		.SB_T1_EAST_SB_OUT_B1_ready(Tile_X02_Y03_SB_T1_WEST_SB_IN_B1_ready),
		.SB_T1_EAST_SB_OUT_B1_valid(Tile_X01_Y03_SB_T1_EAST_SB_OUT_B1_valid),
		.SB_T1_NORTH_SB_IN_B1(Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_IN_B17(Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_IN_B17_ready(Tile_X01_Y03_SB_T1_NORTH_SB_IN_B17_ready),
		.SB_T1_NORTH_SB_IN_B17_valid(Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B17_valid),
		.SB_T1_NORTH_SB_IN_B1_ready(Tile_X01_Y03_SB_T1_NORTH_SB_IN_B1_ready),
		.SB_T1_NORTH_SB_IN_B1_valid(Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B1_valid),
		.SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_OUT_B17(Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_OUT_B17_ready(Tile_X01_Y02_SB_T1_SOUTH_SB_IN_B17_ready),
		.SB_T1_NORTH_SB_OUT_B17_valid(Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B17_valid),
		.SB_T1_NORTH_SB_OUT_B1_ready(Tile_X01_Y02_SB_T1_SOUTH_SB_IN_B1_ready),
		.SB_T1_NORTH_SB_OUT_B1_valid(Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B1_valid),
		.SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_IN_B17(Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_IN_B17_ready(Tile_X01_Y03_SB_T1_SOUTH_SB_IN_B17_ready),
		.SB_T1_SOUTH_SB_IN_B17_valid(Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B17_valid),
		.SB_T1_SOUTH_SB_IN_B1_ready(Tile_X01_Y03_SB_T1_SOUTH_SB_IN_B1_ready),
		.SB_T1_SOUTH_SB_IN_B1_valid(Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B1_valid),
		.SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_OUT_B17(Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_OUT_B17_ready(Tile_X01_Y04_SB_T1_NORTH_SB_IN_B17_ready),
		.SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B17_valid),
		.SB_T1_SOUTH_SB_OUT_B1_ready(Tile_X01_Y04_SB_T1_NORTH_SB_IN_B1_ready),
		.SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B1_valid),
		.SB_T1_WEST_SB_IN_B1(Tile_X00_Y03_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_WEST_SB_IN_B17(Tile_X00_Y03_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_WEST_SB_IN_B17_ready(Tile_X01_Y03_SB_T1_WEST_SB_IN_B17_ready),
		.SB_T1_WEST_SB_IN_B17_valid(Tile_X00_Y03_SB_T1_EAST_SB_OUT_B17_valid),
		.SB_T1_WEST_SB_IN_B1_ready(Tile_X01_Y03_SB_T1_WEST_SB_IN_B1_ready),
		.SB_T1_WEST_SB_IN_B1_valid(Tile_X00_Y03_SB_T1_EAST_SB_OUT_B1_valid),
		.SB_T1_WEST_SB_OUT_B1(Tile_X01_Y03_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_WEST_SB_OUT_B17(Tile_X01_Y03_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_WEST_SB_OUT_B17_ready(Tile_X00_Y03_SB_T1_EAST_SB_IN_B17_ready),
		.SB_T1_WEST_SB_OUT_B17_valid(Tile_X01_Y03_SB_T1_WEST_SB_OUT_B17_valid),
		.SB_T1_WEST_SB_OUT_B1_ready(Tile_X00_Y03_SB_T1_EAST_SB_IN_B1_ready),
		.SB_T1_WEST_SB_OUT_B1_valid(Tile_X01_Y03_SB_T1_WEST_SB_OUT_B1_valid),
		.SB_T2_EAST_SB_IN_B1(Tile_X02_Y03_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_EAST_SB_IN_B17(Tile_X02_Y03_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_EAST_SB_IN_B17_ready(Tile_X01_Y03_SB_T2_EAST_SB_IN_B17_ready),
		.SB_T2_EAST_SB_IN_B17_valid(Tile_X02_Y03_SB_T2_WEST_SB_OUT_B17_valid),
		.SB_T2_EAST_SB_IN_B1_ready(Tile_X01_Y03_SB_T2_EAST_SB_IN_B1_ready),
		.SB_T2_EAST_SB_IN_B1_valid(Tile_X02_Y03_SB_T2_WEST_SB_OUT_B1_valid),
		.SB_T2_EAST_SB_OUT_B1(Tile_X01_Y03_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_EAST_SB_OUT_B17(Tile_X01_Y03_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_EAST_SB_OUT_B17_ready(Tile_X02_Y03_SB_T2_WEST_SB_IN_B17_ready),
		.SB_T2_EAST_SB_OUT_B17_valid(Tile_X01_Y03_SB_T2_EAST_SB_OUT_B17_valid),
		.SB_T2_EAST_SB_OUT_B1_ready(Tile_X02_Y03_SB_T2_WEST_SB_IN_B1_ready),
		.SB_T2_EAST_SB_OUT_B1_valid(Tile_X01_Y03_SB_T2_EAST_SB_OUT_B1_valid),
		.SB_T2_NORTH_SB_IN_B1(Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_IN_B17(Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_IN_B17_ready(Tile_X01_Y03_SB_T2_NORTH_SB_IN_B17_ready),
		.SB_T2_NORTH_SB_IN_B17_valid(Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B17_valid),
		.SB_T2_NORTH_SB_IN_B1_ready(Tile_X01_Y03_SB_T2_NORTH_SB_IN_B1_ready),
		.SB_T2_NORTH_SB_IN_B1_valid(Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B1_valid),
		.SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_OUT_B17(Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_OUT_B17_ready(Tile_X01_Y02_SB_T2_SOUTH_SB_IN_B17_ready),
		.SB_T2_NORTH_SB_OUT_B17_valid(Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B17_valid),
		.SB_T2_NORTH_SB_OUT_B1_ready(Tile_X01_Y02_SB_T2_SOUTH_SB_IN_B1_ready),
		.SB_T2_NORTH_SB_OUT_B1_valid(Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B1_valid),
		.SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_IN_B17(Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_IN_B17_ready(Tile_X01_Y03_SB_T2_SOUTH_SB_IN_B17_ready),
		.SB_T2_SOUTH_SB_IN_B17_valid(Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B17_valid),
		.SB_T2_SOUTH_SB_IN_B1_ready(Tile_X01_Y03_SB_T2_SOUTH_SB_IN_B1_ready),
		.SB_T2_SOUTH_SB_IN_B1_valid(Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B1_valid),
		.SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_OUT_B17(Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_OUT_B17_ready(Tile_X01_Y04_SB_T2_NORTH_SB_IN_B17_ready),
		.SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B17_valid),
		.SB_T2_SOUTH_SB_OUT_B1_ready(Tile_X01_Y04_SB_T2_NORTH_SB_IN_B1_ready),
		.SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B1_valid),
		.SB_T2_WEST_SB_IN_B1(Tile_X00_Y03_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_WEST_SB_IN_B17(Tile_X00_Y03_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_WEST_SB_IN_B17_ready(Tile_X01_Y03_SB_T2_WEST_SB_IN_B17_ready),
		.SB_T2_WEST_SB_IN_B17_valid(Tile_X00_Y03_SB_T2_EAST_SB_OUT_B17_valid),
		.SB_T2_WEST_SB_IN_B1_ready(Tile_X01_Y03_SB_T2_WEST_SB_IN_B1_ready),
		.SB_T2_WEST_SB_IN_B1_valid(Tile_X00_Y03_SB_T2_EAST_SB_OUT_B1_valid),
		.SB_T2_WEST_SB_OUT_B1(Tile_X01_Y03_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_WEST_SB_OUT_B17(Tile_X01_Y03_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_WEST_SB_OUT_B17_ready(Tile_X00_Y03_SB_T2_EAST_SB_IN_B17_ready),
		.SB_T2_WEST_SB_OUT_B17_valid(Tile_X01_Y03_SB_T2_WEST_SB_OUT_B17_valid),
		.SB_T2_WEST_SB_OUT_B1_ready(Tile_X00_Y03_SB_T2_EAST_SB_IN_B1_ready),
		.SB_T2_WEST_SB_OUT_B1_valid(Tile_X01_Y03_SB_T2_WEST_SB_OUT_B1_valid),
		.SB_T3_EAST_SB_IN_B1(Tile_X02_Y03_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_EAST_SB_IN_B17(Tile_X02_Y03_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_EAST_SB_IN_B17_ready(Tile_X01_Y03_SB_T3_EAST_SB_IN_B17_ready),
		.SB_T3_EAST_SB_IN_B17_valid(Tile_X02_Y03_SB_T3_WEST_SB_OUT_B17_valid),
		.SB_T3_EAST_SB_IN_B1_ready(Tile_X01_Y03_SB_T3_EAST_SB_IN_B1_ready),
		.SB_T3_EAST_SB_IN_B1_valid(Tile_X02_Y03_SB_T3_WEST_SB_OUT_B1_valid),
		.SB_T3_EAST_SB_OUT_B1(Tile_X01_Y03_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_EAST_SB_OUT_B17(Tile_X01_Y03_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_EAST_SB_OUT_B17_ready(Tile_X02_Y03_SB_T3_WEST_SB_IN_B17_ready),
		.SB_T3_EAST_SB_OUT_B17_valid(Tile_X01_Y03_SB_T3_EAST_SB_OUT_B17_valid),
		.SB_T3_EAST_SB_OUT_B1_ready(Tile_X02_Y03_SB_T3_WEST_SB_IN_B1_ready),
		.SB_T3_EAST_SB_OUT_B1_valid(Tile_X01_Y03_SB_T3_EAST_SB_OUT_B1_valid),
		.SB_T3_NORTH_SB_IN_B1(Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_IN_B17(Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_IN_B17_ready(Tile_X01_Y03_SB_T3_NORTH_SB_IN_B17_ready),
		.SB_T3_NORTH_SB_IN_B17_valid(Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B17_valid),
		.SB_T3_NORTH_SB_IN_B1_ready(Tile_X01_Y03_SB_T3_NORTH_SB_IN_B1_ready),
		.SB_T3_NORTH_SB_IN_B1_valid(Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B1_valid),
		.SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_OUT_B17(Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_OUT_B17_ready(Tile_X01_Y02_SB_T3_SOUTH_SB_IN_B17_ready),
		.SB_T3_NORTH_SB_OUT_B17_valid(Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B17_valid),
		.SB_T3_NORTH_SB_OUT_B1_ready(Tile_X01_Y02_SB_T3_SOUTH_SB_IN_B1_ready),
		.SB_T3_NORTH_SB_OUT_B1_valid(Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B1_valid),
		.SB_T3_SOUTH_SB_IN_B1(Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_IN_B17(Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_IN_B17_ready(Tile_X01_Y03_SB_T3_SOUTH_SB_IN_B17_ready),
		.SB_T3_SOUTH_SB_IN_B17_valid(Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B17_valid),
		.SB_T3_SOUTH_SB_IN_B1_ready(Tile_X01_Y03_SB_T3_SOUTH_SB_IN_B1_ready),
		.SB_T3_SOUTH_SB_IN_B1_valid(Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B1_valid),
		.SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_OUT_B17(Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_OUT_B17_ready(Tile_X01_Y04_SB_T3_NORTH_SB_IN_B17_ready),
		.SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B17_valid),
		.SB_T3_SOUTH_SB_OUT_B1_ready(Tile_X01_Y04_SB_T3_NORTH_SB_IN_B1_ready),
		.SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B1_valid),
		.SB_T3_WEST_SB_IN_B1(Tile_X00_Y03_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_WEST_SB_IN_B17(Tile_X00_Y03_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_WEST_SB_IN_B17_ready(Tile_X01_Y03_SB_T3_WEST_SB_IN_B17_ready),
		.SB_T3_WEST_SB_IN_B17_valid(Tile_X00_Y03_SB_T3_EAST_SB_OUT_B17_valid),
		.SB_T3_WEST_SB_IN_B1_ready(Tile_X01_Y03_SB_T3_WEST_SB_IN_B1_ready),
		.SB_T3_WEST_SB_IN_B1_valid(Tile_X00_Y03_SB_T3_EAST_SB_OUT_B1_valid),
		.SB_T3_WEST_SB_OUT_B1(Tile_X01_Y03_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_WEST_SB_OUT_B17(Tile_X01_Y03_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_WEST_SB_OUT_B17_ready(Tile_X00_Y03_SB_T3_EAST_SB_IN_B17_ready),
		.SB_T3_WEST_SB_OUT_B17_valid(Tile_X01_Y03_SB_T3_WEST_SB_OUT_B17_valid),
		.SB_T3_WEST_SB_OUT_B1_ready(Tile_X00_Y03_SB_T3_EAST_SB_IN_B1_ready),
		.SB_T3_WEST_SB_OUT_B1_valid(Tile_X01_Y03_SB_T3_WEST_SB_OUT_B1_valid),
		.SB_T4_EAST_SB_IN_B1(Tile_X02_Y03_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_EAST_SB_IN_B17(Tile_X02_Y03_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_EAST_SB_IN_B17_ready(Tile_X01_Y03_SB_T4_EAST_SB_IN_B17_ready),
		.SB_T4_EAST_SB_IN_B17_valid(Tile_X02_Y03_SB_T4_WEST_SB_OUT_B17_valid),
		.SB_T4_EAST_SB_IN_B1_ready(Tile_X01_Y03_SB_T4_EAST_SB_IN_B1_ready),
		.SB_T4_EAST_SB_IN_B1_valid(Tile_X02_Y03_SB_T4_WEST_SB_OUT_B1_valid),
		.SB_T4_EAST_SB_OUT_B1(Tile_X01_Y03_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_EAST_SB_OUT_B17(Tile_X01_Y03_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_EAST_SB_OUT_B17_ready(Tile_X02_Y03_SB_T4_WEST_SB_IN_B17_ready),
		.SB_T4_EAST_SB_OUT_B17_valid(Tile_X01_Y03_SB_T4_EAST_SB_OUT_B17_valid),
		.SB_T4_EAST_SB_OUT_B1_ready(Tile_X02_Y03_SB_T4_WEST_SB_IN_B1_ready),
		.SB_T4_EAST_SB_OUT_B1_valid(Tile_X01_Y03_SB_T4_EAST_SB_OUT_B1_valid),
		.SB_T4_NORTH_SB_IN_B1(Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_IN_B17(Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_IN_B17_ready(Tile_X01_Y03_SB_T4_NORTH_SB_IN_B17_ready),
		.SB_T4_NORTH_SB_IN_B17_valid(Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B17_valid),
		.SB_T4_NORTH_SB_IN_B1_ready(Tile_X01_Y03_SB_T4_NORTH_SB_IN_B1_ready),
		.SB_T4_NORTH_SB_IN_B1_valid(Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B1_valid),
		.SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_OUT_B17(Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_OUT_B17_ready(Tile_X01_Y02_SB_T4_SOUTH_SB_IN_B17_ready),
		.SB_T4_NORTH_SB_OUT_B17_valid(Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B17_valid),
		.SB_T4_NORTH_SB_OUT_B1_ready(Tile_X01_Y02_SB_T4_SOUTH_SB_IN_B1_ready),
		.SB_T4_NORTH_SB_OUT_B1_valid(Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B1_valid),
		.SB_T4_SOUTH_SB_IN_B1(Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_IN_B17(Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_IN_B17_ready(Tile_X01_Y03_SB_T4_SOUTH_SB_IN_B17_ready),
		.SB_T4_SOUTH_SB_IN_B17_valid(Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B17_valid),
		.SB_T4_SOUTH_SB_IN_B1_ready(Tile_X01_Y03_SB_T4_SOUTH_SB_IN_B1_ready),
		.SB_T4_SOUTH_SB_IN_B1_valid(Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B1_valid),
		.SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_OUT_B17(Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_OUT_B17_ready(Tile_X01_Y04_SB_T4_NORTH_SB_IN_B17_ready),
		.SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B17_valid),
		.SB_T4_SOUTH_SB_OUT_B1_ready(Tile_X01_Y04_SB_T4_NORTH_SB_IN_B1_ready),
		.SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B1_valid),
		.SB_T4_WEST_SB_IN_B1(Tile_X00_Y03_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_WEST_SB_IN_B17(Tile_X00_Y03_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_WEST_SB_IN_B17_ready(Tile_X01_Y03_SB_T4_WEST_SB_IN_B17_ready),
		.SB_T4_WEST_SB_IN_B17_valid(Tile_X00_Y03_SB_T4_EAST_SB_OUT_B17_valid),
		.SB_T4_WEST_SB_IN_B1_ready(Tile_X01_Y03_SB_T4_WEST_SB_IN_B1_ready),
		.SB_T4_WEST_SB_IN_B1_valid(Tile_X00_Y03_SB_T4_EAST_SB_OUT_B1_valid),
		.SB_T4_WEST_SB_OUT_B1(Tile_X01_Y03_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_WEST_SB_OUT_B17(Tile_X01_Y03_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_WEST_SB_OUT_B17_ready(Tile_X00_Y03_SB_T4_EAST_SB_IN_B17_ready),
		.SB_T4_WEST_SB_OUT_B17_valid(Tile_X01_Y03_SB_T4_WEST_SB_OUT_B17_valid),
		.SB_T4_WEST_SB_OUT_B1_ready(Tile_X00_Y03_SB_T4_EAST_SB_IN_B1_ready),
		.SB_T4_WEST_SB_OUT_B1_valid(Tile_X01_Y03_SB_T4_WEST_SB_OUT_B1_valid),
		.clk(Tile_X01_Y02_clk_out),
		.clk_out(Tile_X01_Y03_clk_out),
		.clk_pass_through(Tile_X01_Y02_clk_pass_through_out_bot),
		.clk_pass_through_out_bot(Tile_X01_Y03_clk_pass_through_out_bot),
		.clk_pass_through_out_right(Tile_X01_Y03_clk_pass_through_out_right),
		.config_config_addr(Tile_X01_Y02_config_out_config_addr),
		.config_config_data(Tile_X01_Y02_config_out_config_data),
		.config_out_config_addr(Tile_X01_Y03_config_out_config_addr),
		.config_out_config_data(Tile_X01_Y03_config_out_config_data),
		.config_out_read(Tile_X01_Y03_config_out_read),
		.config_out_write(Tile_X01_Y03_config_out_write),
		.config_read(Tile_X01_Y02_config_out_read),
		.config_write(Tile_X01_Y02_config_out_write),
		.flush(Tile_X01_Y02_flush_out),
		.flush_out(Tile_X01_Y03_flush_out),
		.hi(Tile_X01_Y03_hi),
		.lo(Tile_X01_Y03_lo),
		.read_config_data(Tile_X01_Y03_read_config_data),
		.read_config_data_in(Tile_X01_Y02_read_config_data),
		.reset(Tile_X01_Y02_reset_out),
		.reset_out(Tile_X01_Y03_reset_out),
		.stall(Tile_X01_Y02_stall_out),
		.stall_out(Tile_X01_Y03_stall_out),
		.tile_id(Tile_X01_Y03_tile_id)
	);
	wire [15:0] Tile_X01_Y04_tile_id;
	assign Tile_X01_Y04_tile_id = {Tile_X01_Y04_lo[7], Tile_X01_Y04_lo[7], Tile_X01_Y04_lo[6], Tile_X01_Y04_lo[6], Tile_X01_Y04_lo[5], Tile_X01_Y04_lo[5], Tile_X01_Y04_lo[4], Tile_X01_Y04_hi[4], Tile_X01_Y04_lo[3], Tile_X01_Y04_lo[3], Tile_X01_Y04_lo[2], Tile_X01_Y04_lo[2], Tile_X01_Y04_lo[1], Tile_X01_Y04_hi[1], Tile_X01_Y04_lo[0], Tile_X01_Y04_lo[0]};
	Tile_PE Tile_X01_Y04(
		.SB_T0_EAST_SB_IN_B1(Tile_X02_Y04_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_EAST_SB_IN_B17(Tile_X02_Y04_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_EAST_SB_IN_B17_ready(Tile_X01_Y04_SB_T0_EAST_SB_IN_B17_ready),
		.SB_T0_EAST_SB_IN_B17_valid(Tile_X02_Y04_SB_T0_WEST_SB_OUT_B17_valid),
		.SB_T0_EAST_SB_IN_B1_ready(Tile_X01_Y04_SB_T0_EAST_SB_IN_B1_ready),
		.SB_T0_EAST_SB_IN_B1_valid(Tile_X02_Y04_SB_T0_WEST_SB_OUT_B1_valid),
		.SB_T0_EAST_SB_OUT_B1(Tile_X01_Y04_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_EAST_SB_OUT_B17(Tile_X01_Y04_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_EAST_SB_OUT_B17_ready(Tile_X02_Y04_SB_T0_WEST_SB_IN_B17_ready),
		.SB_T0_EAST_SB_OUT_B17_valid(Tile_X01_Y04_SB_T0_EAST_SB_OUT_B17_valid),
		.SB_T0_EAST_SB_OUT_B1_ready(Tile_X02_Y04_SB_T0_WEST_SB_IN_B1_ready),
		.SB_T0_EAST_SB_OUT_B1_valid(Tile_X01_Y04_SB_T0_EAST_SB_OUT_B1_valid),
		.SB_T0_NORTH_SB_IN_B1(Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_IN_B17(Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_IN_B17_ready(Tile_X01_Y04_SB_T0_NORTH_SB_IN_B17_ready),
		.SB_T0_NORTH_SB_IN_B17_valid(Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B17_valid),
		.SB_T0_NORTH_SB_IN_B1_ready(Tile_X01_Y04_SB_T0_NORTH_SB_IN_B1_ready),
		.SB_T0_NORTH_SB_IN_B1_valid(Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B1_valid),
		.SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_OUT_B17(Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_OUT_B17_ready(Tile_X01_Y03_SB_T0_SOUTH_SB_IN_B17_ready),
		.SB_T0_NORTH_SB_OUT_B17_valid(Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B17_valid),
		.SB_T0_NORTH_SB_OUT_B1_ready(Tile_X01_Y03_SB_T0_SOUTH_SB_IN_B1_ready),
		.SB_T0_NORTH_SB_OUT_B1_valid(Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B1_valid),
		.SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
		.SB_T0_SOUTH_SB_IN_B17(const_0_17_out),
		.SB_T0_SOUTH_SB_IN_B17_ready(Tile_X01_Y04_SB_T0_SOUTH_SB_IN_B17_ready),
		.SB_T0_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T0_SOUTH_SB_IN_B1_ready(Tile_X01_Y04_SB_T0_SOUTH_SB_IN_B1_ready),
		.SB_T0_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_OUT_B17(Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B17_valid),
		.SB_T0_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B1_valid),
		.SB_T0_WEST_SB_IN_B1(Tile_X00_Y04_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_WEST_SB_IN_B17(Tile_X00_Y04_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_WEST_SB_IN_B17_ready(Tile_X01_Y04_SB_T0_WEST_SB_IN_B17_ready),
		.SB_T0_WEST_SB_IN_B17_valid(Tile_X00_Y04_SB_T0_EAST_SB_OUT_B17_valid),
		.SB_T0_WEST_SB_IN_B1_ready(Tile_X01_Y04_SB_T0_WEST_SB_IN_B1_ready),
		.SB_T0_WEST_SB_IN_B1_valid(Tile_X00_Y04_SB_T0_EAST_SB_OUT_B1_valid),
		.SB_T0_WEST_SB_OUT_B1(Tile_X01_Y04_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_WEST_SB_OUT_B17(Tile_X01_Y04_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_WEST_SB_OUT_B17_ready(Tile_X00_Y04_SB_T0_EAST_SB_IN_B17_ready),
		.SB_T0_WEST_SB_OUT_B17_valid(Tile_X01_Y04_SB_T0_WEST_SB_OUT_B17_valid),
		.SB_T0_WEST_SB_OUT_B1_ready(Tile_X00_Y04_SB_T0_EAST_SB_IN_B1_ready),
		.SB_T0_WEST_SB_OUT_B1_valid(Tile_X01_Y04_SB_T0_WEST_SB_OUT_B1_valid),
		.SB_T1_EAST_SB_IN_B1(Tile_X02_Y04_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_EAST_SB_IN_B17(Tile_X02_Y04_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_EAST_SB_IN_B17_ready(Tile_X01_Y04_SB_T1_EAST_SB_IN_B17_ready),
		.SB_T1_EAST_SB_IN_B17_valid(Tile_X02_Y04_SB_T1_WEST_SB_OUT_B17_valid),
		.SB_T1_EAST_SB_IN_B1_ready(Tile_X01_Y04_SB_T1_EAST_SB_IN_B1_ready),
		.SB_T1_EAST_SB_IN_B1_valid(Tile_X02_Y04_SB_T1_WEST_SB_OUT_B1_valid),
		.SB_T1_EAST_SB_OUT_B1(Tile_X01_Y04_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_EAST_SB_OUT_B17(Tile_X01_Y04_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_EAST_SB_OUT_B17_ready(Tile_X02_Y04_SB_T1_WEST_SB_IN_B17_ready),
		.SB_T1_EAST_SB_OUT_B17_valid(Tile_X01_Y04_SB_T1_EAST_SB_OUT_B17_valid),
		.SB_T1_EAST_SB_OUT_B1_ready(Tile_X02_Y04_SB_T1_WEST_SB_IN_B1_ready),
		.SB_T1_EAST_SB_OUT_B1_valid(Tile_X01_Y04_SB_T1_EAST_SB_OUT_B1_valid),
		.SB_T1_NORTH_SB_IN_B1(Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_IN_B17(Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_IN_B17_ready(Tile_X01_Y04_SB_T1_NORTH_SB_IN_B17_ready),
		.SB_T1_NORTH_SB_IN_B17_valid(Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B17_valid),
		.SB_T1_NORTH_SB_IN_B1_ready(Tile_X01_Y04_SB_T1_NORTH_SB_IN_B1_ready),
		.SB_T1_NORTH_SB_IN_B1_valid(Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B1_valid),
		.SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_OUT_B17(Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_OUT_B17_ready(Tile_X01_Y03_SB_T1_SOUTH_SB_IN_B17_ready),
		.SB_T1_NORTH_SB_OUT_B17_valid(Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B17_valid),
		.SB_T1_NORTH_SB_OUT_B1_ready(Tile_X01_Y03_SB_T1_SOUTH_SB_IN_B1_ready),
		.SB_T1_NORTH_SB_OUT_B1_valid(Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B1_valid),
		.SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
		.SB_T1_SOUTH_SB_IN_B17(const_0_17_out),
		.SB_T1_SOUTH_SB_IN_B17_ready(Tile_X01_Y04_SB_T1_SOUTH_SB_IN_B17_ready),
		.SB_T1_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T1_SOUTH_SB_IN_B1_ready(Tile_X01_Y04_SB_T1_SOUTH_SB_IN_B1_ready),
		.SB_T1_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_OUT_B17(Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B17_valid),
		.SB_T1_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B1_valid),
		.SB_T1_WEST_SB_IN_B1(Tile_X00_Y04_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_WEST_SB_IN_B17(Tile_X00_Y04_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_WEST_SB_IN_B17_ready(Tile_X01_Y04_SB_T1_WEST_SB_IN_B17_ready),
		.SB_T1_WEST_SB_IN_B17_valid(Tile_X00_Y04_SB_T1_EAST_SB_OUT_B17_valid),
		.SB_T1_WEST_SB_IN_B1_ready(Tile_X01_Y04_SB_T1_WEST_SB_IN_B1_ready),
		.SB_T1_WEST_SB_IN_B1_valid(Tile_X00_Y04_SB_T1_EAST_SB_OUT_B1_valid),
		.SB_T1_WEST_SB_OUT_B1(Tile_X01_Y04_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_WEST_SB_OUT_B17(Tile_X01_Y04_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_WEST_SB_OUT_B17_ready(Tile_X00_Y04_SB_T1_EAST_SB_IN_B17_ready),
		.SB_T1_WEST_SB_OUT_B17_valid(Tile_X01_Y04_SB_T1_WEST_SB_OUT_B17_valid),
		.SB_T1_WEST_SB_OUT_B1_ready(Tile_X00_Y04_SB_T1_EAST_SB_IN_B1_ready),
		.SB_T1_WEST_SB_OUT_B1_valid(Tile_X01_Y04_SB_T1_WEST_SB_OUT_B1_valid),
		.SB_T2_EAST_SB_IN_B1(Tile_X02_Y04_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_EAST_SB_IN_B17(Tile_X02_Y04_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_EAST_SB_IN_B17_ready(Tile_X01_Y04_SB_T2_EAST_SB_IN_B17_ready),
		.SB_T2_EAST_SB_IN_B17_valid(Tile_X02_Y04_SB_T2_WEST_SB_OUT_B17_valid),
		.SB_T2_EAST_SB_IN_B1_ready(Tile_X01_Y04_SB_T2_EAST_SB_IN_B1_ready),
		.SB_T2_EAST_SB_IN_B1_valid(Tile_X02_Y04_SB_T2_WEST_SB_OUT_B1_valid),
		.SB_T2_EAST_SB_OUT_B1(Tile_X01_Y04_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_EAST_SB_OUT_B17(Tile_X01_Y04_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_EAST_SB_OUT_B17_ready(Tile_X02_Y04_SB_T2_WEST_SB_IN_B17_ready),
		.SB_T2_EAST_SB_OUT_B17_valid(Tile_X01_Y04_SB_T2_EAST_SB_OUT_B17_valid),
		.SB_T2_EAST_SB_OUT_B1_ready(Tile_X02_Y04_SB_T2_WEST_SB_IN_B1_ready),
		.SB_T2_EAST_SB_OUT_B1_valid(Tile_X01_Y04_SB_T2_EAST_SB_OUT_B1_valid),
		.SB_T2_NORTH_SB_IN_B1(Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_IN_B17(Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_IN_B17_ready(Tile_X01_Y04_SB_T2_NORTH_SB_IN_B17_ready),
		.SB_T2_NORTH_SB_IN_B17_valid(Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B17_valid),
		.SB_T2_NORTH_SB_IN_B1_ready(Tile_X01_Y04_SB_T2_NORTH_SB_IN_B1_ready),
		.SB_T2_NORTH_SB_IN_B1_valid(Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B1_valid),
		.SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_OUT_B17(Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_OUT_B17_ready(Tile_X01_Y03_SB_T2_SOUTH_SB_IN_B17_ready),
		.SB_T2_NORTH_SB_OUT_B17_valid(Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B17_valid),
		.SB_T2_NORTH_SB_OUT_B1_ready(Tile_X01_Y03_SB_T2_SOUTH_SB_IN_B1_ready),
		.SB_T2_NORTH_SB_OUT_B1_valid(Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B1_valid),
		.SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
		.SB_T2_SOUTH_SB_IN_B17(const_0_17_out),
		.SB_T2_SOUTH_SB_IN_B17_ready(Tile_X01_Y04_SB_T2_SOUTH_SB_IN_B17_ready),
		.SB_T2_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T2_SOUTH_SB_IN_B1_ready(Tile_X01_Y04_SB_T2_SOUTH_SB_IN_B1_ready),
		.SB_T2_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_OUT_B17(Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B17_valid),
		.SB_T2_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B1_valid),
		.SB_T2_WEST_SB_IN_B1(Tile_X00_Y04_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_WEST_SB_IN_B17(Tile_X00_Y04_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_WEST_SB_IN_B17_ready(Tile_X01_Y04_SB_T2_WEST_SB_IN_B17_ready),
		.SB_T2_WEST_SB_IN_B17_valid(Tile_X00_Y04_SB_T2_EAST_SB_OUT_B17_valid),
		.SB_T2_WEST_SB_IN_B1_ready(Tile_X01_Y04_SB_T2_WEST_SB_IN_B1_ready),
		.SB_T2_WEST_SB_IN_B1_valid(Tile_X00_Y04_SB_T2_EAST_SB_OUT_B1_valid),
		.SB_T2_WEST_SB_OUT_B1(Tile_X01_Y04_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_WEST_SB_OUT_B17(Tile_X01_Y04_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_WEST_SB_OUT_B17_ready(Tile_X00_Y04_SB_T2_EAST_SB_IN_B17_ready),
		.SB_T2_WEST_SB_OUT_B17_valid(Tile_X01_Y04_SB_T2_WEST_SB_OUT_B17_valid),
		.SB_T2_WEST_SB_OUT_B1_ready(Tile_X00_Y04_SB_T2_EAST_SB_IN_B1_ready),
		.SB_T2_WEST_SB_OUT_B1_valid(Tile_X01_Y04_SB_T2_WEST_SB_OUT_B1_valid),
		.SB_T3_EAST_SB_IN_B1(Tile_X02_Y04_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_EAST_SB_IN_B17(Tile_X02_Y04_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_EAST_SB_IN_B17_ready(Tile_X01_Y04_SB_T3_EAST_SB_IN_B17_ready),
		.SB_T3_EAST_SB_IN_B17_valid(Tile_X02_Y04_SB_T3_WEST_SB_OUT_B17_valid),
		.SB_T3_EAST_SB_IN_B1_ready(Tile_X01_Y04_SB_T3_EAST_SB_IN_B1_ready),
		.SB_T3_EAST_SB_IN_B1_valid(Tile_X02_Y04_SB_T3_WEST_SB_OUT_B1_valid),
		.SB_T3_EAST_SB_OUT_B1(Tile_X01_Y04_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_EAST_SB_OUT_B17(Tile_X01_Y04_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_EAST_SB_OUT_B17_ready(Tile_X02_Y04_SB_T3_WEST_SB_IN_B17_ready),
		.SB_T3_EAST_SB_OUT_B17_valid(Tile_X01_Y04_SB_T3_EAST_SB_OUT_B17_valid),
		.SB_T3_EAST_SB_OUT_B1_ready(Tile_X02_Y04_SB_T3_WEST_SB_IN_B1_ready),
		.SB_T3_EAST_SB_OUT_B1_valid(Tile_X01_Y04_SB_T3_EAST_SB_OUT_B1_valid),
		.SB_T3_NORTH_SB_IN_B1(Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_IN_B17(Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_IN_B17_ready(Tile_X01_Y04_SB_T3_NORTH_SB_IN_B17_ready),
		.SB_T3_NORTH_SB_IN_B17_valid(Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B17_valid),
		.SB_T3_NORTH_SB_IN_B1_ready(Tile_X01_Y04_SB_T3_NORTH_SB_IN_B1_ready),
		.SB_T3_NORTH_SB_IN_B1_valid(Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B1_valid),
		.SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_OUT_B17(Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_OUT_B17_ready(Tile_X01_Y03_SB_T3_SOUTH_SB_IN_B17_ready),
		.SB_T3_NORTH_SB_OUT_B17_valid(Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B17_valid),
		.SB_T3_NORTH_SB_OUT_B1_ready(Tile_X01_Y03_SB_T3_SOUTH_SB_IN_B1_ready),
		.SB_T3_NORTH_SB_OUT_B1_valid(Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B1_valid),
		.SB_T3_SOUTH_SB_IN_B1(const_0_1_out),
		.SB_T3_SOUTH_SB_IN_B17(const_0_17_out),
		.SB_T3_SOUTH_SB_IN_B17_ready(Tile_X01_Y04_SB_T3_SOUTH_SB_IN_B17_ready),
		.SB_T3_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T3_SOUTH_SB_IN_B1_ready(Tile_X01_Y04_SB_T3_SOUTH_SB_IN_B1_ready),
		.SB_T3_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y04_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_OUT_B17(Tile_X01_Y04_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X01_Y04_SB_T3_SOUTH_SB_OUT_B17_valid),
		.SB_T3_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X01_Y04_SB_T3_SOUTH_SB_OUT_B1_valid),
		.SB_T3_WEST_SB_IN_B1(Tile_X00_Y04_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_WEST_SB_IN_B17(Tile_X00_Y04_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_WEST_SB_IN_B17_ready(Tile_X01_Y04_SB_T3_WEST_SB_IN_B17_ready),
		.SB_T3_WEST_SB_IN_B17_valid(Tile_X00_Y04_SB_T3_EAST_SB_OUT_B17_valid),
		.SB_T3_WEST_SB_IN_B1_ready(Tile_X01_Y04_SB_T3_WEST_SB_IN_B1_ready),
		.SB_T3_WEST_SB_IN_B1_valid(Tile_X00_Y04_SB_T3_EAST_SB_OUT_B1_valid),
		.SB_T3_WEST_SB_OUT_B1(Tile_X01_Y04_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_WEST_SB_OUT_B17(Tile_X01_Y04_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_WEST_SB_OUT_B17_ready(Tile_X00_Y04_SB_T3_EAST_SB_IN_B17_ready),
		.SB_T3_WEST_SB_OUT_B17_valid(Tile_X01_Y04_SB_T3_WEST_SB_OUT_B17_valid),
		.SB_T3_WEST_SB_OUT_B1_ready(Tile_X00_Y04_SB_T3_EAST_SB_IN_B1_ready),
		.SB_T3_WEST_SB_OUT_B1_valid(Tile_X01_Y04_SB_T3_WEST_SB_OUT_B1_valid),
		.SB_T4_EAST_SB_IN_B1(Tile_X02_Y04_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_EAST_SB_IN_B17(Tile_X02_Y04_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_EAST_SB_IN_B17_ready(Tile_X01_Y04_SB_T4_EAST_SB_IN_B17_ready),
		.SB_T4_EAST_SB_IN_B17_valid(Tile_X02_Y04_SB_T4_WEST_SB_OUT_B17_valid),
		.SB_T4_EAST_SB_IN_B1_ready(Tile_X01_Y04_SB_T4_EAST_SB_IN_B1_ready),
		.SB_T4_EAST_SB_IN_B1_valid(Tile_X02_Y04_SB_T4_WEST_SB_OUT_B1_valid),
		.SB_T4_EAST_SB_OUT_B1(Tile_X01_Y04_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_EAST_SB_OUT_B17(Tile_X01_Y04_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_EAST_SB_OUT_B17_ready(Tile_X02_Y04_SB_T4_WEST_SB_IN_B17_ready),
		.SB_T4_EAST_SB_OUT_B17_valid(Tile_X01_Y04_SB_T4_EAST_SB_OUT_B17_valid),
		.SB_T4_EAST_SB_OUT_B1_ready(Tile_X02_Y04_SB_T4_WEST_SB_IN_B1_ready),
		.SB_T4_EAST_SB_OUT_B1_valid(Tile_X01_Y04_SB_T4_EAST_SB_OUT_B1_valid),
		.SB_T4_NORTH_SB_IN_B1(Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_IN_B17(Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_IN_B17_ready(Tile_X01_Y04_SB_T4_NORTH_SB_IN_B17_ready),
		.SB_T4_NORTH_SB_IN_B17_valid(Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B17_valid),
		.SB_T4_NORTH_SB_IN_B1_ready(Tile_X01_Y04_SB_T4_NORTH_SB_IN_B1_ready),
		.SB_T4_NORTH_SB_IN_B1_valid(Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B1_valid),
		.SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_OUT_B17(Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_OUT_B17_ready(Tile_X01_Y03_SB_T4_SOUTH_SB_IN_B17_ready),
		.SB_T4_NORTH_SB_OUT_B17_valid(Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B17_valid),
		.SB_T4_NORTH_SB_OUT_B1_ready(Tile_X01_Y03_SB_T4_SOUTH_SB_IN_B1_ready),
		.SB_T4_NORTH_SB_OUT_B1_valid(Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B1_valid),
		.SB_T4_SOUTH_SB_IN_B1(const_0_1_out),
		.SB_T4_SOUTH_SB_IN_B17(const_0_17_out),
		.SB_T4_SOUTH_SB_IN_B17_ready(Tile_X01_Y04_SB_T4_SOUTH_SB_IN_B17_ready),
		.SB_T4_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T4_SOUTH_SB_IN_B1_ready(Tile_X01_Y04_SB_T4_SOUTH_SB_IN_B1_ready),
		.SB_T4_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y04_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_OUT_B17(Tile_X01_Y04_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X01_Y04_SB_T4_SOUTH_SB_OUT_B17_valid),
		.SB_T4_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X01_Y04_SB_T4_SOUTH_SB_OUT_B1_valid),
		.SB_T4_WEST_SB_IN_B1(Tile_X00_Y04_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_WEST_SB_IN_B17(Tile_X00_Y04_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_WEST_SB_IN_B17_ready(Tile_X01_Y04_SB_T4_WEST_SB_IN_B17_ready),
		.SB_T4_WEST_SB_IN_B17_valid(Tile_X00_Y04_SB_T4_EAST_SB_OUT_B17_valid),
		.SB_T4_WEST_SB_IN_B1_ready(Tile_X01_Y04_SB_T4_WEST_SB_IN_B1_ready),
		.SB_T4_WEST_SB_IN_B1_valid(Tile_X00_Y04_SB_T4_EAST_SB_OUT_B1_valid),
		.SB_T4_WEST_SB_OUT_B1(Tile_X01_Y04_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_WEST_SB_OUT_B17(Tile_X01_Y04_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_WEST_SB_OUT_B17_ready(Tile_X00_Y04_SB_T4_EAST_SB_IN_B17_ready),
		.SB_T4_WEST_SB_OUT_B17_valid(Tile_X01_Y04_SB_T4_WEST_SB_OUT_B17_valid),
		.SB_T4_WEST_SB_OUT_B1_ready(Tile_X00_Y04_SB_T4_EAST_SB_IN_B1_ready),
		.SB_T4_WEST_SB_OUT_B1_valid(Tile_X01_Y04_SB_T4_WEST_SB_OUT_B1_valid),
		.clk(Tile_X01_Y03_clk_out),
		.clk_out(Tile_X01_Y04_clk_out),
		.clk_pass_through(Tile_X01_Y03_clk_pass_through_out_bot),
		.clk_pass_through_out_bot(Tile_X01_Y04_clk_pass_through_out_bot),
		.clk_pass_through_out_right(Tile_X01_Y04_clk_pass_through_out_right),
		.config_config_addr(Tile_X01_Y03_config_out_config_addr),
		.config_config_data(Tile_X01_Y03_config_out_config_data),
		.config_out_config_addr(Tile_X01_Y04_config_out_config_addr),
		.config_out_config_data(Tile_X01_Y04_config_out_config_data),
		.config_out_read(Tile_X01_Y04_config_out_read),
		.config_out_write(Tile_X01_Y04_config_out_write),
		.config_read(Tile_X01_Y03_config_out_read),
		.config_write(Tile_X01_Y03_config_out_write),
		.flush(Tile_X01_Y03_flush_out),
		.flush_out(Tile_X01_Y04_flush_out),
		.hi(Tile_X01_Y04_hi),
		.lo(Tile_X01_Y04_lo),
		.read_config_data(Tile_X01_Y04_read_config_data),
		.read_config_data_in(Tile_X01_Y03_read_config_data),
		.reset(Tile_X01_Y03_reset_out),
		.reset_out(Tile_X01_Y04_reset_out),
		.stall(Tile_X01_Y03_stall_out),
		.stall_out(Tile_X01_Y04_stall_out),
		.tile_id(Tile_X01_Y04_tile_id)
	);
	wire [31:0] Tile_X02_Y00_config_config_addr;
	assign Tile_X02_Y00_config_config_addr = {PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[31], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[30], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[29], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[28], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[27], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[26], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[25], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[24], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[23], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[22], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[21], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[20], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[19], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[18], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[17], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[16], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[15], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[14], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[13], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[12], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[11], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[10], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[9], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[8], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[7], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[6], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[5], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[4], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[3], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[2], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[1], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[0]};
	wire [31:0] Tile_X02_Y00_config_config_data;
	assign Tile_X02_Y00_config_config_data = {PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[63], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[62], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[61], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[60], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[59], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[58], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[57], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[56], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[55], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[54], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[53], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[52], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[51], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[50], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[49], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[48], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[47], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[46], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[45], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[44], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[43], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[42], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[41], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[40], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[39], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[38], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[37], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[36], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[35], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[34], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[33], PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[32]};
	wire [4:0] Tile_X02_Y00_io2f_17_ready;
	assign Tile_X02_Y00_io2f_17_ready = {Tile_X02_Y01_SB_T4_NORTH_SB_IN_B17_ready, Tile_X02_Y01_SB_T3_NORTH_SB_IN_B17_ready, Tile_X02_Y01_SB_T2_NORTH_SB_IN_B17_ready, Tile_X02_Y01_SB_T1_NORTH_SB_IN_B17_ready, Tile_X02_Y01_SB_T0_NORTH_SB_IN_B17_ready};
	wire [4:0] Tile_X02_Y00_io2f_1_ready;
	assign Tile_X02_Y00_io2f_1_ready = {Tile_X02_Y01_SB_T4_NORTH_SB_IN_B1_ready, Tile_X02_Y01_SB_T3_NORTH_SB_IN_B1_ready, Tile_X02_Y01_SB_T2_NORTH_SB_IN_B1_ready, Tile_X02_Y01_SB_T1_NORTH_SB_IN_B1_ready, Tile_X02_Y01_SB_T0_NORTH_SB_IN_B1_ready};
	wire [15:0] Tile_X02_Y00_tile_id;
	assign Tile_X02_Y00_tile_id = {Tile_X02_Y00_lo[7], Tile_X02_Y00_lo[7], Tile_X02_Y00_lo[6], Tile_X02_Y00_lo[6], Tile_X02_Y00_lo[5], Tile_X02_Y00_lo[5], Tile_X02_Y00_hi[5], Tile_X02_Y00_lo[4], Tile_X02_Y00_lo[3], Tile_X02_Y00_lo[3], Tile_X02_Y00_lo[2], Tile_X02_Y00_lo[2], Tile_X02_Y00_lo[1], Tile_X02_Y00_lo[1], Tile_X02_Y00_lo[0], Tile_X02_Y00_lo[0]};
	Tile_IOCoreReadyValid Tile_X02_Y00(
		.clk(clk),
		.clk_out(Tile_X02_Y00_clk_out),
		.config_config_addr(Tile_X02_Y00_config_config_addr),
		.config_config_data(Tile_X02_Y00_config_config_data),
		.config_out_config_addr(Tile_X02_Y00_config_out_config_addr),
		.config_out_config_data(Tile_X02_Y00_config_out_config_data),
		.config_out_read(Tile_X02_Y00_config_out_read),
		.config_out_write(Tile_X02_Y00_config_out_write),
		.config_read(PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[64]),
		.config_write(PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[65]),
		.f2io_1(Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B1),
		.f2io_17(Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B17),
		.f2io_17_ready(Tile_X02_Y00_f2io_17_ready),
		.f2io_17_valid(Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B17_valid),
		.f2io_1_ready(Tile_X02_Y00_f2io_1_ready),
		.f2io_1_valid(Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B1_valid),
		.flush(PipelineRegister_inst2$Register_inst0$reg_P1_inst0_out),
		.flush_out(Tile_X02_Y00_flush_out),
		.glb2io_1(glb2io_1_X02_Y00),
		.glb2io_17(glb2io_17_X02_Y00),
		.glb2io_17_ready(Tile_X02_Y00_glb2io_17_ready),
		.glb2io_17_valid(glb2io_17_X02_Y00_valid),
		.glb2io_1_ready(Tile_X02_Y00_glb2io_1_ready),
		.glb2io_1_valid(glb2io_1_X02_Y00_valid),
		.hi(Tile_X02_Y00_hi),
		.io2f_1(Tile_X02_Y00_io2f_1),
		.io2f_17(Tile_X02_Y00_io2f_17),
		.io2f_17_ready(Tile_X02_Y00_io2f_17_ready),
		.io2f_17_valid(Tile_X02_Y00_io2f_17_valid),
		.io2f_1_ready(Tile_X02_Y00_io2f_1_ready),
		.io2f_1_valid(Tile_X02_Y00_io2f_1_valid),
		.io2glb_1(Tile_X02_Y00_io2glb_1),
		.io2glb_17(Tile_X02_Y00_io2glb_17),
		.io2glb_17_ready(io2glb_17_X02_Y00_ready),
		.io2glb_17_valid(Tile_X02_Y00_io2glb_17_valid),
		.io2glb_1_ready(io2glb_1_X02_Y00_ready),
		.io2glb_1_valid(Tile_X02_Y00_io2glb_1_valid),
		.lo(Tile_X02_Y00_lo),
		.read_config_data(Tile_X02_Y00_read_config_data),
		.read_config_data_in(const_0_32_out),
		.reset(reset),
		.reset_out(Tile_X02_Y00_reset_out),
		.stall(self_stall_out[2:2]),
		.stall_out(Tile_X02_Y00_stall_out),
		.tile_id(Tile_X02_Y00_tile_id)
	);
	wire [15:0] Tile_X02_Y01_tile_id;
	assign Tile_X02_Y01_tile_id = {Tile_X02_Y01_lo[7], Tile_X02_Y01_lo[7], Tile_X02_Y01_lo[6], Tile_X02_Y01_lo[6], Tile_X02_Y01_lo[5], Tile_X02_Y01_lo[5], Tile_X02_Y01_hi[5], Tile_X02_Y01_lo[4], Tile_X02_Y01_lo[3], Tile_X02_Y01_lo[3], Tile_X02_Y01_lo[2], Tile_X02_Y01_lo[2], Tile_X02_Y01_lo[1], Tile_X02_Y01_lo[1], Tile_X02_Y01_lo[0], Tile_X02_Y01_hi[0]};
	Tile_PE Tile_X02_Y01(
		.SB_T0_EAST_SB_IN_B1(Tile_X03_Y01_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_EAST_SB_IN_B17(Tile_X03_Y01_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_EAST_SB_IN_B17_ready(Tile_X02_Y01_SB_T0_EAST_SB_IN_B17_ready),
		.SB_T0_EAST_SB_IN_B17_valid(Tile_X03_Y01_SB_T0_WEST_SB_OUT_B17_valid),
		.SB_T0_EAST_SB_IN_B1_ready(Tile_X02_Y01_SB_T0_EAST_SB_IN_B1_ready),
		.SB_T0_EAST_SB_IN_B1_valid(Tile_X03_Y01_SB_T0_WEST_SB_OUT_B1_valid),
		.SB_T0_EAST_SB_OUT_B1(Tile_X02_Y01_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_EAST_SB_OUT_B17(Tile_X02_Y01_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_EAST_SB_OUT_B17_ready(Tile_X03_Y01_SB_T0_WEST_SB_IN_B17_ready),
		.SB_T0_EAST_SB_OUT_B17_valid(Tile_X02_Y01_SB_T0_EAST_SB_OUT_B17_valid),
		.SB_T0_EAST_SB_OUT_B1_ready(Tile_X03_Y01_SB_T0_WEST_SB_IN_B1_ready),
		.SB_T0_EAST_SB_OUT_B1_valid(Tile_X02_Y01_SB_T0_EAST_SB_OUT_B1_valid),
		.SB_T0_NORTH_SB_IN_B1(Tile_X02_Y00_io2f_1),
		.SB_T0_NORTH_SB_IN_B17(Tile_X02_Y00_io2f_17),
		.SB_T0_NORTH_SB_IN_B17_ready(Tile_X02_Y01_SB_T0_NORTH_SB_IN_B17_ready),
		.SB_T0_NORTH_SB_IN_B17_valid(Tile_X02_Y00_io2f_17_valid),
		.SB_T0_NORTH_SB_IN_B1_ready(Tile_X02_Y01_SB_T0_NORTH_SB_IN_B1_ready),
		.SB_T0_NORTH_SB_IN_B1_valid(Tile_X02_Y00_io2f_1_valid),
		.SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_OUT_B17(Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_OUT_B17_ready(Tile_X02_Y00_f2io_17_ready),
		.SB_T0_NORTH_SB_OUT_B17_valid(Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B17_valid),
		.SB_T0_NORTH_SB_OUT_B1_ready(Tile_X02_Y00_f2io_1_ready),
		.SB_T0_NORTH_SB_OUT_B1_valid(Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B1_valid),
		.SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_IN_B17(Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_IN_B17_ready(Tile_X02_Y01_SB_T0_SOUTH_SB_IN_B17_ready),
		.SB_T0_SOUTH_SB_IN_B17_valid(Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B17_valid),
		.SB_T0_SOUTH_SB_IN_B1_ready(Tile_X02_Y01_SB_T0_SOUTH_SB_IN_B1_ready),
		.SB_T0_SOUTH_SB_IN_B1_valid(Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B1_valid),
		.SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_OUT_B17(Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_OUT_B17_ready(Tile_X02_Y02_SB_T0_NORTH_SB_IN_B17_ready),
		.SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B17_valid),
		.SB_T0_SOUTH_SB_OUT_B1_ready(Tile_X02_Y02_SB_T0_NORTH_SB_IN_B1_ready),
		.SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B1_valid),
		.SB_T0_WEST_SB_IN_B1(Tile_X01_Y01_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_WEST_SB_IN_B17(Tile_X01_Y01_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_WEST_SB_IN_B17_ready(Tile_X02_Y01_SB_T0_WEST_SB_IN_B17_ready),
		.SB_T0_WEST_SB_IN_B17_valid(Tile_X01_Y01_SB_T0_EAST_SB_OUT_B17_valid),
		.SB_T0_WEST_SB_IN_B1_ready(Tile_X02_Y01_SB_T0_WEST_SB_IN_B1_ready),
		.SB_T0_WEST_SB_IN_B1_valid(Tile_X01_Y01_SB_T0_EAST_SB_OUT_B1_valid),
		.SB_T0_WEST_SB_OUT_B1(Tile_X02_Y01_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_WEST_SB_OUT_B17(Tile_X02_Y01_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_WEST_SB_OUT_B17_ready(Tile_X01_Y01_SB_T0_EAST_SB_IN_B17_ready),
		.SB_T0_WEST_SB_OUT_B17_valid(Tile_X02_Y01_SB_T0_WEST_SB_OUT_B17_valid),
		.SB_T0_WEST_SB_OUT_B1_ready(Tile_X01_Y01_SB_T0_EAST_SB_IN_B1_ready),
		.SB_T0_WEST_SB_OUT_B1_valid(Tile_X02_Y01_SB_T0_WEST_SB_OUT_B1_valid),
		.SB_T1_EAST_SB_IN_B1(Tile_X03_Y01_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_EAST_SB_IN_B17(Tile_X03_Y01_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_EAST_SB_IN_B17_ready(Tile_X02_Y01_SB_T1_EAST_SB_IN_B17_ready),
		.SB_T1_EAST_SB_IN_B17_valid(Tile_X03_Y01_SB_T1_WEST_SB_OUT_B17_valid),
		.SB_T1_EAST_SB_IN_B1_ready(Tile_X02_Y01_SB_T1_EAST_SB_IN_B1_ready),
		.SB_T1_EAST_SB_IN_B1_valid(Tile_X03_Y01_SB_T1_WEST_SB_OUT_B1_valid),
		.SB_T1_EAST_SB_OUT_B1(Tile_X02_Y01_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_EAST_SB_OUT_B17(Tile_X02_Y01_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_EAST_SB_OUT_B17_ready(Tile_X03_Y01_SB_T1_WEST_SB_IN_B17_ready),
		.SB_T1_EAST_SB_OUT_B17_valid(Tile_X02_Y01_SB_T1_EAST_SB_OUT_B17_valid),
		.SB_T1_EAST_SB_OUT_B1_ready(Tile_X03_Y01_SB_T1_WEST_SB_IN_B1_ready),
		.SB_T1_EAST_SB_OUT_B1_valid(Tile_X02_Y01_SB_T1_EAST_SB_OUT_B1_valid),
		.SB_T1_NORTH_SB_IN_B1(Tile_X02_Y00_io2f_1),
		.SB_T1_NORTH_SB_IN_B17(Tile_X02_Y00_io2f_17),
		.SB_T1_NORTH_SB_IN_B17_ready(Tile_X02_Y01_SB_T1_NORTH_SB_IN_B17_ready),
		.SB_T1_NORTH_SB_IN_B17_valid(Tile_X02_Y00_io2f_17_valid),
		.SB_T1_NORTH_SB_IN_B1_ready(Tile_X02_Y01_SB_T1_NORTH_SB_IN_B1_ready),
		.SB_T1_NORTH_SB_IN_B1_valid(Tile_X02_Y00_io2f_1_valid),
		.SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y01_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_OUT_B17(Tile_X02_Y01_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T1_NORTH_SB_OUT_B17_valid(Tile_X02_Y01_SB_T1_NORTH_SB_OUT_B17_valid),
		.SB_T1_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T1_NORTH_SB_OUT_B1_valid(Tile_X02_Y01_SB_T1_NORTH_SB_OUT_B1_valid),
		.SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_IN_B17(Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_IN_B17_ready(Tile_X02_Y01_SB_T1_SOUTH_SB_IN_B17_ready),
		.SB_T1_SOUTH_SB_IN_B17_valid(Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B17_valid),
		.SB_T1_SOUTH_SB_IN_B1_ready(Tile_X02_Y01_SB_T1_SOUTH_SB_IN_B1_ready),
		.SB_T1_SOUTH_SB_IN_B1_valid(Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B1_valid),
		.SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_OUT_B17(Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_OUT_B17_ready(Tile_X02_Y02_SB_T1_NORTH_SB_IN_B17_ready),
		.SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B17_valid),
		.SB_T1_SOUTH_SB_OUT_B1_ready(Tile_X02_Y02_SB_T1_NORTH_SB_IN_B1_ready),
		.SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B1_valid),
		.SB_T1_WEST_SB_IN_B1(Tile_X01_Y01_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_WEST_SB_IN_B17(Tile_X01_Y01_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_WEST_SB_IN_B17_ready(Tile_X02_Y01_SB_T1_WEST_SB_IN_B17_ready),
		.SB_T1_WEST_SB_IN_B17_valid(Tile_X01_Y01_SB_T1_EAST_SB_OUT_B17_valid),
		.SB_T1_WEST_SB_IN_B1_ready(Tile_X02_Y01_SB_T1_WEST_SB_IN_B1_ready),
		.SB_T1_WEST_SB_IN_B1_valid(Tile_X01_Y01_SB_T1_EAST_SB_OUT_B1_valid),
		.SB_T1_WEST_SB_OUT_B1(Tile_X02_Y01_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_WEST_SB_OUT_B17(Tile_X02_Y01_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_WEST_SB_OUT_B17_ready(Tile_X01_Y01_SB_T1_EAST_SB_IN_B17_ready),
		.SB_T1_WEST_SB_OUT_B17_valid(Tile_X02_Y01_SB_T1_WEST_SB_OUT_B17_valid),
		.SB_T1_WEST_SB_OUT_B1_ready(Tile_X01_Y01_SB_T1_EAST_SB_IN_B1_ready),
		.SB_T1_WEST_SB_OUT_B1_valid(Tile_X02_Y01_SB_T1_WEST_SB_OUT_B1_valid),
		.SB_T2_EAST_SB_IN_B1(Tile_X03_Y01_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_EAST_SB_IN_B17(Tile_X03_Y01_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_EAST_SB_IN_B17_ready(Tile_X02_Y01_SB_T2_EAST_SB_IN_B17_ready),
		.SB_T2_EAST_SB_IN_B17_valid(Tile_X03_Y01_SB_T2_WEST_SB_OUT_B17_valid),
		.SB_T2_EAST_SB_IN_B1_ready(Tile_X02_Y01_SB_T2_EAST_SB_IN_B1_ready),
		.SB_T2_EAST_SB_IN_B1_valid(Tile_X03_Y01_SB_T2_WEST_SB_OUT_B1_valid),
		.SB_T2_EAST_SB_OUT_B1(Tile_X02_Y01_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_EAST_SB_OUT_B17(Tile_X02_Y01_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_EAST_SB_OUT_B17_ready(Tile_X03_Y01_SB_T2_WEST_SB_IN_B17_ready),
		.SB_T2_EAST_SB_OUT_B17_valid(Tile_X02_Y01_SB_T2_EAST_SB_OUT_B17_valid),
		.SB_T2_EAST_SB_OUT_B1_ready(Tile_X03_Y01_SB_T2_WEST_SB_IN_B1_ready),
		.SB_T2_EAST_SB_OUT_B1_valid(Tile_X02_Y01_SB_T2_EAST_SB_OUT_B1_valid),
		.SB_T2_NORTH_SB_IN_B1(Tile_X02_Y00_io2f_1),
		.SB_T2_NORTH_SB_IN_B17(Tile_X02_Y00_io2f_17),
		.SB_T2_NORTH_SB_IN_B17_ready(Tile_X02_Y01_SB_T2_NORTH_SB_IN_B17_ready),
		.SB_T2_NORTH_SB_IN_B17_valid(Tile_X02_Y00_io2f_17_valid),
		.SB_T2_NORTH_SB_IN_B1_ready(Tile_X02_Y01_SB_T2_NORTH_SB_IN_B1_ready),
		.SB_T2_NORTH_SB_IN_B1_valid(Tile_X02_Y00_io2f_1_valid),
		.SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y01_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_OUT_B17(Tile_X02_Y01_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T2_NORTH_SB_OUT_B17_valid(Tile_X02_Y01_SB_T2_NORTH_SB_OUT_B17_valid),
		.SB_T2_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T2_NORTH_SB_OUT_B1_valid(Tile_X02_Y01_SB_T2_NORTH_SB_OUT_B1_valid),
		.SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_IN_B17(Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_IN_B17_ready(Tile_X02_Y01_SB_T2_SOUTH_SB_IN_B17_ready),
		.SB_T2_SOUTH_SB_IN_B17_valid(Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B17_valid),
		.SB_T2_SOUTH_SB_IN_B1_ready(Tile_X02_Y01_SB_T2_SOUTH_SB_IN_B1_ready),
		.SB_T2_SOUTH_SB_IN_B1_valid(Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B1_valid),
		.SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_OUT_B17(Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_OUT_B17_ready(Tile_X02_Y02_SB_T2_NORTH_SB_IN_B17_ready),
		.SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B17_valid),
		.SB_T2_SOUTH_SB_OUT_B1_ready(Tile_X02_Y02_SB_T2_NORTH_SB_IN_B1_ready),
		.SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B1_valid),
		.SB_T2_WEST_SB_IN_B1(Tile_X01_Y01_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_WEST_SB_IN_B17(Tile_X01_Y01_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_WEST_SB_IN_B17_ready(Tile_X02_Y01_SB_T2_WEST_SB_IN_B17_ready),
		.SB_T2_WEST_SB_IN_B17_valid(Tile_X01_Y01_SB_T2_EAST_SB_OUT_B17_valid),
		.SB_T2_WEST_SB_IN_B1_ready(Tile_X02_Y01_SB_T2_WEST_SB_IN_B1_ready),
		.SB_T2_WEST_SB_IN_B1_valid(Tile_X01_Y01_SB_T2_EAST_SB_OUT_B1_valid),
		.SB_T2_WEST_SB_OUT_B1(Tile_X02_Y01_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_WEST_SB_OUT_B17(Tile_X02_Y01_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_WEST_SB_OUT_B17_ready(Tile_X01_Y01_SB_T2_EAST_SB_IN_B17_ready),
		.SB_T2_WEST_SB_OUT_B17_valid(Tile_X02_Y01_SB_T2_WEST_SB_OUT_B17_valid),
		.SB_T2_WEST_SB_OUT_B1_ready(Tile_X01_Y01_SB_T2_EAST_SB_IN_B1_ready),
		.SB_T2_WEST_SB_OUT_B1_valid(Tile_X02_Y01_SB_T2_WEST_SB_OUT_B1_valid),
		.SB_T3_EAST_SB_IN_B1(Tile_X03_Y01_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_EAST_SB_IN_B17(Tile_X03_Y01_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_EAST_SB_IN_B17_ready(Tile_X02_Y01_SB_T3_EAST_SB_IN_B17_ready),
		.SB_T3_EAST_SB_IN_B17_valid(Tile_X03_Y01_SB_T3_WEST_SB_OUT_B17_valid),
		.SB_T3_EAST_SB_IN_B1_ready(Tile_X02_Y01_SB_T3_EAST_SB_IN_B1_ready),
		.SB_T3_EAST_SB_IN_B1_valid(Tile_X03_Y01_SB_T3_WEST_SB_OUT_B1_valid),
		.SB_T3_EAST_SB_OUT_B1(Tile_X02_Y01_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_EAST_SB_OUT_B17(Tile_X02_Y01_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_EAST_SB_OUT_B17_ready(Tile_X03_Y01_SB_T3_WEST_SB_IN_B17_ready),
		.SB_T3_EAST_SB_OUT_B17_valid(Tile_X02_Y01_SB_T3_EAST_SB_OUT_B17_valid),
		.SB_T3_EAST_SB_OUT_B1_ready(Tile_X03_Y01_SB_T3_WEST_SB_IN_B1_ready),
		.SB_T3_EAST_SB_OUT_B1_valid(Tile_X02_Y01_SB_T3_EAST_SB_OUT_B1_valid),
		.SB_T3_NORTH_SB_IN_B1(Tile_X02_Y00_io2f_1),
		.SB_T3_NORTH_SB_IN_B17(Tile_X02_Y00_io2f_17),
		.SB_T3_NORTH_SB_IN_B17_ready(Tile_X02_Y01_SB_T3_NORTH_SB_IN_B17_ready),
		.SB_T3_NORTH_SB_IN_B17_valid(Tile_X02_Y00_io2f_17_valid),
		.SB_T3_NORTH_SB_IN_B1_ready(Tile_X02_Y01_SB_T3_NORTH_SB_IN_B1_ready),
		.SB_T3_NORTH_SB_IN_B1_valid(Tile_X02_Y00_io2f_1_valid),
		.SB_T3_NORTH_SB_OUT_B1(Tile_X02_Y01_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_OUT_B17(Tile_X02_Y01_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T3_NORTH_SB_OUT_B17_valid(Tile_X02_Y01_SB_T3_NORTH_SB_OUT_B17_valid),
		.SB_T3_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T3_NORTH_SB_OUT_B1_valid(Tile_X02_Y01_SB_T3_NORTH_SB_OUT_B1_valid),
		.SB_T3_SOUTH_SB_IN_B1(Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_IN_B17(Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_IN_B17_ready(Tile_X02_Y01_SB_T3_SOUTH_SB_IN_B17_ready),
		.SB_T3_SOUTH_SB_IN_B17_valid(Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B17_valid),
		.SB_T3_SOUTH_SB_IN_B1_ready(Tile_X02_Y01_SB_T3_SOUTH_SB_IN_B1_ready),
		.SB_T3_SOUTH_SB_IN_B1_valid(Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B1_valid),
		.SB_T3_SOUTH_SB_OUT_B1(Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_OUT_B17(Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_OUT_B17_ready(Tile_X02_Y02_SB_T3_NORTH_SB_IN_B17_ready),
		.SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B17_valid),
		.SB_T3_SOUTH_SB_OUT_B1_ready(Tile_X02_Y02_SB_T3_NORTH_SB_IN_B1_ready),
		.SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B1_valid),
		.SB_T3_WEST_SB_IN_B1(Tile_X01_Y01_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_WEST_SB_IN_B17(Tile_X01_Y01_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_WEST_SB_IN_B17_ready(Tile_X02_Y01_SB_T3_WEST_SB_IN_B17_ready),
		.SB_T3_WEST_SB_IN_B17_valid(Tile_X01_Y01_SB_T3_EAST_SB_OUT_B17_valid),
		.SB_T3_WEST_SB_IN_B1_ready(Tile_X02_Y01_SB_T3_WEST_SB_IN_B1_ready),
		.SB_T3_WEST_SB_IN_B1_valid(Tile_X01_Y01_SB_T3_EAST_SB_OUT_B1_valid),
		.SB_T3_WEST_SB_OUT_B1(Tile_X02_Y01_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_WEST_SB_OUT_B17(Tile_X02_Y01_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_WEST_SB_OUT_B17_ready(Tile_X01_Y01_SB_T3_EAST_SB_IN_B17_ready),
		.SB_T3_WEST_SB_OUT_B17_valid(Tile_X02_Y01_SB_T3_WEST_SB_OUT_B17_valid),
		.SB_T3_WEST_SB_OUT_B1_ready(Tile_X01_Y01_SB_T3_EAST_SB_IN_B1_ready),
		.SB_T3_WEST_SB_OUT_B1_valid(Tile_X02_Y01_SB_T3_WEST_SB_OUT_B1_valid),
		.SB_T4_EAST_SB_IN_B1(Tile_X03_Y01_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_EAST_SB_IN_B17(Tile_X03_Y01_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_EAST_SB_IN_B17_ready(Tile_X02_Y01_SB_T4_EAST_SB_IN_B17_ready),
		.SB_T4_EAST_SB_IN_B17_valid(Tile_X03_Y01_SB_T4_WEST_SB_OUT_B17_valid),
		.SB_T4_EAST_SB_IN_B1_ready(Tile_X02_Y01_SB_T4_EAST_SB_IN_B1_ready),
		.SB_T4_EAST_SB_IN_B1_valid(Tile_X03_Y01_SB_T4_WEST_SB_OUT_B1_valid),
		.SB_T4_EAST_SB_OUT_B1(Tile_X02_Y01_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_EAST_SB_OUT_B17(Tile_X02_Y01_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_EAST_SB_OUT_B17_ready(Tile_X03_Y01_SB_T4_WEST_SB_IN_B17_ready),
		.SB_T4_EAST_SB_OUT_B17_valid(Tile_X02_Y01_SB_T4_EAST_SB_OUT_B17_valid),
		.SB_T4_EAST_SB_OUT_B1_ready(Tile_X03_Y01_SB_T4_WEST_SB_IN_B1_ready),
		.SB_T4_EAST_SB_OUT_B1_valid(Tile_X02_Y01_SB_T4_EAST_SB_OUT_B1_valid),
		.SB_T4_NORTH_SB_IN_B1(Tile_X02_Y00_io2f_1),
		.SB_T4_NORTH_SB_IN_B17(Tile_X02_Y00_io2f_17),
		.SB_T4_NORTH_SB_IN_B17_ready(Tile_X02_Y01_SB_T4_NORTH_SB_IN_B17_ready),
		.SB_T4_NORTH_SB_IN_B17_valid(Tile_X02_Y00_io2f_17_valid),
		.SB_T4_NORTH_SB_IN_B1_ready(Tile_X02_Y01_SB_T4_NORTH_SB_IN_B1_ready),
		.SB_T4_NORTH_SB_IN_B1_valid(Tile_X02_Y00_io2f_1_valid),
		.SB_T4_NORTH_SB_OUT_B1(Tile_X02_Y01_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_OUT_B17(Tile_X02_Y01_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T4_NORTH_SB_OUT_B17_valid(Tile_X02_Y01_SB_T4_NORTH_SB_OUT_B17_valid),
		.SB_T4_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T4_NORTH_SB_OUT_B1_valid(Tile_X02_Y01_SB_T4_NORTH_SB_OUT_B1_valid),
		.SB_T4_SOUTH_SB_IN_B1(Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_IN_B17(Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_IN_B17_ready(Tile_X02_Y01_SB_T4_SOUTH_SB_IN_B17_ready),
		.SB_T4_SOUTH_SB_IN_B17_valid(Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B17_valid),
		.SB_T4_SOUTH_SB_IN_B1_ready(Tile_X02_Y01_SB_T4_SOUTH_SB_IN_B1_ready),
		.SB_T4_SOUTH_SB_IN_B1_valid(Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B1_valid),
		.SB_T4_SOUTH_SB_OUT_B1(Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_OUT_B17(Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_OUT_B17_ready(Tile_X02_Y02_SB_T4_NORTH_SB_IN_B17_ready),
		.SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B17_valid),
		.SB_T4_SOUTH_SB_OUT_B1_ready(Tile_X02_Y02_SB_T4_NORTH_SB_IN_B1_ready),
		.SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B1_valid),
		.SB_T4_WEST_SB_IN_B1(Tile_X01_Y01_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_WEST_SB_IN_B17(Tile_X01_Y01_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_WEST_SB_IN_B17_ready(Tile_X02_Y01_SB_T4_WEST_SB_IN_B17_ready),
		.SB_T4_WEST_SB_IN_B17_valid(Tile_X01_Y01_SB_T4_EAST_SB_OUT_B17_valid),
		.SB_T4_WEST_SB_IN_B1_ready(Tile_X02_Y01_SB_T4_WEST_SB_IN_B1_ready),
		.SB_T4_WEST_SB_IN_B1_valid(Tile_X01_Y01_SB_T4_EAST_SB_OUT_B1_valid),
		.SB_T4_WEST_SB_OUT_B1(Tile_X02_Y01_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_WEST_SB_OUT_B17(Tile_X02_Y01_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_WEST_SB_OUT_B17_ready(Tile_X01_Y01_SB_T4_EAST_SB_IN_B17_ready),
		.SB_T4_WEST_SB_OUT_B17_valid(Tile_X02_Y01_SB_T4_WEST_SB_OUT_B17_valid),
		.SB_T4_WEST_SB_OUT_B1_ready(Tile_X01_Y01_SB_T4_EAST_SB_IN_B1_ready),
		.SB_T4_WEST_SB_OUT_B1_valid(Tile_X02_Y01_SB_T4_WEST_SB_OUT_B1_valid),
		.clk(Tile_X02_Y00_clk_out),
		.clk_out(Tile_X02_Y01_clk_out),
		.clk_pass_through(coreir_wrapInClock_inst2_out),
		.clk_pass_through_out_bot(Tile_X02_Y01_clk_pass_through_out_bot),
		.clk_pass_through_out_right(Tile_X02_Y01_clk_pass_through_out_right),
		.config_config_addr(Tile_X02_Y00_config_out_config_addr),
		.config_config_data(Tile_X02_Y00_config_out_config_data),
		.config_out_config_addr(Tile_X02_Y01_config_out_config_addr),
		.config_out_config_data(Tile_X02_Y01_config_out_config_data),
		.config_out_read(Tile_X02_Y01_config_out_read),
		.config_out_write(Tile_X02_Y01_config_out_write),
		.config_read(Tile_X02_Y00_config_out_read),
		.config_write(Tile_X02_Y00_config_out_write),
		.flush(Tile_X02_Y00_flush_out),
		.flush_out(Tile_X02_Y01_flush_out),
		.hi(Tile_X02_Y01_hi),
		.lo(Tile_X02_Y01_lo),
		.read_config_data(Tile_X02_Y01_read_config_data),
		.read_config_data_in(Tile_X02_Y00_read_config_data),
		.reset(Tile_X02_Y00_reset_out),
		.reset_out(Tile_X02_Y01_reset_out),
		.stall(Tile_X02_Y00_stall_out),
		.stall_out(Tile_X02_Y01_stall_out),
		.tile_id(Tile_X02_Y01_tile_id)
	);
	wire [15:0] Tile_X02_Y02_tile_id;
	assign Tile_X02_Y02_tile_id = {Tile_X02_Y02_lo[7], Tile_X02_Y02_lo[7], Tile_X02_Y02_lo[6], Tile_X02_Y02_lo[6], Tile_X02_Y02_lo[5], Tile_X02_Y02_lo[5], Tile_X02_Y02_hi[5], Tile_X02_Y02_lo[4], Tile_X02_Y02_lo[3], Tile_X02_Y02_lo[3], Tile_X02_Y02_lo[2], Tile_X02_Y02_lo[2], Tile_X02_Y02_lo[1], Tile_X02_Y02_lo[1], Tile_X02_Y02_hi[1], Tile_X02_Y02_lo[0]};
	Tile_PE Tile_X02_Y02(
		.SB_T0_EAST_SB_IN_B1(Tile_X03_Y02_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_EAST_SB_IN_B17(Tile_X03_Y02_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_EAST_SB_IN_B17_ready(Tile_X02_Y02_SB_T0_EAST_SB_IN_B17_ready),
		.SB_T0_EAST_SB_IN_B17_valid(Tile_X03_Y02_SB_T0_WEST_SB_OUT_B17_valid),
		.SB_T0_EAST_SB_IN_B1_ready(Tile_X02_Y02_SB_T0_EAST_SB_IN_B1_ready),
		.SB_T0_EAST_SB_IN_B1_valid(Tile_X03_Y02_SB_T0_WEST_SB_OUT_B1_valid),
		.SB_T0_EAST_SB_OUT_B1(Tile_X02_Y02_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_EAST_SB_OUT_B17(Tile_X02_Y02_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_EAST_SB_OUT_B17_ready(Tile_X03_Y02_SB_T0_WEST_SB_IN_B17_ready),
		.SB_T0_EAST_SB_OUT_B17_valid(Tile_X02_Y02_SB_T0_EAST_SB_OUT_B17_valid),
		.SB_T0_EAST_SB_OUT_B1_ready(Tile_X03_Y02_SB_T0_WEST_SB_IN_B1_ready),
		.SB_T0_EAST_SB_OUT_B1_valid(Tile_X02_Y02_SB_T0_EAST_SB_OUT_B1_valid),
		.SB_T0_NORTH_SB_IN_B1(Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_IN_B17(Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_IN_B17_ready(Tile_X02_Y02_SB_T0_NORTH_SB_IN_B17_ready),
		.SB_T0_NORTH_SB_IN_B17_valid(Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B17_valid),
		.SB_T0_NORTH_SB_IN_B1_ready(Tile_X02_Y02_SB_T0_NORTH_SB_IN_B1_ready),
		.SB_T0_NORTH_SB_IN_B1_valid(Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B1_valid),
		.SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_OUT_B17(Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_OUT_B17_ready(Tile_X02_Y01_SB_T0_SOUTH_SB_IN_B17_ready),
		.SB_T0_NORTH_SB_OUT_B17_valid(Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B17_valid),
		.SB_T0_NORTH_SB_OUT_B1_ready(Tile_X02_Y01_SB_T0_SOUTH_SB_IN_B1_ready),
		.SB_T0_NORTH_SB_OUT_B1_valid(Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B1_valid),
		.SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_IN_B17(Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_IN_B17_ready(Tile_X02_Y02_SB_T0_SOUTH_SB_IN_B17_ready),
		.SB_T0_SOUTH_SB_IN_B17_valid(Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B17_valid),
		.SB_T0_SOUTH_SB_IN_B1_ready(Tile_X02_Y02_SB_T0_SOUTH_SB_IN_B1_ready),
		.SB_T0_SOUTH_SB_IN_B1_valid(Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B1_valid),
		.SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_OUT_B17(Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_OUT_B17_ready(Tile_X02_Y03_SB_T0_NORTH_SB_IN_B17_ready),
		.SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B17_valid),
		.SB_T0_SOUTH_SB_OUT_B1_ready(Tile_X02_Y03_SB_T0_NORTH_SB_IN_B1_ready),
		.SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B1_valid),
		.SB_T0_WEST_SB_IN_B1(Tile_X01_Y02_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_WEST_SB_IN_B17(Tile_X01_Y02_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_WEST_SB_IN_B17_ready(Tile_X02_Y02_SB_T0_WEST_SB_IN_B17_ready),
		.SB_T0_WEST_SB_IN_B17_valid(Tile_X01_Y02_SB_T0_EAST_SB_OUT_B17_valid),
		.SB_T0_WEST_SB_IN_B1_ready(Tile_X02_Y02_SB_T0_WEST_SB_IN_B1_ready),
		.SB_T0_WEST_SB_IN_B1_valid(Tile_X01_Y02_SB_T0_EAST_SB_OUT_B1_valid),
		.SB_T0_WEST_SB_OUT_B1(Tile_X02_Y02_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_WEST_SB_OUT_B17(Tile_X02_Y02_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_WEST_SB_OUT_B17_ready(Tile_X01_Y02_SB_T0_EAST_SB_IN_B17_ready),
		.SB_T0_WEST_SB_OUT_B17_valid(Tile_X02_Y02_SB_T0_WEST_SB_OUT_B17_valid),
		.SB_T0_WEST_SB_OUT_B1_ready(Tile_X01_Y02_SB_T0_EAST_SB_IN_B1_ready),
		.SB_T0_WEST_SB_OUT_B1_valid(Tile_X02_Y02_SB_T0_WEST_SB_OUT_B1_valid),
		.SB_T1_EAST_SB_IN_B1(Tile_X03_Y02_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_EAST_SB_IN_B17(Tile_X03_Y02_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_EAST_SB_IN_B17_ready(Tile_X02_Y02_SB_T1_EAST_SB_IN_B17_ready),
		.SB_T1_EAST_SB_IN_B17_valid(Tile_X03_Y02_SB_T1_WEST_SB_OUT_B17_valid),
		.SB_T1_EAST_SB_IN_B1_ready(Tile_X02_Y02_SB_T1_EAST_SB_IN_B1_ready),
		.SB_T1_EAST_SB_IN_B1_valid(Tile_X03_Y02_SB_T1_WEST_SB_OUT_B1_valid),
		.SB_T1_EAST_SB_OUT_B1(Tile_X02_Y02_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_EAST_SB_OUT_B17(Tile_X02_Y02_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_EAST_SB_OUT_B17_ready(Tile_X03_Y02_SB_T1_WEST_SB_IN_B17_ready),
		.SB_T1_EAST_SB_OUT_B17_valid(Tile_X02_Y02_SB_T1_EAST_SB_OUT_B17_valid),
		.SB_T1_EAST_SB_OUT_B1_ready(Tile_X03_Y02_SB_T1_WEST_SB_IN_B1_ready),
		.SB_T1_EAST_SB_OUT_B1_valid(Tile_X02_Y02_SB_T1_EAST_SB_OUT_B1_valid),
		.SB_T1_NORTH_SB_IN_B1(Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_IN_B17(Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_IN_B17_ready(Tile_X02_Y02_SB_T1_NORTH_SB_IN_B17_ready),
		.SB_T1_NORTH_SB_IN_B17_valid(Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B17_valid),
		.SB_T1_NORTH_SB_IN_B1_ready(Tile_X02_Y02_SB_T1_NORTH_SB_IN_B1_ready),
		.SB_T1_NORTH_SB_IN_B1_valid(Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B1_valid),
		.SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_OUT_B17(Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_OUT_B17_ready(Tile_X02_Y01_SB_T1_SOUTH_SB_IN_B17_ready),
		.SB_T1_NORTH_SB_OUT_B17_valid(Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B17_valid),
		.SB_T1_NORTH_SB_OUT_B1_ready(Tile_X02_Y01_SB_T1_SOUTH_SB_IN_B1_ready),
		.SB_T1_NORTH_SB_OUT_B1_valid(Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B1_valid),
		.SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_IN_B17(Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_IN_B17_ready(Tile_X02_Y02_SB_T1_SOUTH_SB_IN_B17_ready),
		.SB_T1_SOUTH_SB_IN_B17_valid(Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B17_valid),
		.SB_T1_SOUTH_SB_IN_B1_ready(Tile_X02_Y02_SB_T1_SOUTH_SB_IN_B1_ready),
		.SB_T1_SOUTH_SB_IN_B1_valid(Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B1_valid),
		.SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_OUT_B17(Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_OUT_B17_ready(Tile_X02_Y03_SB_T1_NORTH_SB_IN_B17_ready),
		.SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B17_valid),
		.SB_T1_SOUTH_SB_OUT_B1_ready(Tile_X02_Y03_SB_T1_NORTH_SB_IN_B1_ready),
		.SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B1_valid),
		.SB_T1_WEST_SB_IN_B1(Tile_X01_Y02_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_WEST_SB_IN_B17(Tile_X01_Y02_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_WEST_SB_IN_B17_ready(Tile_X02_Y02_SB_T1_WEST_SB_IN_B17_ready),
		.SB_T1_WEST_SB_IN_B17_valid(Tile_X01_Y02_SB_T1_EAST_SB_OUT_B17_valid),
		.SB_T1_WEST_SB_IN_B1_ready(Tile_X02_Y02_SB_T1_WEST_SB_IN_B1_ready),
		.SB_T1_WEST_SB_IN_B1_valid(Tile_X01_Y02_SB_T1_EAST_SB_OUT_B1_valid),
		.SB_T1_WEST_SB_OUT_B1(Tile_X02_Y02_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_WEST_SB_OUT_B17(Tile_X02_Y02_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_WEST_SB_OUT_B17_ready(Tile_X01_Y02_SB_T1_EAST_SB_IN_B17_ready),
		.SB_T1_WEST_SB_OUT_B17_valid(Tile_X02_Y02_SB_T1_WEST_SB_OUT_B17_valid),
		.SB_T1_WEST_SB_OUT_B1_ready(Tile_X01_Y02_SB_T1_EAST_SB_IN_B1_ready),
		.SB_T1_WEST_SB_OUT_B1_valid(Tile_X02_Y02_SB_T1_WEST_SB_OUT_B1_valid),
		.SB_T2_EAST_SB_IN_B1(Tile_X03_Y02_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_EAST_SB_IN_B17(Tile_X03_Y02_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_EAST_SB_IN_B17_ready(Tile_X02_Y02_SB_T2_EAST_SB_IN_B17_ready),
		.SB_T2_EAST_SB_IN_B17_valid(Tile_X03_Y02_SB_T2_WEST_SB_OUT_B17_valid),
		.SB_T2_EAST_SB_IN_B1_ready(Tile_X02_Y02_SB_T2_EAST_SB_IN_B1_ready),
		.SB_T2_EAST_SB_IN_B1_valid(Tile_X03_Y02_SB_T2_WEST_SB_OUT_B1_valid),
		.SB_T2_EAST_SB_OUT_B1(Tile_X02_Y02_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_EAST_SB_OUT_B17(Tile_X02_Y02_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_EAST_SB_OUT_B17_ready(Tile_X03_Y02_SB_T2_WEST_SB_IN_B17_ready),
		.SB_T2_EAST_SB_OUT_B17_valid(Tile_X02_Y02_SB_T2_EAST_SB_OUT_B17_valid),
		.SB_T2_EAST_SB_OUT_B1_ready(Tile_X03_Y02_SB_T2_WEST_SB_IN_B1_ready),
		.SB_T2_EAST_SB_OUT_B1_valid(Tile_X02_Y02_SB_T2_EAST_SB_OUT_B1_valid),
		.SB_T2_NORTH_SB_IN_B1(Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_IN_B17(Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_IN_B17_ready(Tile_X02_Y02_SB_T2_NORTH_SB_IN_B17_ready),
		.SB_T2_NORTH_SB_IN_B17_valid(Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B17_valid),
		.SB_T2_NORTH_SB_IN_B1_ready(Tile_X02_Y02_SB_T2_NORTH_SB_IN_B1_ready),
		.SB_T2_NORTH_SB_IN_B1_valid(Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B1_valid),
		.SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_OUT_B17(Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_OUT_B17_ready(Tile_X02_Y01_SB_T2_SOUTH_SB_IN_B17_ready),
		.SB_T2_NORTH_SB_OUT_B17_valid(Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B17_valid),
		.SB_T2_NORTH_SB_OUT_B1_ready(Tile_X02_Y01_SB_T2_SOUTH_SB_IN_B1_ready),
		.SB_T2_NORTH_SB_OUT_B1_valid(Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B1_valid),
		.SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_IN_B17(Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_IN_B17_ready(Tile_X02_Y02_SB_T2_SOUTH_SB_IN_B17_ready),
		.SB_T2_SOUTH_SB_IN_B17_valid(Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B17_valid),
		.SB_T2_SOUTH_SB_IN_B1_ready(Tile_X02_Y02_SB_T2_SOUTH_SB_IN_B1_ready),
		.SB_T2_SOUTH_SB_IN_B1_valid(Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B1_valid),
		.SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_OUT_B17(Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_OUT_B17_ready(Tile_X02_Y03_SB_T2_NORTH_SB_IN_B17_ready),
		.SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B17_valid),
		.SB_T2_SOUTH_SB_OUT_B1_ready(Tile_X02_Y03_SB_T2_NORTH_SB_IN_B1_ready),
		.SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B1_valid),
		.SB_T2_WEST_SB_IN_B1(Tile_X01_Y02_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_WEST_SB_IN_B17(Tile_X01_Y02_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_WEST_SB_IN_B17_ready(Tile_X02_Y02_SB_T2_WEST_SB_IN_B17_ready),
		.SB_T2_WEST_SB_IN_B17_valid(Tile_X01_Y02_SB_T2_EAST_SB_OUT_B17_valid),
		.SB_T2_WEST_SB_IN_B1_ready(Tile_X02_Y02_SB_T2_WEST_SB_IN_B1_ready),
		.SB_T2_WEST_SB_IN_B1_valid(Tile_X01_Y02_SB_T2_EAST_SB_OUT_B1_valid),
		.SB_T2_WEST_SB_OUT_B1(Tile_X02_Y02_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_WEST_SB_OUT_B17(Tile_X02_Y02_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_WEST_SB_OUT_B17_ready(Tile_X01_Y02_SB_T2_EAST_SB_IN_B17_ready),
		.SB_T2_WEST_SB_OUT_B17_valid(Tile_X02_Y02_SB_T2_WEST_SB_OUT_B17_valid),
		.SB_T2_WEST_SB_OUT_B1_ready(Tile_X01_Y02_SB_T2_EAST_SB_IN_B1_ready),
		.SB_T2_WEST_SB_OUT_B1_valid(Tile_X02_Y02_SB_T2_WEST_SB_OUT_B1_valid),
		.SB_T3_EAST_SB_IN_B1(Tile_X03_Y02_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_EAST_SB_IN_B17(Tile_X03_Y02_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_EAST_SB_IN_B17_ready(Tile_X02_Y02_SB_T3_EAST_SB_IN_B17_ready),
		.SB_T3_EAST_SB_IN_B17_valid(Tile_X03_Y02_SB_T3_WEST_SB_OUT_B17_valid),
		.SB_T3_EAST_SB_IN_B1_ready(Tile_X02_Y02_SB_T3_EAST_SB_IN_B1_ready),
		.SB_T3_EAST_SB_IN_B1_valid(Tile_X03_Y02_SB_T3_WEST_SB_OUT_B1_valid),
		.SB_T3_EAST_SB_OUT_B1(Tile_X02_Y02_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_EAST_SB_OUT_B17(Tile_X02_Y02_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_EAST_SB_OUT_B17_ready(Tile_X03_Y02_SB_T3_WEST_SB_IN_B17_ready),
		.SB_T3_EAST_SB_OUT_B17_valid(Tile_X02_Y02_SB_T3_EAST_SB_OUT_B17_valid),
		.SB_T3_EAST_SB_OUT_B1_ready(Tile_X03_Y02_SB_T3_WEST_SB_IN_B1_ready),
		.SB_T3_EAST_SB_OUT_B1_valid(Tile_X02_Y02_SB_T3_EAST_SB_OUT_B1_valid),
		.SB_T3_NORTH_SB_IN_B1(Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_IN_B17(Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_IN_B17_ready(Tile_X02_Y02_SB_T3_NORTH_SB_IN_B17_ready),
		.SB_T3_NORTH_SB_IN_B17_valid(Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B17_valid),
		.SB_T3_NORTH_SB_IN_B1_ready(Tile_X02_Y02_SB_T3_NORTH_SB_IN_B1_ready),
		.SB_T3_NORTH_SB_IN_B1_valid(Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B1_valid),
		.SB_T3_NORTH_SB_OUT_B1(Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_OUT_B17(Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_OUT_B17_ready(Tile_X02_Y01_SB_T3_SOUTH_SB_IN_B17_ready),
		.SB_T3_NORTH_SB_OUT_B17_valid(Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B17_valid),
		.SB_T3_NORTH_SB_OUT_B1_ready(Tile_X02_Y01_SB_T3_SOUTH_SB_IN_B1_ready),
		.SB_T3_NORTH_SB_OUT_B1_valid(Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B1_valid),
		.SB_T3_SOUTH_SB_IN_B1(Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_IN_B17(Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_IN_B17_ready(Tile_X02_Y02_SB_T3_SOUTH_SB_IN_B17_ready),
		.SB_T3_SOUTH_SB_IN_B17_valid(Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B17_valid),
		.SB_T3_SOUTH_SB_IN_B1_ready(Tile_X02_Y02_SB_T3_SOUTH_SB_IN_B1_ready),
		.SB_T3_SOUTH_SB_IN_B1_valid(Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B1_valid),
		.SB_T3_SOUTH_SB_OUT_B1(Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_OUT_B17(Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_OUT_B17_ready(Tile_X02_Y03_SB_T3_NORTH_SB_IN_B17_ready),
		.SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B17_valid),
		.SB_T3_SOUTH_SB_OUT_B1_ready(Tile_X02_Y03_SB_T3_NORTH_SB_IN_B1_ready),
		.SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B1_valid),
		.SB_T3_WEST_SB_IN_B1(Tile_X01_Y02_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_WEST_SB_IN_B17(Tile_X01_Y02_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_WEST_SB_IN_B17_ready(Tile_X02_Y02_SB_T3_WEST_SB_IN_B17_ready),
		.SB_T3_WEST_SB_IN_B17_valid(Tile_X01_Y02_SB_T3_EAST_SB_OUT_B17_valid),
		.SB_T3_WEST_SB_IN_B1_ready(Tile_X02_Y02_SB_T3_WEST_SB_IN_B1_ready),
		.SB_T3_WEST_SB_IN_B1_valid(Tile_X01_Y02_SB_T3_EAST_SB_OUT_B1_valid),
		.SB_T3_WEST_SB_OUT_B1(Tile_X02_Y02_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_WEST_SB_OUT_B17(Tile_X02_Y02_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_WEST_SB_OUT_B17_ready(Tile_X01_Y02_SB_T3_EAST_SB_IN_B17_ready),
		.SB_T3_WEST_SB_OUT_B17_valid(Tile_X02_Y02_SB_T3_WEST_SB_OUT_B17_valid),
		.SB_T3_WEST_SB_OUT_B1_ready(Tile_X01_Y02_SB_T3_EAST_SB_IN_B1_ready),
		.SB_T3_WEST_SB_OUT_B1_valid(Tile_X02_Y02_SB_T3_WEST_SB_OUT_B1_valid),
		.SB_T4_EAST_SB_IN_B1(Tile_X03_Y02_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_EAST_SB_IN_B17(Tile_X03_Y02_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_EAST_SB_IN_B17_ready(Tile_X02_Y02_SB_T4_EAST_SB_IN_B17_ready),
		.SB_T4_EAST_SB_IN_B17_valid(Tile_X03_Y02_SB_T4_WEST_SB_OUT_B17_valid),
		.SB_T4_EAST_SB_IN_B1_ready(Tile_X02_Y02_SB_T4_EAST_SB_IN_B1_ready),
		.SB_T4_EAST_SB_IN_B1_valid(Tile_X03_Y02_SB_T4_WEST_SB_OUT_B1_valid),
		.SB_T4_EAST_SB_OUT_B1(Tile_X02_Y02_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_EAST_SB_OUT_B17(Tile_X02_Y02_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_EAST_SB_OUT_B17_ready(Tile_X03_Y02_SB_T4_WEST_SB_IN_B17_ready),
		.SB_T4_EAST_SB_OUT_B17_valid(Tile_X02_Y02_SB_T4_EAST_SB_OUT_B17_valid),
		.SB_T4_EAST_SB_OUT_B1_ready(Tile_X03_Y02_SB_T4_WEST_SB_IN_B1_ready),
		.SB_T4_EAST_SB_OUT_B1_valid(Tile_X02_Y02_SB_T4_EAST_SB_OUT_B1_valid),
		.SB_T4_NORTH_SB_IN_B1(Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_IN_B17(Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_IN_B17_ready(Tile_X02_Y02_SB_T4_NORTH_SB_IN_B17_ready),
		.SB_T4_NORTH_SB_IN_B17_valid(Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B17_valid),
		.SB_T4_NORTH_SB_IN_B1_ready(Tile_X02_Y02_SB_T4_NORTH_SB_IN_B1_ready),
		.SB_T4_NORTH_SB_IN_B1_valid(Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B1_valid),
		.SB_T4_NORTH_SB_OUT_B1(Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_OUT_B17(Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_OUT_B17_ready(Tile_X02_Y01_SB_T4_SOUTH_SB_IN_B17_ready),
		.SB_T4_NORTH_SB_OUT_B17_valid(Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B17_valid),
		.SB_T4_NORTH_SB_OUT_B1_ready(Tile_X02_Y01_SB_T4_SOUTH_SB_IN_B1_ready),
		.SB_T4_NORTH_SB_OUT_B1_valid(Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B1_valid),
		.SB_T4_SOUTH_SB_IN_B1(Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_IN_B17(Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_IN_B17_ready(Tile_X02_Y02_SB_T4_SOUTH_SB_IN_B17_ready),
		.SB_T4_SOUTH_SB_IN_B17_valid(Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B17_valid),
		.SB_T4_SOUTH_SB_IN_B1_ready(Tile_X02_Y02_SB_T4_SOUTH_SB_IN_B1_ready),
		.SB_T4_SOUTH_SB_IN_B1_valid(Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B1_valid),
		.SB_T4_SOUTH_SB_OUT_B1(Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_OUT_B17(Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_OUT_B17_ready(Tile_X02_Y03_SB_T4_NORTH_SB_IN_B17_ready),
		.SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B17_valid),
		.SB_T4_SOUTH_SB_OUT_B1_ready(Tile_X02_Y03_SB_T4_NORTH_SB_IN_B1_ready),
		.SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B1_valid),
		.SB_T4_WEST_SB_IN_B1(Tile_X01_Y02_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_WEST_SB_IN_B17(Tile_X01_Y02_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_WEST_SB_IN_B17_ready(Tile_X02_Y02_SB_T4_WEST_SB_IN_B17_ready),
		.SB_T4_WEST_SB_IN_B17_valid(Tile_X01_Y02_SB_T4_EAST_SB_OUT_B17_valid),
		.SB_T4_WEST_SB_IN_B1_ready(Tile_X02_Y02_SB_T4_WEST_SB_IN_B1_ready),
		.SB_T4_WEST_SB_IN_B1_valid(Tile_X01_Y02_SB_T4_EAST_SB_OUT_B1_valid),
		.SB_T4_WEST_SB_OUT_B1(Tile_X02_Y02_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_WEST_SB_OUT_B17(Tile_X02_Y02_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_WEST_SB_OUT_B17_ready(Tile_X01_Y02_SB_T4_EAST_SB_IN_B17_ready),
		.SB_T4_WEST_SB_OUT_B17_valid(Tile_X02_Y02_SB_T4_WEST_SB_OUT_B17_valid),
		.SB_T4_WEST_SB_OUT_B1_ready(Tile_X01_Y02_SB_T4_EAST_SB_IN_B1_ready),
		.SB_T4_WEST_SB_OUT_B1_valid(Tile_X02_Y02_SB_T4_WEST_SB_OUT_B1_valid),
		.clk(Tile_X02_Y01_clk_out),
		.clk_out(Tile_X02_Y02_clk_out),
		.clk_pass_through(Tile_X02_Y01_clk_pass_through_out_bot),
		.clk_pass_through_out_bot(Tile_X02_Y02_clk_pass_through_out_bot),
		.clk_pass_through_out_right(Tile_X02_Y02_clk_pass_through_out_right),
		.config_config_addr(Tile_X02_Y01_config_out_config_addr),
		.config_config_data(Tile_X02_Y01_config_out_config_data),
		.config_out_config_addr(Tile_X02_Y02_config_out_config_addr),
		.config_out_config_data(Tile_X02_Y02_config_out_config_data),
		.config_out_read(Tile_X02_Y02_config_out_read),
		.config_out_write(Tile_X02_Y02_config_out_write),
		.config_read(Tile_X02_Y01_config_out_read),
		.config_write(Tile_X02_Y01_config_out_write),
		.flush(Tile_X02_Y01_flush_out),
		.flush_out(Tile_X02_Y02_flush_out),
		.hi(Tile_X02_Y02_hi),
		.lo(Tile_X02_Y02_lo),
		.read_config_data(Tile_X02_Y02_read_config_data),
		.read_config_data_in(Tile_X02_Y01_read_config_data),
		.reset(Tile_X02_Y01_reset_out),
		.reset_out(Tile_X02_Y02_reset_out),
		.stall(Tile_X02_Y01_stall_out),
		.stall_out(Tile_X02_Y02_stall_out),
		.tile_id(Tile_X02_Y02_tile_id)
	);
	wire [15:0] Tile_X02_Y03_tile_id;
	assign Tile_X02_Y03_tile_id = {Tile_X02_Y03_lo[7], Tile_X02_Y03_lo[7], Tile_X02_Y03_lo[6], Tile_X02_Y03_lo[6], Tile_X02_Y03_lo[5], Tile_X02_Y03_lo[5], Tile_X02_Y03_hi[5], Tile_X02_Y03_lo[4], Tile_X02_Y03_lo[3], Tile_X02_Y03_lo[3], Tile_X02_Y03_lo[2], Tile_X02_Y03_lo[2], Tile_X02_Y03_lo[1], Tile_X02_Y03_lo[1], Tile_X02_Y03_hi[1], Tile_X02_Y03_hi[0]};
	Tile_PE Tile_X02_Y03(
		.SB_T0_EAST_SB_IN_B1(Tile_X03_Y03_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_EAST_SB_IN_B17(Tile_X03_Y03_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_EAST_SB_IN_B17_ready(Tile_X02_Y03_SB_T0_EAST_SB_IN_B17_ready),
		.SB_T0_EAST_SB_IN_B17_valid(Tile_X03_Y03_SB_T0_WEST_SB_OUT_B17_valid),
		.SB_T0_EAST_SB_IN_B1_ready(Tile_X02_Y03_SB_T0_EAST_SB_IN_B1_ready),
		.SB_T0_EAST_SB_IN_B1_valid(Tile_X03_Y03_SB_T0_WEST_SB_OUT_B1_valid),
		.SB_T0_EAST_SB_OUT_B1(Tile_X02_Y03_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_EAST_SB_OUT_B17(Tile_X02_Y03_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_EAST_SB_OUT_B17_ready(Tile_X03_Y03_SB_T0_WEST_SB_IN_B17_ready),
		.SB_T0_EAST_SB_OUT_B17_valid(Tile_X02_Y03_SB_T0_EAST_SB_OUT_B17_valid),
		.SB_T0_EAST_SB_OUT_B1_ready(Tile_X03_Y03_SB_T0_WEST_SB_IN_B1_ready),
		.SB_T0_EAST_SB_OUT_B1_valid(Tile_X02_Y03_SB_T0_EAST_SB_OUT_B1_valid),
		.SB_T0_NORTH_SB_IN_B1(Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_IN_B17(Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_IN_B17_ready(Tile_X02_Y03_SB_T0_NORTH_SB_IN_B17_ready),
		.SB_T0_NORTH_SB_IN_B17_valid(Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B17_valid),
		.SB_T0_NORTH_SB_IN_B1_ready(Tile_X02_Y03_SB_T0_NORTH_SB_IN_B1_ready),
		.SB_T0_NORTH_SB_IN_B1_valid(Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B1_valid),
		.SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_OUT_B17(Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_OUT_B17_ready(Tile_X02_Y02_SB_T0_SOUTH_SB_IN_B17_ready),
		.SB_T0_NORTH_SB_OUT_B17_valid(Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B17_valid),
		.SB_T0_NORTH_SB_OUT_B1_ready(Tile_X02_Y02_SB_T0_SOUTH_SB_IN_B1_ready),
		.SB_T0_NORTH_SB_OUT_B1_valid(Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B1_valid),
		.SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_IN_B17(Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_IN_B17_ready(Tile_X02_Y03_SB_T0_SOUTH_SB_IN_B17_ready),
		.SB_T0_SOUTH_SB_IN_B17_valid(Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B17_valid),
		.SB_T0_SOUTH_SB_IN_B1_ready(Tile_X02_Y03_SB_T0_SOUTH_SB_IN_B1_ready),
		.SB_T0_SOUTH_SB_IN_B1_valid(Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B1_valid),
		.SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_OUT_B17(Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_OUT_B17_ready(Tile_X02_Y04_SB_T0_NORTH_SB_IN_B17_ready),
		.SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B17_valid),
		.SB_T0_SOUTH_SB_OUT_B1_ready(Tile_X02_Y04_SB_T0_NORTH_SB_IN_B1_ready),
		.SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B1_valid),
		.SB_T0_WEST_SB_IN_B1(Tile_X01_Y03_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_WEST_SB_IN_B17(Tile_X01_Y03_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_WEST_SB_IN_B17_ready(Tile_X02_Y03_SB_T0_WEST_SB_IN_B17_ready),
		.SB_T0_WEST_SB_IN_B17_valid(Tile_X01_Y03_SB_T0_EAST_SB_OUT_B17_valid),
		.SB_T0_WEST_SB_IN_B1_ready(Tile_X02_Y03_SB_T0_WEST_SB_IN_B1_ready),
		.SB_T0_WEST_SB_IN_B1_valid(Tile_X01_Y03_SB_T0_EAST_SB_OUT_B1_valid),
		.SB_T0_WEST_SB_OUT_B1(Tile_X02_Y03_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_WEST_SB_OUT_B17(Tile_X02_Y03_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_WEST_SB_OUT_B17_ready(Tile_X01_Y03_SB_T0_EAST_SB_IN_B17_ready),
		.SB_T0_WEST_SB_OUT_B17_valid(Tile_X02_Y03_SB_T0_WEST_SB_OUT_B17_valid),
		.SB_T0_WEST_SB_OUT_B1_ready(Tile_X01_Y03_SB_T0_EAST_SB_IN_B1_ready),
		.SB_T0_WEST_SB_OUT_B1_valid(Tile_X02_Y03_SB_T0_WEST_SB_OUT_B1_valid),
		.SB_T1_EAST_SB_IN_B1(Tile_X03_Y03_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_EAST_SB_IN_B17(Tile_X03_Y03_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_EAST_SB_IN_B17_ready(Tile_X02_Y03_SB_T1_EAST_SB_IN_B17_ready),
		.SB_T1_EAST_SB_IN_B17_valid(Tile_X03_Y03_SB_T1_WEST_SB_OUT_B17_valid),
		.SB_T1_EAST_SB_IN_B1_ready(Tile_X02_Y03_SB_T1_EAST_SB_IN_B1_ready),
		.SB_T1_EAST_SB_IN_B1_valid(Tile_X03_Y03_SB_T1_WEST_SB_OUT_B1_valid),
		.SB_T1_EAST_SB_OUT_B1(Tile_X02_Y03_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_EAST_SB_OUT_B17(Tile_X02_Y03_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_EAST_SB_OUT_B17_ready(Tile_X03_Y03_SB_T1_WEST_SB_IN_B17_ready),
		.SB_T1_EAST_SB_OUT_B17_valid(Tile_X02_Y03_SB_T1_EAST_SB_OUT_B17_valid),
		.SB_T1_EAST_SB_OUT_B1_ready(Tile_X03_Y03_SB_T1_WEST_SB_IN_B1_ready),
		.SB_T1_EAST_SB_OUT_B1_valid(Tile_X02_Y03_SB_T1_EAST_SB_OUT_B1_valid),
		.SB_T1_NORTH_SB_IN_B1(Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_IN_B17(Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_IN_B17_ready(Tile_X02_Y03_SB_T1_NORTH_SB_IN_B17_ready),
		.SB_T1_NORTH_SB_IN_B17_valid(Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B17_valid),
		.SB_T1_NORTH_SB_IN_B1_ready(Tile_X02_Y03_SB_T1_NORTH_SB_IN_B1_ready),
		.SB_T1_NORTH_SB_IN_B1_valid(Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B1_valid),
		.SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_OUT_B17(Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_OUT_B17_ready(Tile_X02_Y02_SB_T1_SOUTH_SB_IN_B17_ready),
		.SB_T1_NORTH_SB_OUT_B17_valid(Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B17_valid),
		.SB_T1_NORTH_SB_OUT_B1_ready(Tile_X02_Y02_SB_T1_SOUTH_SB_IN_B1_ready),
		.SB_T1_NORTH_SB_OUT_B1_valid(Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B1_valid),
		.SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_IN_B17(Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_IN_B17_ready(Tile_X02_Y03_SB_T1_SOUTH_SB_IN_B17_ready),
		.SB_T1_SOUTH_SB_IN_B17_valid(Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B17_valid),
		.SB_T1_SOUTH_SB_IN_B1_ready(Tile_X02_Y03_SB_T1_SOUTH_SB_IN_B1_ready),
		.SB_T1_SOUTH_SB_IN_B1_valid(Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B1_valid),
		.SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_OUT_B17(Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_OUT_B17_ready(Tile_X02_Y04_SB_T1_NORTH_SB_IN_B17_ready),
		.SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B17_valid),
		.SB_T1_SOUTH_SB_OUT_B1_ready(Tile_X02_Y04_SB_T1_NORTH_SB_IN_B1_ready),
		.SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B1_valid),
		.SB_T1_WEST_SB_IN_B1(Tile_X01_Y03_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_WEST_SB_IN_B17(Tile_X01_Y03_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_WEST_SB_IN_B17_ready(Tile_X02_Y03_SB_T1_WEST_SB_IN_B17_ready),
		.SB_T1_WEST_SB_IN_B17_valid(Tile_X01_Y03_SB_T1_EAST_SB_OUT_B17_valid),
		.SB_T1_WEST_SB_IN_B1_ready(Tile_X02_Y03_SB_T1_WEST_SB_IN_B1_ready),
		.SB_T1_WEST_SB_IN_B1_valid(Tile_X01_Y03_SB_T1_EAST_SB_OUT_B1_valid),
		.SB_T1_WEST_SB_OUT_B1(Tile_X02_Y03_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_WEST_SB_OUT_B17(Tile_X02_Y03_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_WEST_SB_OUT_B17_ready(Tile_X01_Y03_SB_T1_EAST_SB_IN_B17_ready),
		.SB_T1_WEST_SB_OUT_B17_valid(Tile_X02_Y03_SB_T1_WEST_SB_OUT_B17_valid),
		.SB_T1_WEST_SB_OUT_B1_ready(Tile_X01_Y03_SB_T1_EAST_SB_IN_B1_ready),
		.SB_T1_WEST_SB_OUT_B1_valid(Tile_X02_Y03_SB_T1_WEST_SB_OUT_B1_valid),
		.SB_T2_EAST_SB_IN_B1(Tile_X03_Y03_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_EAST_SB_IN_B17(Tile_X03_Y03_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_EAST_SB_IN_B17_ready(Tile_X02_Y03_SB_T2_EAST_SB_IN_B17_ready),
		.SB_T2_EAST_SB_IN_B17_valid(Tile_X03_Y03_SB_T2_WEST_SB_OUT_B17_valid),
		.SB_T2_EAST_SB_IN_B1_ready(Tile_X02_Y03_SB_T2_EAST_SB_IN_B1_ready),
		.SB_T2_EAST_SB_IN_B1_valid(Tile_X03_Y03_SB_T2_WEST_SB_OUT_B1_valid),
		.SB_T2_EAST_SB_OUT_B1(Tile_X02_Y03_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_EAST_SB_OUT_B17(Tile_X02_Y03_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_EAST_SB_OUT_B17_ready(Tile_X03_Y03_SB_T2_WEST_SB_IN_B17_ready),
		.SB_T2_EAST_SB_OUT_B17_valid(Tile_X02_Y03_SB_T2_EAST_SB_OUT_B17_valid),
		.SB_T2_EAST_SB_OUT_B1_ready(Tile_X03_Y03_SB_T2_WEST_SB_IN_B1_ready),
		.SB_T2_EAST_SB_OUT_B1_valid(Tile_X02_Y03_SB_T2_EAST_SB_OUT_B1_valid),
		.SB_T2_NORTH_SB_IN_B1(Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_IN_B17(Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_IN_B17_ready(Tile_X02_Y03_SB_T2_NORTH_SB_IN_B17_ready),
		.SB_T2_NORTH_SB_IN_B17_valid(Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B17_valid),
		.SB_T2_NORTH_SB_IN_B1_ready(Tile_X02_Y03_SB_T2_NORTH_SB_IN_B1_ready),
		.SB_T2_NORTH_SB_IN_B1_valid(Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B1_valid),
		.SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_OUT_B17(Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_OUT_B17_ready(Tile_X02_Y02_SB_T2_SOUTH_SB_IN_B17_ready),
		.SB_T2_NORTH_SB_OUT_B17_valid(Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B17_valid),
		.SB_T2_NORTH_SB_OUT_B1_ready(Tile_X02_Y02_SB_T2_SOUTH_SB_IN_B1_ready),
		.SB_T2_NORTH_SB_OUT_B1_valid(Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B1_valid),
		.SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_IN_B17(Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_IN_B17_ready(Tile_X02_Y03_SB_T2_SOUTH_SB_IN_B17_ready),
		.SB_T2_SOUTH_SB_IN_B17_valid(Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B17_valid),
		.SB_T2_SOUTH_SB_IN_B1_ready(Tile_X02_Y03_SB_T2_SOUTH_SB_IN_B1_ready),
		.SB_T2_SOUTH_SB_IN_B1_valid(Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B1_valid),
		.SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_OUT_B17(Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_OUT_B17_ready(Tile_X02_Y04_SB_T2_NORTH_SB_IN_B17_ready),
		.SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B17_valid),
		.SB_T2_SOUTH_SB_OUT_B1_ready(Tile_X02_Y04_SB_T2_NORTH_SB_IN_B1_ready),
		.SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B1_valid),
		.SB_T2_WEST_SB_IN_B1(Tile_X01_Y03_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_WEST_SB_IN_B17(Tile_X01_Y03_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_WEST_SB_IN_B17_ready(Tile_X02_Y03_SB_T2_WEST_SB_IN_B17_ready),
		.SB_T2_WEST_SB_IN_B17_valid(Tile_X01_Y03_SB_T2_EAST_SB_OUT_B17_valid),
		.SB_T2_WEST_SB_IN_B1_ready(Tile_X02_Y03_SB_T2_WEST_SB_IN_B1_ready),
		.SB_T2_WEST_SB_IN_B1_valid(Tile_X01_Y03_SB_T2_EAST_SB_OUT_B1_valid),
		.SB_T2_WEST_SB_OUT_B1(Tile_X02_Y03_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_WEST_SB_OUT_B17(Tile_X02_Y03_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_WEST_SB_OUT_B17_ready(Tile_X01_Y03_SB_T2_EAST_SB_IN_B17_ready),
		.SB_T2_WEST_SB_OUT_B17_valid(Tile_X02_Y03_SB_T2_WEST_SB_OUT_B17_valid),
		.SB_T2_WEST_SB_OUT_B1_ready(Tile_X01_Y03_SB_T2_EAST_SB_IN_B1_ready),
		.SB_T2_WEST_SB_OUT_B1_valid(Tile_X02_Y03_SB_T2_WEST_SB_OUT_B1_valid),
		.SB_T3_EAST_SB_IN_B1(Tile_X03_Y03_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_EAST_SB_IN_B17(Tile_X03_Y03_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_EAST_SB_IN_B17_ready(Tile_X02_Y03_SB_T3_EAST_SB_IN_B17_ready),
		.SB_T3_EAST_SB_IN_B17_valid(Tile_X03_Y03_SB_T3_WEST_SB_OUT_B17_valid),
		.SB_T3_EAST_SB_IN_B1_ready(Tile_X02_Y03_SB_T3_EAST_SB_IN_B1_ready),
		.SB_T3_EAST_SB_IN_B1_valid(Tile_X03_Y03_SB_T3_WEST_SB_OUT_B1_valid),
		.SB_T3_EAST_SB_OUT_B1(Tile_X02_Y03_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_EAST_SB_OUT_B17(Tile_X02_Y03_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_EAST_SB_OUT_B17_ready(Tile_X03_Y03_SB_T3_WEST_SB_IN_B17_ready),
		.SB_T3_EAST_SB_OUT_B17_valid(Tile_X02_Y03_SB_T3_EAST_SB_OUT_B17_valid),
		.SB_T3_EAST_SB_OUT_B1_ready(Tile_X03_Y03_SB_T3_WEST_SB_IN_B1_ready),
		.SB_T3_EAST_SB_OUT_B1_valid(Tile_X02_Y03_SB_T3_EAST_SB_OUT_B1_valid),
		.SB_T3_NORTH_SB_IN_B1(Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_IN_B17(Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_IN_B17_ready(Tile_X02_Y03_SB_T3_NORTH_SB_IN_B17_ready),
		.SB_T3_NORTH_SB_IN_B17_valid(Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B17_valid),
		.SB_T3_NORTH_SB_IN_B1_ready(Tile_X02_Y03_SB_T3_NORTH_SB_IN_B1_ready),
		.SB_T3_NORTH_SB_IN_B1_valid(Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B1_valid),
		.SB_T3_NORTH_SB_OUT_B1(Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_OUT_B17(Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_OUT_B17_ready(Tile_X02_Y02_SB_T3_SOUTH_SB_IN_B17_ready),
		.SB_T3_NORTH_SB_OUT_B17_valid(Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B17_valid),
		.SB_T3_NORTH_SB_OUT_B1_ready(Tile_X02_Y02_SB_T3_SOUTH_SB_IN_B1_ready),
		.SB_T3_NORTH_SB_OUT_B1_valid(Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B1_valid),
		.SB_T3_SOUTH_SB_IN_B1(Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_IN_B17(Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_IN_B17_ready(Tile_X02_Y03_SB_T3_SOUTH_SB_IN_B17_ready),
		.SB_T3_SOUTH_SB_IN_B17_valid(Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B17_valid),
		.SB_T3_SOUTH_SB_IN_B1_ready(Tile_X02_Y03_SB_T3_SOUTH_SB_IN_B1_ready),
		.SB_T3_SOUTH_SB_IN_B1_valid(Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B1_valid),
		.SB_T3_SOUTH_SB_OUT_B1(Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_OUT_B17(Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_OUT_B17_ready(Tile_X02_Y04_SB_T3_NORTH_SB_IN_B17_ready),
		.SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B17_valid),
		.SB_T3_SOUTH_SB_OUT_B1_ready(Tile_X02_Y04_SB_T3_NORTH_SB_IN_B1_ready),
		.SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B1_valid),
		.SB_T3_WEST_SB_IN_B1(Tile_X01_Y03_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_WEST_SB_IN_B17(Tile_X01_Y03_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_WEST_SB_IN_B17_ready(Tile_X02_Y03_SB_T3_WEST_SB_IN_B17_ready),
		.SB_T3_WEST_SB_IN_B17_valid(Tile_X01_Y03_SB_T3_EAST_SB_OUT_B17_valid),
		.SB_T3_WEST_SB_IN_B1_ready(Tile_X02_Y03_SB_T3_WEST_SB_IN_B1_ready),
		.SB_T3_WEST_SB_IN_B1_valid(Tile_X01_Y03_SB_T3_EAST_SB_OUT_B1_valid),
		.SB_T3_WEST_SB_OUT_B1(Tile_X02_Y03_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_WEST_SB_OUT_B17(Tile_X02_Y03_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_WEST_SB_OUT_B17_ready(Tile_X01_Y03_SB_T3_EAST_SB_IN_B17_ready),
		.SB_T3_WEST_SB_OUT_B17_valid(Tile_X02_Y03_SB_T3_WEST_SB_OUT_B17_valid),
		.SB_T3_WEST_SB_OUT_B1_ready(Tile_X01_Y03_SB_T3_EAST_SB_IN_B1_ready),
		.SB_T3_WEST_SB_OUT_B1_valid(Tile_X02_Y03_SB_T3_WEST_SB_OUT_B1_valid),
		.SB_T4_EAST_SB_IN_B1(Tile_X03_Y03_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_EAST_SB_IN_B17(Tile_X03_Y03_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_EAST_SB_IN_B17_ready(Tile_X02_Y03_SB_T4_EAST_SB_IN_B17_ready),
		.SB_T4_EAST_SB_IN_B17_valid(Tile_X03_Y03_SB_T4_WEST_SB_OUT_B17_valid),
		.SB_T4_EAST_SB_IN_B1_ready(Tile_X02_Y03_SB_T4_EAST_SB_IN_B1_ready),
		.SB_T4_EAST_SB_IN_B1_valid(Tile_X03_Y03_SB_T4_WEST_SB_OUT_B1_valid),
		.SB_T4_EAST_SB_OUT_B1(Tile_X02_Y03_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_EAST_SB_OUT_B17(Tile_X02_Y03_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_EAST_SB_OUT_B17_ready(Tile_X03_Y03_SB_T4_WEST_SB_IN_B17_ready),
		.SB_T4_EAST_SB_OUT_B17_valid(Tile_X02_Y03_SB_T4_EAST_SB_OUT_B17_valid),
		.SB_T4_EAST_SB_OUT_B1_ready(Tile_X03_Y03_SB_T4_WEST_SB_IN_B1_ready),
		.SB_T4_EAST_SB_OUT_B1_valid(Tile_X02_Y03_SB_T4_EAST_SB_OUT_B1_valid),
		.SB_T4_NORTH_SB_IN_B1(Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_IN_B17(Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_IN_B17_ready(Tile_X02_Y03_SB_T4_NORTH_SB_IN_B17_ready),
		.SB_T4_NORTH_SB_IN_B17_valid(Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B17_valid),
		.SB_T4_NORTH_SB_IN_B1_ready(Tile_X02_Y03_SB_T4_NORTH_SB_IN_B1_ready),
		.SB_T4_NORTH_SB_IN_B1_valid(Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B1_valid),
		.SB_T4_NORTH_SB_OUT_B1(Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_OUT_B17(Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_OUT_B17_ready(Tile_X02_Y02_SB_T4_SOUTH_SB_IN_B17_ready),
		.SB_T4_NORTH_SB_OUT_B17_valid(Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B17_valid),
		.SB_T4_NORTH_SB_OUT_B1_ready(Tile_X02_Y02_SB_T4_SOUTH_SB_IN_B1_ready),
		.SB_T4_NORTH_SB_OUT_B1_valid(Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B1_valid),
		.SB_T4_SOUTH_SB_IN_B1(Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_IN_B17(Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_IN_B17_ready(Tile_X02_Y03_SB_T4_SOUTH_SB_IN_B17_ready),
		.SB_T4_SOUTH_SB_IN_B17_valid(Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B17_valid),
		.SB_T4_SOUTH_SB_IN_B1_ready(Tile_X02_Y03_SB_T4_SOUTH_SB_IN_B1_ready),
		.SB_T4_SOUTH_SB_IN_B1_valid(Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B1_valid),
		.SB_T4_SOUTH_SB_OUT_B1(Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_OUT_B17(Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_OUT_B17_ready(Tile_X02_Y04_SB_T4_NORTH_SB_IN_B17_ready),
		.SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B17_valid),
		.SB_T4_SOUTH_SB_OUT_B1_ready(Tile_X02_Y04_SB_T4_NORTH_SB_IN_B1_ready),
		.SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B1_valid),
		.SB_T4_WEST_SB_IN_B1(Tile_X01_Y03_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_WEST_SB_IN_B17(Tile_X01_Y03_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_WEST_SB_IN_B17_ready(Tile_X02_Y03_SB_T4_WEST_SB_IN_B17_ready),
		.SB_T4_WEST_SB_IN_B17_valid(Tile_X01_Y03_SB_T4_EAST_SB_OUT_B17_valid),
		.SB_T4_WEST_SB_IN_B1_ready(Tile_X02_Y03_SB_T4_WEST_SB_IN_B1_ready),
		.SB_T4_WEST_SB_IN_B1_valid(Tile_X01_Y03_SB_T4_EAST_SB_OUT_B1_valid),
		.SB_T4_WEST_SB_OUT_B1(Tile_X02_Y03_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_WEST_SB_OUT_B17(Tile_X02_Y03_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_WEST_SB_OUT_B17_ready(Tile_X01_Y03_SB_T4_EAST_SB_IN_B17_ready),
		.SB_T4_WEST_SB_OUT_B17_valid(Tile_X02_Y03_SB_T4_WEST_SB_OUT_B17_valid),
		.SB_T4_WEST_SB_OUT_B1_ready(Tile_X01_Y03_SB_T4_EAST_SB_IN_B1_ready),
		.SB_T4_WEST_SB_OUT_B1_valid(Tile_X02_Y03_SB_T4_WEST_SB_OUT_B1_valid),
		.clk(Tile_X02_Y02_clk_out),
		.clk_out(Tile_X02_Y03_clk_out),
		.clk_pass_through(Tile_X02_Y02_clk_pass_through_out_bot),
		.clk_pass_through_out_bot(Tile_X02_Y03_clk_pass_through_out_bot),
		.clk_pass_through_out_right(Tile_X02_Y03_clk_pass_through_out_right),
		.config_config_addr(Tile_X02_Y02_config_out_config_addr),
		.config_config_data(Tile_X02_Y02_config_out_config_data),
		.config_out_config_addr(Tile_X02_Y03_config_out_config_addr),
		.config_out_config_data(Tile_X02_Y03_config_out_config_data),
		.config_out_read(Tile_X02_Y03_config_out_read),
		.config_out_write(Tile_X02_Y03_config_out_write),
		.config_read(Tile_X02_Y02_config_out_read),
		.config_write(Tile_X02_Y02_config_out_write),
		.flush(Tile_X02_Y02_flush_out),
		.flush_out(Tile_X02_Y03_flush_out),
		.hi(Tile_X02_Y03_hi),
		.lo(Tile_X02_Y03_lo),
		.read_config_data(Tile_X02_Y03_read_config_data),
		.read_config_data_in(Tile_X02_Y02_read_config_data),
		.reset(Tile_X02_Y02_reset_out),
		.reset_out(Tile_X02_Y03_reset_out),
		.stall(Tile_X02_Y02_stall_out),
		.stall_out(Tile_X02_Y03_stall_out),
		.tile_id(Tile_X02_Y03_tile_id)
	);
	wire [15:0] Tile_X02_Y04_tile_id;
	assign Tile_X02_Y04_tile_id = {Tile_X02_Y04_lo[7], Tile_X02_Y04_lo[7], Tile_X02_Y04_lo[6], Tile_X02_Y04_lo[6], Tile_X02_Y04_lo[5], Tile_X02_Y04_lo[5], Tile_X02_Y04_hi[5], Tile_X02_Y04_lo[4], Tile_X02_Y04_lo[3], Tile_X02_Y04_lo[3], Tile_X02_Y04_lo[2], Tile_X02_Y04_lo[2], Tile_X02_Y04_lo[1], Tile_X02_Y04_hi[1], Tile_X02_Y04_lo[0], Tile_X02_Y04_lo[0]};
	Tile_PE Tile_X02_Y04(
		.SB_T0_EAST_SB_IN_B1(Tile_X03_Y04_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_EAST_SB_IN_B17(Tile_X03_Y04_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_EAST_SB_IN_B17_ready(Tile_X02_Y04_SB_T0_EAST_SB_IN_B17_ready),
		.SB_T0_EAST_SB_IN_B17_valid(Tile_X03_Y04_SB_T0_WEST_SB_OUT_B17_valid),
		.SB_T0_EAST_SB_IN_B1_ready(Tile_X02_Y04_SB_T0_EAST_SB_IN_B1_ready),
		.SB_T0_EAST_SB_IN_B1_valid(Tile_X03_Y04_SB_T0_WEST_SB_OUT_B1_valid),
		.SB_T0_EAST_SB_OUT_B1(Tile_X02_Y04_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_EAST_SB_OUT_B17(Tile_X02_Y04_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_EAST_SB_OUT_B17_ready(Tile_X03_Y04_SB_T0_WEST_SB_IN_B17_ready),
		.SB_T0_EAST_SB_OUT_B17_valid(Tile_X02_Y04_SB_T0_EAST_SB_OUT_B17_valid),
		.SB_T0_EAST_SB_OUT_B1_ready(Tile_X03_Y04_SB_T0_WEST_SB_IN_B1_ready),
		.SB_T0_EAST_SB_OUT_B1_valid(Tile_X02_Y04_SB_T0_EAST_SB_OUT_B1_valid),
		.SB_T0_NORTH_SB_IN_B1(Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_IN_B17(Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_IN_B17_ready(Tile_X02_Y04_SB_T0_NORTH_SB_IN_B17_ready),
		.SB_T0_NORTH_SB_IN_B17_valid(Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B17_valid),
		.SB_T0_NORTH_SB_IN_B1_ready(Tile_X02_Y04_SB_T0_NORTH_SB_IN_B1_ready),
		.SB_T0_NORTH_SB_IN_B1_valid(Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B1_valid),
		.SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_OUT_B17(Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_OUT_B17_ready(Tile_X02_Y03_SB_T0_SOUTH_SB_IN_B17_ready),
		.SB_T0_NORTH_SB_OUT_B17_valid(Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B17_valid),
		.SB_T0_NORTH_SB_OUT_B1_ready(Tile_X02_Y03_SB_T0_SOUTH_SB_IN_B1_ready),
		.SB_T0_NORTH_SB_OUT_B1_valid(Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B1_valid),
		.SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
		.SB_T0_SOUTH_SB_IN_B17(const_0_17_out),
		.SB_T0_SOUTH_SB_IN_B17_ready(Tile_X02_Y04_SB_T0_SOUTH_SB_IN_B17_ready),
		.SB_T0_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T0_SOUTH_SB_IN_B1_ready(Tile_X02_Y04_SB_T0_SOUTH_SB_IN_B1_ready),
		.SB_T0_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_OUT_B17(Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B17_valid),
		.SB_T0_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B1_valid),
		.SB_T0_WEST_SB_IN_B1(Tile_X01_Y04_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_WEST_SB_IN_B17(Tile_X01_Y04_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_WEST_SB_IN_B17_ready(Tile_X02_Y04_SB_T0_WEST_SB_IN_B17_ready),
		.SB_T0_WEST_SB_IN_B17_valid(Tile_X01_Y04_SB_T0_EAST_SB_OUT_B17_valid),
		.SB_T0_WEST_SB_IN_B1_ready(Tile_X02_Y04_SB_T0_WEST_SB_IN_B1_ready),
		.SB_T0_WEST_SB_IN_B1_valid(Tile_X01_Y04_SB_T0_EAST_SB_OUT_B1_valid),
		.SB_T0_WEST_SB_OUT_B1(Tile_X02_Y04_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_WEST_SB_OUT_B17(Tile_X02_Y04_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_WEST_SB_OUT_B17_ready(Tile_X01_Y04_SB_T0_EAST_SB_IN_B17_ready),
		.SB_T0_WEST_SB_OUT_B17_valid(Tile_X02_Y04_SB_T0_WEST_SB_OUT_B17_valid),
		.SB_T0_WEST_SB_OUT_B1_ready(Tile_X01_Y04_SB_T0_EAST_SB_IN_B1_ready),
		.SB_T0_WEST_SB_OUT_B1_valid(Tile_X02_Y04_SB_T0_WEST_SB_OUT_B1_valid),
		.SB_T1_EAST_SB_IN_B1(Tile_X03_Y04_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_EAST_SB_IN_B17(Tile_X03_Y04_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_EAST_SB_IN_B17_ready(Tile_X02_Y04_SB_T1_EAST_SB_IN_B17_ready),
		.SB_T1_EAST_SB_IN_B17_valid(Tile_X03_Y04_SB_T1_WEST_SB_OUT_B17_valid),
		.SB_T1_EAST_SB_IN_B1_ready(Tile_X02_Y04_SB_T1_EAST_SB_IN_B1_ready),
		.SB_T1_EAST_SB_IN_B1_valid(Tile_X03_Y04_SB_T1_WEST_SB_OUT_B1_valid),
		.SB_T1_EAST_SB_OUT_B1(Tile_X02_Y04_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_EAST_SB_OUT_B17(Tile_X02_Y04_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_EAST_SB_OUT_B17_ready(Tile_X03_Y04_SB_T1_WEST_SB_IN_B17_ready),
		.SB_T1_EAST_SB_OUT_B17_valid(Tile_X02_Y04_SB_T1_EAST_SB_OUT_B17_valid),
		.SB_T1_EAST_SB_OUT_B1_ready(Tile_X03_Y04_SB_T1_WEST_SB_IN_B1_ready),
		.SB_T1_EAST_SB_OUT_B1_valid(Tile_X02_Y04_SB_T1_EAST_SB_OUT_B1_valid),
		.SB_T1_NORTH_SB_IN_B1(Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_IN_B17(Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_IN_B17_ready(Tile_X02_Y04_SB_T1_NORTH_SB_IN_B17_ready),
		.SB_T1_NORTH_SB_IN_B17_valid(Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B17_valid),
		.SB_T1_NORTH_SB_IN_B1_ready(Tile_X02_Y04_SB_T1_NORTH_SB_IN_B1_ready),
		.SB_T1_NORTH_SB_IN_B1_valid(Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B1_valid),
		.SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_OUT_B17(Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_OUT_B17_ready(Tile_X02_Y03_SB_T1_SOUTH_SB_IN_B17_ready),
		.SB_T1_NORTH_SB_OUT_B17_valid(Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B17_valid),
		.SB_T1_NORTH_SB_OUT_B1_ready(Tile_X02_Y03_SB_T1_SOUTH_SB_IN_B1_ready),
		.SB_T1_NORTH_SB_OUT_B1_valid(Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B1_valid),
		.SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
		.SB_T1_SOUTH_SB_IN_B17(const_0_17_out),
		.SB_T1_SOUTH_SB_IN_B17_ready(Tile_X02_Y04_SB_T1_SOUTH_SB_IN_B17_ready),
		.SB_T1_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T1_SOUTH_SB_IN_B1_ready(Tile_X02_Y04_SB_T1_SOUTH_SB_IN_B1_ready),
		.SB_T1_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_OUT_B17(Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B17_valid),
		.SB_T1_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B1_valid),
		.SB_T1_WEST_SB_IN_B1(Tile_X01_Y04_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_WEST_SB_IN_B17(Tile_X01_Y04_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_WEST_SB_IN_B17_ready(Tile_X02_Y04_SB_T1_WEST_SB_IN_B17_ready),
		.SB_T1_WEST_SB_IN_B17_valid(Tile_X01_Y04_SB_T1_EAST_SB_OUT_B17_valid),
		.SB_T1_WEST_SB_IN_B1_ready(Tile_X02_Y04_SB_T1_WEST_SB_IN_B1_ready),
		.SB_T1_WEST_SB_IN_B1_valid(Tile_X01_Y04_SB_T1_EAST_SB_OUT_B1_valid),
		.SB_T1_WEST_SB_OUT_B1(Tile_X02_Y04_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_WEST_SB_OUT_B17(Tile_X02_Y04_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_WEST_SB_OUT_B17_ready(Tile_X01_Y04_SB_T1_EAST_SB_IN_B17_ready),
		.SB_T1_WEST_SB_OUT_B17_valid(Tile_X02_Y04_SB_T1_WEST_SB_OUT_B17_valid),
		.SB_T1_WEST_SB_OUT_B1_ready(Tile_X01_Y04_SB_T1_EAST_SB_IN_B1_ready),
		.SB_T1_WEST_SB_OUT_B1_valid(Tile_X02_Y04_SB_T1_WEST_SB_OUT_B1_valid),
		.SB_T2_EAST_SB_IN_B1(Tile_X03_Y04_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_EAST_SB_IN_B17(Tile_X03_Y04_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_EAST_SB_IN_B17_ready(Tile_X02_Y04_SB_T2_EAST_SB_IN_B17_ready),
		.SB_T2_EAST_SB_IN_B17_valid(Tile_X03_Y04_SB_T2_WEST_SB_OUT_B17_valid),
		.SB_T2_EAST_SB_IN_B1_ready(Tile_X02_Y04_SB_T2_EAST_SB_IN_B1_ready),
		.SB_T2_EAST_SB_IN_B1_valid(Tile_X03_Y04_SB_T2_WEST_SB_OUT_B1_valid),
		.SB_T2_EAST_SB_OUT_B1(Tile_X02_Y04_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_EAST_SB_OUT_B17(Tile_X02_Y04_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_EAST_SB_OUT_B17_ready(Tile_X03_Y04_SB_T2_WEST_SB_IN_B17_ready),
		.SB_T2_EAST_SB_OUT_B17_valid(Tile_X02_Y04_SB_T2_EAST_SB_OUT_B17_valid),
		.SB_T2_EAST_SB_OUT_B1_ready(Tile_X03_Y04_SB_T2_WEST_SB_IN_B1_ready),
		.SB_T2_EAST_SB_OUT_B1_valid(Tile_X02_Y04_SB_T2_EAST_SB_OUT_B1_valid),
		.SB_T2_NORTH_SB_IN_B1(Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_IN_B17(Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_IN_B17_ready(Tile_X02_Y04_SB_T2_NORTH_SB_IN_B17_ready),
		.SB_T2_NORTH_SB_IN_B17_valid(Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B17_valid),
		.SB_T2_NORTH_SB_IN_B1_ready(Tile_X02_Y04_SB_T2_NORTH_SB_IN_B1_ready),
		.SB_T2_NORTH_SB_IN_B1_valid(Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B1_valid),
		.SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_OUT_B17(Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_OUT_B17_ready(Tile_X02_Y03_SB_T2_SOUTH_SB_IN_B17_ready),
		.SB_T2_NORTH_SB_OUT_B17_valid(Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B17_valid),
		.SB_T2_NORTH_SB_OUT_B1_ready(Tile_X02_Y03_SB_T2_SOUTH_SB_IN_B1_ready),
		.SB_T2_NORTH_SB_OUT_B1_valid(Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B1_valid),
		.SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
		.SB_T2_SOUTH_SB_IN_B17(const_0_17_out),
		.SB_T2_SOUTH_SB_IN_B17_ready(Tile_X02_Y04_SB_T2_SOUTH_SB_IN_B17_ready),
		.SB_T2_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T2_SOUTH_SB_IN_B1_ready(Tile_X02_Y04_SB_T2_SOUTH_SB_IN_B1_ready),
		.SB_T2_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_OUT_B17(Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B17_valid),
		.SB_T2_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B1_valid),
		.SB_T2_WEST_SB_IN_B1(Tile_X01_Y04_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_WEST_SB_IN_B17(Tile_X01_Y04_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_WEST_SB_IN_B17_ready(Tile_X02_Y04_SB_T2_WEST_SB_IN_B17_ready),
		.SB_T2_WEST_SB_IN_B17_valid(Tile_X01_Y04_SB_T2_EAST_SB_OUT_B17_valid),
		.SB_T2_WEST_SB_IN_B1_ready(Tile_X02_Y04_SB_T2_WEST_SB_IN_B1_ready),
		.SB_T2_WEST_SB_IN_B1_valid(Tile_X01_Y04_SB_T2_EAST_SB_OUT_B1_valid),
		.SB_T2_WEST_SB_OUT_B1(Tile_X02_Y04_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_WEST_SB_OUT_B17(Tile_X02_Y04_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_WEST_SB_OUT_B17_ready(Tile_X01_Y04_SB_T2_EAST_SB_IN_B17_ready),
		.SB_T2_WEST_SB_OUT_B17_valid(Tile_X02_Y04_SB_T2_WEST_SB_OUT_B17_valid),
		.SB_T2_WEST_SB_OUT_B1_ready(Tile_X01_Y04_SB_T2_EAST_SB_IN_B1_ready),
		.SB_T2_WEST_SB_OUT_B1_valid(Tile_X02_Y04_SB_T2_WEST_SB_OUT_B1_valid),
		.SB_T3_EAST_SB_IN_B1(Tile_X03_Y04_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_EAST_SB_IN_B17(Tile_X03_Y04_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_EAST_SB_IN_B17_ready(Tile_X02_Y04_SB_T3_EAST_SB_IN_B17_ready),
		.SB_T3_EAST_SB_IN_B17_valid(Tile_X03_Y04_SB_T3_WEST_SB_OUT_B17_valid),
		.SB_T3_EAST_SB_IN_B1_ready(Tile_X02_Y04_SB_T3_EAST_SB_IN_B1_ready),
		.SB_T3_EAST_SB_IN_B1_valid(Tile_X03_Y04_SB_T3_WEST_SB_OUT_B1_valid),
		.SB_T3_EAST_SB_OUT_B1(Tile_X02_Y04_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_EAST_SB_OUT_B17(Tile_X02_Y04_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_EAST_SB_OUT_B17_ready(Tile_X03_Y04_SB_T3_WEST_SB_IN_B17_ready),
		.SB_T3_EAST_SB_OUT_B17_valid(Tile_X02_Y04_SB_T3_EAST_SB_OUT_B17_valid),
		.SB_T3_EAST_SB_OUT_B1_ready(Tile_X03_Y04_SB_T3_WEST_SB_IN_B1_ready),
		.SB_T3_EAST_SB_OUT_B1_valid(Tile_X02_Y04_SB_T3_EAST_SB_OUT_B1_valid),
		.SB_T3_NORTH_SB_IN_B1(Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_IN_B17(Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_IN_B17_ready(Tile_X02_Y04_SB_T3_NORTH_SB_IN_B17_ready),
		.SB_T3_NORTH_SB_IN_B17_valid(Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B17_valid),
		.SB_T3_NORTH_SB_IN_B1_ready(Tile_X02_Y04_SB_T3_NORTH_SB_IN_B1_ready),
		.SB_T3_NORTH_SB_IN_B1_valid(Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B1_valid),
		.SB_T3_NORTH_SB_OUT_B1(Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_OUT_B17(Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_OUT_B17_ready(Tile_X02_Y03_SB_T3_SOUTH_SB_IN_B17_ready),
		.SB_T3_NORTH_SB_OUT_B17_valid(Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B17_valid),
		.SB_T3_NORTH_SB_OUT_B1_ready(Tile_X02_Y03_SB_T3_SOUTH_SB_IN_B1_ready),
		.SB_T3_NORTH_SB_OUT_B1_valid(Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B1_valid),
		.SB_T3_SOUTH_SB_IN_B1(const_0_1_out),
		.SB_T3_SOUTH_SB_IN_B17(const_0_17_out),
		.SB_T3_SOUTH_SB_IN_B17_ready(Tile_X02_Y04_SB_T3_SOUTH_SB_IN_B17_ready),
		.SB_T3_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T3_SOUTH_SB_IN_B1_ready(Tile_X02_Y04_SB_T3_SOUTH_SB_IN_B1_ready),
		.SB_T3_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T3_SOUTH_SB_OUT_B1(Tile_X02_Y04_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_OUT_B17(Tile_X02_Y04_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X02_Y04_SB_T3_SOUTH_SB_OUT_B17_valid),
		.SB_T3_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X02_Y04_SB_T3_SOUTH_SB_OUT_B1_valid),
		.SB_T3_WEST_SB_IN_B1(Tile_X01_Y04_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_WEST_SB_IN_B17(Tile_X01_Y04_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_WEST_SB_IN_B17_ready(Tile_X02_Y04_SB_T3_WEST_SB_IN_B17_ready),
		.SB_T3_WEST_SB_IN_B17_valid(Tile_X01_Y04_SB_T3_EAST_SB_OUT_B17_valid),
		.SB_T3_WEST_SB_IN_B1_ready(Tile_X02_Y04_SB_T3_WEST_SB_IN_B1_ready),
		.SB_T3_WEST_SB_IN_B1_valid(Tile_X01_Y04_SB_T3_EAST_SB_OUT_B1_valid),
		.SB_T3_WEST_SB_OUT_B1(Tile_X02_Y04_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_WEST_SB_OUT_B17(Tile_X02_Y04_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_WEST_SB_OUT_B17_ready(Tile_X01_Y04_SB_T3_EAST_SB_IN_B17_ready),
		.SB_T3_WEST_SB_OUT_B17_valid(Tile_X02_Y04_SB_T3_WEST_SB_OUT_B17_valid),
		.SB_T3_WEST_SB_OUT_B1_ready(Tile_X01_Y04_SB_T3_EAST_SB_IN_B1_ready),
		.SB_T3_WEST_SB_OUT_B1_valid(Tile_X02_Y04_SB_T3_WEST_SB_OUT_B1_valid),
		.SB_T4_EAST_SB_IN_B1(Tile_X03_Y04_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_EAST_SB_IN_B17(Tile_X03_Y04_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_EAST_SB_IN_B17_ready(Tile_X02_Y04_SB_T4_EAST_SB_IN_B17_ready),
		.SB_T4_EAST_SB_IN_B17_valid(Tile_X03_Y04_SB_T4_WEST_SB_OUT_B17_valid),
		.SB_T4_EAST_SB_IN_B1_ready(Tile_X02_Y04_SB_T4_EAST_SB_IN_B1_ready),
		.SB_T4_EAST_SB_IN_B1_valid(Tile_X03_Y04_SB_T4_WEST_SB_OUT_B1_valid),
		.SB_T4_EAST_SB_OUT_B1(Tile_X02_Y04_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_EAST_SB_OUT_B17(Tile_X02_Y04_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_EAST_SB_OUT_B17_ready(Tile_X03_Y04_SB_T4_WEST_SB_IN_B17_ready),
		.SB_T4_EAST_SB_OUT_B17_valid(Tile_X02_Y04_SB_T4_EAST_SB_OUT_B17_valid),
		.SB_T4_EAST_SB_OUT_B1_ready(Tile_X03_Y04_SB_T4_WEST_SB_IN_B1_ready),
		.SB_T4_EAST_SB_OUT_B1_valid(Tile_X02_Y04_SB_T4_EAST_SB_OUT_B1_valid),
		.SB_T4_NORTH_SB_IN_B1(Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_IN_B17(Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_IN_B17_ready(Tile_X02_Y04_SB_T4_NORTH_SB_IN_B17_ready),
		.SB_T4_NORTH_SB_IN_B17_valid(Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B17_valid),
		.SB_T4_NORTH_SB_IN_B1_ready(Tile_X02_Y04_SB_T4_NORTH_SB_IN_B1_ready),
		.SB_T4_NORTH_SB_IN_B1_valid(Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B1_valid),
		.SB_T4_NORTH_SB_OUT_B1(Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_OUT_B17(Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_OUT_B17_ready(Tile_X02_Y03_SB_T4_SOUTH_SB_IN_B17_ready),
		.SB_T4_NORTH_SB_OUT_B17_valid(Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B17_valid),
		.SB_T4_NORTH_SB_OUT_B1_ready(Tile_X02_Y03_SB_T4_SOUTH_SB_IN_B1_ready),
		.SB_T4_NORTH_SB_OUT_B1_valid(Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B1_valid),
		.SB_T4_SOUTH_SB_IN_B1(const_0_1_out),
		.SB_T4_SOUTH_SB_IN_B17(const_0_17_out),
		.SB_T4_SOUTH_SB_IN_B17_ready(Tile_X02_Y04_SB_T4_SOUTH_SB_IN_B17_ready),
		.SB_T4_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T4_SOUTH_SB_IN_B1_ready(Tile_X02_Y04_SB_T4_SOUTH_SB_IN_B1_ready),
		.SB_T4_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T4_SOUTH_SB_OUT_B1(Tile_X02_Y04_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_OUT_B17(Tile_X02_Y04_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X02_Y04_SB_T4_SOUTH_SB_OUT_B17_valid),
		.SB_T4_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X02_Y04_SB_T4_SOUTH_SB_OUT_B1_valid),
		.SB_T4_WEST_SB_IN_B1(Tile_X01_Y04_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_WEST_SB_IN_B17(Tile_X01_Y04_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_WEST_SB_IN_B17_ready(Tile_X02_Y04_SB_T4_WEST_SB_IN_B17_ready),
		.SB_T4_WEST_SB_IN_B17_valid(Tile_X01_Y04_SB_T4_EAST_SB_OUT_B17_valid),
		.SB_T4_WEST_SB_IN_B1_ready(Tile_X02_Y04_SB_T4_WEST_SB_IN_B1_ready),
		.SB_T4_WEST_SB_IN_B1_valid(Tile_X01_Y04_SB_T4_EAST_SB_OUT_B1_valid),
		.SB_T4_WEST_SB_OUT_B1(Tile_X02_Y04_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_WEST_SB_OUT_B17(Tile_X02_Y04_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_WEST_SB_OUT_B17_ready(Tile_X01_Y04_SB_T4_EAST_SB_IN_B17_ready),
		.SB_T4_WEST_SB_OUT_B17_valid(Tile_X02_Y04_SB_T4_WEST_SB_OUT_B17_valid),
		.SB_T4_WEST_SB_OUT_B1_ready(Tile_X01_Y04_SB_T4_EAST_SB_IN_B1_ready),
		.SB_T4_WEST_SB_OUT_B1_valid(Tile_X02_Y04_SB_T4_WEST_SB_OUT_B1_valid),
		.clk(Tile_X02_Y03_clk_out),
		.clk_out(Tile_X02_Y04_clk_out),
		.clk_pass_through(Tile_X02_Y03_clk_pass_through_out_bot),
		.clk_pass_through_out_bot(Tile_X02_Y04_clk_pass_through_out_bot),
		.clk_pass_through_out_right(Tile_X02_Y04_clk_pass_through_out_right),
		.config_config_addr(Tile_X02_Y03_config_out_config_addr),
		.config_config_data(Tile_X02_Y03_config_out_config_data),
		.config_out_config_addr(Tile_X02_Y04_config_out_config_addr),
		.config_out_config_data(Tile_X02_Y04_config_out_config_data),
		.config_out_read(Tile_X02_Y04_config_out_read),
		.config_out_write(Tile_X02_Y04_config_out_write),
		.config_read(Tile_X02_Y03_config_out_read),
		.config_write(Tile_X02_Y03_config_out_write),
		.flush(Tile_X02_Y03_flush_out),
		.flush_out(Tile_X02_Y04_flush_out),
		.hi(Tile_X02_Y04_hi),
		.lo(Tile_X02_Y04_lo),
		.read_config_data(Tile_X02_Y04_read_config_data),
		.read_config_data_in(Tile_X02_Y03_read_config_data),
		.reset(Tile_X02_Y03_reset_out),
		.reset_out(Tile_X02_Y04_reset_out),
		.stall(Tile_X02_Y03_stall_out),
		.stall_out(Tile_X02_Y04_stall_out),
		.tile_id(Tile_X02_Y04_tile_id)
	);
	wire [31:0] Tile_X03_Y00_config_config_addr;
	assign Tile_X03_Y00_config_config_addr = {PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[31], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[30], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[29], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[28], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[27], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[26], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[25], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[24], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[23], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[22], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[21], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[20], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[19], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[18], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[17], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[16], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[15], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[14], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[13], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[12], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[11], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[10], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[9], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[8], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[7], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[6], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[5], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[4], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[3], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[2], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[1], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[0]};
	wire [31:0] Tile_X03_Y00_config_config_data;
	assign Tile_X03_Y00_config_config_data = {PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[63], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[62], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[61], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[60], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[59], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[58], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[57], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[56], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[55], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[54], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[53], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[52], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[51], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[50], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[49], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[48], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[47], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[46], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[45], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[44], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[43], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[42], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[41], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[40], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[39], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[38], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[37], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[36], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[35], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[34], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[33], PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[32]};
	wire [4:0] Tile_X03_Y00_io2f_17_ready;
	assign Tile_X03_Y00_io2f_17_ready = {Tile_X03_Y01_SB_T4_NORTH_SB_IN_B17_ready, Tile_X03_Y01_SB_T3_NORTH_SB_IN_B17_ready, Tile_X03_Y01_SB_T2_NORTH_SB_IN_B17_ready, Tile_X03_Y01_SB_T1_NORTH_SB_IN_B17_ready, Tile_X03_Y01_SB_T0_NORTH_SB_IN_B17_ready};
	wire [4:0] Tile_X03_Y00_io2f_1_ready;
	assign Tile_X03_Y00_io2f_1_ready = {Tile_X03_Y01_SB_T4_NORTH_SB_IN_B1_ready, Tile_X03_Y01_SB_T3_NORTH_SB_IN_B1_ready, Tile_X03_Y01_SB_T2_NORTH_SB_IN_B1_ready, Tile_X03_Y01_SB_T1_NORTH_SB_IN_B1_ready, Tile_X03_Y01_SB_T0_NORTH_SB_IN_B1_ready};
	wire [15:0] Tile_X03_Y00_tile_id;
	assign Tile_X03_Y00_tile_id = {Tile_X03_Y00_lo[7], Tile_X03_Y00_lo[7], Tile_X03_Y00_lo[6], Tile_X03_Y00_lo[6], Tile_X03_Y00_lo[5], Tile_X03_Y00_lo[5], Tile_X03_Y00_hi[5], Tile_X03_Y00_hi[4], Tile_X03_Y00_lo[3], Tile_X03_Y00_lo[3], Tile_X03_Y00_lo[2], Tile_X03_Y00_lo[2], Tile_X03_Y00_lo[1], Tile_X03_Y00_lo[1], Tile_X03_Y00_lo[0], Tile_X03_Y00_lo[0]};
	Tile_IOCoreReadyValid Tile_X03_Y00(
		.clk(clk),
		.clk_out(Tile_X03_Y00_clk_out),
		.config_config_addr(Tile_X03_Y00_config_config_addr),
		.config_config_data(Tile_X03_Y00_config_config_data),
		.config_out_config_addr(Tile_X03_Y00_config_out_config_addr),
		.config_out_config_data(Tile_X03_Y00_config_out_config_data),
		.config_out_read(Tile_X03_Y00_config_out_read),
		.config_out_write(Tile_X03_Y00_config_out_write),
		.config_read(PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[64]),
		.config_write(PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[65]),
		.f2io_1(Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B1),
		.f2io_17(Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B17),
		.f2io_17_ready(Tile_X03_Y00_f2io_17_ready),
		.f2io_17_valid(Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B17_valid),
		.f2io_1_ready(Tile_X03_Y00_f2io_1_ready),
		.f2io_1_valid(Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B1_valid),
		.flush(PipelineRegister_inst3$Register_inst0$reg_P1_inst0_out),
		.flush_out(Tile_X03_Y00_flush_out),
		.glb2io_1(glb2io_1_X03_Y00),
		.glb2io_17(glb2io_17_X03_Y00),
		.glb2io_17_ready(Tile_X03_Y00_glb2io_17_ready),
		.glb2io_17_valid(glb2io_17_X03_Y00_valid),
		.glb2io_1_ready(Tile_X03_Y00_glb2io_1_ready),
		.glb2io_1_valid(glb2io_1_X03_Y00_valid),
		.hi(Tile_X03_Y00_hi),
		.io2f_1(Tile_X03_Y00_io2f_1),
		.io2f_17(Tile_X03_Y00_io2f_17),
		.io2f_17_ready(Tile_X03_Y00_io2f_17_ready),
		.io2f_17_valid(Tile_X03_Y00_io2f_17_valid),
		.io2f_1_ready(Tile_X03_Y00_io2f_1_ready),
		.io2f_1_valid(Tile_X03_Y00_io2f_1_valid),
		.io2glb_1(Tile_X03_Y00_io2glb_1),
		.io2glb_17(Tile_X03_Y00_io2glb_17),
		.io2glb_17_ready(io2glb_17_X03_Y00_ready),
		.io2glb_17_valid(Tile_X03_Y00_io2glb_17_valid),
		.io2glb_1_ready(io2glb_1_X03_Y00_ready),
		.io2glb_1_valid(Tile_X03_Y00_io2glb_1_valid),
		.lo(Tile_X03_Y00_lo),
		.read_config_data(Tile_X03_Y00_read_config_data),
		.read_config_data_in(const_0_32_out),
		.reset(reset),
		.reset_out(Tile_X03_Y00_reset_out),
		.stall(self_stall_out[3:3]),
		.stall_out(Tile_X03_Y00_stall_out),
		.tile_id(Tile_X03_Y00_tile_id)
	);
	wire [15:0] Tile_X03_Y01_tile_id;
	assign Tile_X03_Y01_tile_id = {Tile_X03_Y01_lo[7], Tile_X03_Y01_lo[7], Tile_X03_Y01_lo[6], Tile_X03_Y01_lo[6], Tile_X03_Y01_lo[5], Tile_X03_Y01_lo[5], Tile_X03_Y01_hi[5], Tile_X03_Y01_hi[4], Tile_X03_Y01_lo[3], Tile_X03_Y01_lo[3], Tile_X03_Y01_lo[2], Tile_X03_Y01_lo[2], Tile_X03_Y01_lo[1], Tile_X03_Y01_lo[1], Tile_X03_Y01_lo[0], Tile_X03_Y01_hi[0]};
	Tile_MemCore Tile_X03_Y01(
		.SB_T0_EAST_SB_IN_B1(const_0_1_out),
		.SB_T0_EAST_SB_IN_B17(const_0_17_out),
		.SB_T0_EAST_SB_IN_B17_ready(Tile_X03_Y01_SB_T0_EAST_SB_IN_B17_ready),
		.SB_T0_EAST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T0_EAST_SB_IN_B1_ready(Tile_X03_Y01_SB_T0_EAST_SB_IN_B1_ready),
		.SB_T0_EAST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T0_EAST_SB_OUT_B1(Tile_X03_Y01_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_EAST_SB_OUT_B17(Tile_X03_Y01_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T0_EAST_SB_OUT_B17_valid(Tile_X03_Y01_SB_T0_EAST_SB_OUT_B17_valid),
		.SB_T0_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T0_EAST_SB_OUT_B1_valid(Tile_X03_Y01_SB_T0_EAST_SB_OUT_B1_valid),
		.SB_T0_NORTH_SB_IN_B1(Tile_X03_Y00_io2f_1),
		.SB_T0_NORTH_SB_IN_B17(Tile_X03_Y00_io2f_17),
		.SB_T0_NORTH_SB_IN_B17_ready(Tile_X03_Y01_SB_T0_NORTH_SB_IN_B17_ready),
		.SB_T0_NORTH_SB_IN_B17_valid(Tile_X03_Y00_io2f_17_valid),
		.SB_T0_NORTH_SB_IN_B1_ready(Tile_X03_Y01_SB_T0_NORTH_SB_IN_B1_ready),
		.SB_T0_NORTH_SB_IN_B1_valid(Tile_X03_Y00_io2f_1_valid),
		.SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_OUT_B17(Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_OUT_B17_ready(Tile_X03_Y00_f2io_17_ready),
		.SB_T0_NORTH_SB_OUT_B17_valid(Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B17_valid),
		.SB_T0_NORTH_SB_OUT_B1_ready(Tile_X03_Y00_f2io_1_ready),
		.SB_T0_NORTH_SB_OUT_B1_valid(Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B1_valid),
		.SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_IN_B17(Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_IN_B17_ready(Tile_X03_Y01_SB_T0_SOUTH_SB_IN_B17_ready),
		.SB_T0_SOUTH_SB_IN_B17_valid(Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B17_valid),
		.SB_T0_SOUTH_SB_IN_B1_ready(Tile_X03_Y01_SB_T0_SOUTH_SB_IN_B1_ready),
		.SB_T0_SOUTH_SB_IN_B1_valid(Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B1_valid),
		.SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_OUT_B17(Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_OUT_B17_ready(Tile_X03_Y02_SB_T0_NORTH_SB_IN_B17_ready),
		.SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B17_valid),
		.SB_T0_SOUTH_SB_OUT_B1_ready(Tile_X03_Y02_SB_T0_NORTH_SB_IN_B1_ready),
		.SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B1_valid),
		.SB_T0_WEST_SB_IN_B1(Tile_X02_Y01_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_WEST_SB_IN_B17(Tile_X02_Y01_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_WEST_SB_IN_B17_ready(Tile_X03_Y01_SB_T0_WEST_SB_IN_B17_ready),
		.SB_T0_WEST_SB_IN_B17_valid(Tile_X02_Y01_SB_T0_EAST_SB_OUT_B17_valid),
		.SB_T0_WEST_SB_IN_B1_ready(Tile_X03_Y01_SB_T0_WEST_SB_IN_B1_ready),
		.SB_T0_WEST_SB_IN_B1_valid(Tile_X02_Y01_SB_T0_EAST_SB_OUT_B1_valid),
		.SB_T0_WEST_SB_OUT_B1(Tile_X03_Y01_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_WEST_SB_OUT_B17(Tile_X03_Y01_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_WEST_SB_OUT_B17_ready(Tile_X02_Y01_SB_T0_EAST_SB_IN_B17_ready),
		.SB_T0_WEST_SB_OUT_B17_valid(Tile_X03_Y01_SB_T0_WEST_SB_OUT_B17_valid),
		.SB_T0_WEST_SB_OUT_B1_ready(Tile_X02_Y01_SB_T0_EAST_SB_IN_B1_ready),
		.SB_T0_WEST_SB_OUT_B1_valid(Tile_X03_Y01_SB_T0_WEST_SB_OUT_B1_valid),
		.SB_T1_EAST_SB_IN_B1(const_0_1_out),
		.SB_T1_EAST_SB_IN_B17(const_0_17_out),
		.SB_T1_EAST_SB_IN_B17_ready(Tile_X03_Y01_SB_T1_EAST_SB_IN_B17_ready),
		.SB_T1_EAST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T1_EAST_SB_IN_B1_ready(Tile_X03_Y01_SB_T1_EAST_SB_IN_B1_ready),
		.SB_T1_EAST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T1_EAST_SB_OUT_B1(Tile_X03_Y01_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_EAST_SB_OUT_B17(Tile_X03_Y01_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T1_EAST_SB_OUT_B17_valid(Tile_X03_Y01_SB_T1_EAST_SB_OUT_B17_valid),
		.SB_T1_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T1_EAST_SB_OUT_B1_valid(Tile_X03_Y01_SB_T1_EAST_SB_OUT_B1_valid),
		.SB_T1_NORTH_SB_IN_B1(Tile_X03_Y00_io2f_1),
		.SB_T1_NORTH_SB_IN_B17(Tile_X03_Y00_io2f_17),
		.SB_T1_NORTH_SB_IN_B17_ready(Tile_X03_Y01_SB_T1_NORTH_SB_IN_B17_ready),
		.SB_T1_NORTH_SB_IN_B17_valid(Tile_X03_Y00_io2f_17_valid),
		.SB_T1_NORTH_SB_IN_B1_ready(Tile_X03_Y01_SB_T1_NORTH_SB_IN_B1_ready),
		.SB_T1_NORTH_SB_IN_B1_valid(Tile_X03_Y00_io2f_1_valid),
		.SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y01_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_OUT_B17(Tile_X03_Y01_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T1_NORTH_SB_OUT_B17_valid(Tile_X03_Y01_SB_T1_NORTH_SB_OUT_B17_valid),
		.SB_T1_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T1_NORTH_SB_OUT_B1_valid(Tile_X03_Y01_SB_T1_NORTH_SB_OUT_B1_valid),
		.SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_IN_B17(Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_IN_B17_ready(Tile_X03_Y01_SB_T1_SOUTH_SB_IN_B17_ready),
		.SB_T1_SOUTH_SB_IN_B17_valid(Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B17_valid),
		.SB_T1_SOUTH_SB_IN_B1_ready(Tile_X03_Y01_SB_T1_SOUTH_SB_IN_B1_ready),
		.SB_T1_SOUTH_SB_IN_B1_valid(Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B1_valid),
		.SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_OUT_B17(Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_OUT_B17_ready(Tile_X03_Y02_SB_T1_NORTH_SB_IN_B17_ready),
		.SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B17_valid),
		.SB_T1_SOUTH_SB_OUT_B1_ready(Tile_X03_Y02_SB_T1_NORTH_SB_IN_B1_ready),
		.SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B1_valid),
		.SB_T1_WEST_SB_IN_B1(Tile_X02_Y01_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_WEST_SB_IN_B17(Tile_X02_Y01_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_WEST_SB_IN_B17_ready(Tile_X03_Y01_SB_T1_WEST_SB_IN_B17_ready),
		.SB_T1_WEST_SB_IN_B17_valid(Tile_X02_Y01_SB_T1_EAST_SB_OUT_B17_valid),
		.SB_T1_WEST_SB_IN_B1_ready(Tile_X03_Y01_SB_T1_WEST_SB_IN_B1_ready),
		.SB_T1_WEST_SB_IN_B1_valid(Tile_X02_Y01_SB_T1_EAST_SB_OUT_B1_valid),
		.SB_T1_WEST_SB_OUT_B1(Tile_X03_Y01_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_WEST_SB_OUT_B17(Tile_X03_Y01_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_WEST_SB_OUT_B17_ready(Tile_X02_Y01_SB_T1_EAST_SB_IN_B17_ready),
		.SB_T1_WEST_SB_OUT_B17_valid(Tile_X03_Y01_SB_T1_WEST_SB_OUT_B17_valid),
		.SB_T1_WEST_SB_OUT_B1_ready(Tile_X02_Y01_SB_T1_EAST_SB_IN_B1_ready),
		.SB_T1_WEST_SB_OUT_B1_valid(Tile_X03_Y01_SB_T1_WEST_SB_OUT_B1_valid),
		.SB_T2_EAST_SB_IN_B1(const_0_1_out),
		.SB_T2_EAST_SB_IN_B17(const_0_17_out),
		.SB_T2_EAST_SB_IN_B17_ready(Tile_X03_Y01_SB_T2_EAST_SB_IN_B17_ready),
		.SB_T2_EAST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T2_EAST_SB_IN_B1_ready(Tile_X03_Y01_SB_T2_EAST_SB_IN_B1_ready),
		.SB_T2_EAST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T2_EAST_SB_OUT_B1(Tile_X03_Y01_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_EAST_SB_OUT_B17(Tile_X03_Y01_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T2_EAST_SB_OUT_B17_valid(Tile_X03_Y01_SB_T2_EAST_SB_OUT_B17_valid),
		.SB_T2_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T2_EAST_SB_OUT_B1_valid(Tile_X03_Y01_SB_T2_EAST_SB_OUT_B1_valid),
		.SB_T2_NORTH_SB_IN_B1(Tile_X03_Y00_io2f_1),
		.SB_T2_NORTH_SB_IN_B17(Tile_X03_Y00_io2f_17),
		.SB_T2_NORTH_SB_IN_B17_ready(Tile_X03_Y01_SB_T2_NORTH_SB_IN_B17_ready),
		.SB_T2_NORTH_SB_IN_B17_valid(Tile_X03_Y00_io2f_17_valid),
		.SB_T2_NORTH_SB_IN_B1_ready(Tile_X03_Y01_SB_T2_NORTH_SB_IN_B1_ready),
		.SB_T2_NORTH_SB_IN_B1_valid(Tile_X03_Y00_io2f_1_valid),
		.SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y01_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_OUT_B17(Tile_X03_Y01_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T2_NORTH_SB_OUT_B17_valid(Tile_X03_Y01_SB_T2_NORTH_SB_OUT_B17_valid),
		.SB_T2_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T2_NORTH_SB_OUT_B1_valid(Tile_X03_Y01_SB_T2_NORTH_SB_OUT_B1_valid),
		.SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_IN_B17(Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_IN_B17_ready(Tile_X03_Y01_SB_T2_SOUTH_SB_IN_B17_ready),
		.SB_T2_SOUTH_SB_IN_B17_valid(Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B17_valid),
		.SB_T2_SOUTH_SB_IN_B1_ready(Tile_X03_Y01_SB_T2_SOUTH_SB_IN_B1_ready),
		.SB_T2_SOUTH_SB_IN_B1_valid(Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B1_valid),
		.SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_OUT_B17(Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_OUT_B17_ready(Tile_X03_Y02_SB_T2_NORTH_SB_IN_B17_ready),
		.SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B17_valid),
		.SB_T2_SOUTH_SB_OUT_B1_ready(Tile_X03_Y02_SB_T2_NORTH_SB_IN_B1_ready),
		.SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B1_valid),
		.SB_T2_WEST_SB_IN_B1(Tile_X02_Y01_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_WEST_SB_IN_B17(Tile_X02_Y01_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_WEST_SB_IN_B17_ready(Tile_X03_Y01_SB_T2_WEST_SB_IN_B17_ready),
		.SB_T2_WEST_SB_IN_B17_valid(Tile_X02_Y01_SB_T2_EAST_SB_OUT_B17_valid),
		.SB_T2_WEST_SB_IN_B1_ready(Tile_X03_Y01_SB_T2_WEST_SB_IN_B1_ready),
		.SB_T2_WEST_SB_IN_B1_valid(Tile_X02_Y01_SB_T2_EAST_SB_OUT_B1_valid),
		.SB_T2_WEST_SB_OUT_B1(Tile_X03_Y01_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_WEST_SB_OUT_B17(Tile_X03_Y01_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_WEST_SB_OUT_B17_ready(Tile_X02_Y01_SB_T2_EAST_SB_IN_B17_ready),
		.SB_T2_WEST_SB_OUT_B17_valid(Tile_X03_Y01_SB_T2_WEST_SB_OUT_B17_valid),
		.SB_T2_WEST_SB_OUT_B1_ready(Tile_X02_Y01_SB_T2_EAST_SB_IN_B1_ready),
		.SB_T2_WEST_SB_OUT_B1_valid(Tile_X03_Y01_SB_T2_WEST_SB_OUT_B1_valid),
		.SB_T3_EAST_SB_IN_B1(const_0_1_out),
		.SB_T3_EAST_SB_IN_B17(const_0_17_out),
		.SB_T3_EAST_SB_IN_B17_ready(Tile_X03_Y01_SB_T3_EAST_SB_IN_B17_ready),
		.SB_T3_EAST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T3_EAST_SB_IN_B1_ready(Tile_X03_Y01_SB_T3_EAST_SB_IN_B1_ready),
		.SB_T3_EAST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T3_EAST_SB_OUT_B1(Tile_X03_Y01_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_EAST_SB_OUT_B17(Tile_X03_Y01_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T3_EAST_SB_OUT_B17_valid(Tile_X03_Y01_SB_T3_EAST_SB_OUT_B17_valid),
		.SB_T3_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T3_EAST_SB_OUT_B1_valid(Tile_X03_Y01_SB_T3_EAST_SB_OUT_B1_valid),
		.SB_T3_NORTH_SB_IN_B1(Tile_X03_Y00_io2f_1),
		.SB_T3_NORTH_SB_IN_B17(Tile_X03_Y00_io2f_17),
		.SB_T3_NORTH_SB_IN_B17_ready(Tile_X03_Y01_SB_T3_NORTH_SB_IN_B17_ready),
		.SB_T3_NORTH_SB_IN_B17_valid(Tile_X03_Y00_io2f_17_valid),
		.SB_T3_NORTH_SB_IN_B1_ready(Tile_X03_Y01_SB_T3_NORTH_SB_IN_B1_ready),
		.SB_T3_NORTH_SB_IN_B1_valid(Tile_X03_Y00_io2f_1_valid),
		.SB_T3_NORTH_SB_OUT_B1(Tile_X03_Y01_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_OUT_B17(Tile_X03_Y01_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T3_NORTH_SB_OUT_B17_valid(Tile_X03_Y01_SB_T3_NORTH_SB_OUT_B17_valid),
		.SB_T3_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T3_NORTH_SB_OUT_B1_valid(Tile_X03_Y01_SB_T3_NORTH_SB_OUT_B1_valid),
		.SB_T3_SOUTH_SB_IN_B1(Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_IN_B17(Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_IN_B17_ready(Tile_X03_Y01_SB_T3_SOUTH_SB_IN_B17_ready),
		.SB_T3_SOUTH_SB_IN_B17_valid(Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B17_valid),
		.SB_T3_SOUTH_SB_IN_B1_ready(Tile_X03_Y01_SB_T3_SOUTH_SB_IN_B1_ready),
		.SB_T3_SOUTH_SB_IN_B1_valid(Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B1_valid),
		.SB_T3_SOUTH_SB_OUT_B1(Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_OUT_B17(Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_OUT_B17_ready(Tile_X03_Y02_SB_T3_NORTH_SB_IN_B17_ready),
		.SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B17_valid),
		.SB_T3_SOUTH_SB_OUT_B1_ready(Tile_X03_Y02_SB_T3_NORTH_SB_IN_B1_ready),
		.SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B1_valid),
		.SB_T3_WEST_SB_IN_B1(Tile_X02_Y01_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_WEST_SB_IN_B17(Tile_X02_Y01_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_WEST_SB_IN_B17_ready(Tile_X03_Y01_SB_T3_WEST_SB_IN_B17_ready),
		.SB_T3_WEST_SB_IN_B17_valid(Tile_X02_Y01_SB_T3_EAST_SB_OUT_B17_valid),
		.SB_T3_WEST_SB_IN_B1_ready(Tile_X03_Y01_SB_T3_WEST_SB_IN_B1_ready),
		.SB_T3_WEST_SB_IN_B1_valid(Tile_X02_Y01_SB_T3_EAST_SB_OUT_B1_valid),
		.SB_T3_WEST_SB_OUT_B1(Tile_X03_Y01_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_WEST_SB_OUT_B17(Tile_X03_Y01_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_WEST_SB_OUT_B17_ready(Tile_X02_Y01_SB_T3_EAST_SB_IN_B17_ready),
		.SB_T3_WEST_SB_OUT_B17_valid(Tile_X03_Y01_SB_T3_WEST_SB_OUT_B17_valid),
		.SB_T3_WEST_SB_OUT_B1_ready(Tile_X02_Y01_SB_T3_EAST_SB_IN_B1_ready),
		.SB_T3_WEST_SB_OUT_B1_valid(Tile_X03_Y01_SB_T3_WEST_SB_OUT_B1_valid),
		.SB_T4_EAST_SB_IN_B1(const_0_1_out),
		.SB_T4_EAST_SB_IN_B17(const_0_17_out),
		.SB_T4_EAST_SB_IN_B17_ready(Tile_X03_Y01_SB_T4_EAST_SB_IN_B17_ready),
		.SB_T4_EAST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T4_EAST_SB_IN_B1_ready(Tile_X03_Y01_SB_T4_EAST_SB_IN_B1_ready),
		.SB_T4_EAST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T4_EAST_SB_OUT_B1(Tile_X03_Y01_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_EAST_SB_OUT_B17(Tile_X03_Y01_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T4_EAST_SB_OUT_B17_valid(Tile_X03_Y01_SB_T4_EAST_SB_OUT_B17_valid),
		.SB_T4_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T4_EAST_SB_OUT_B1_valid(Tile_X03_Y01_SB_T4_EAST_SB_OUT_B1_valid),
		.SB_T4_NORTH_SB_IN_B1(Tile_X03_Y00_io2f_1),
		.SB_T4_NORTH_SB_IN_B17(Tile_X03_Y00_io2f_17),
		.SB_T4_NORTH_SB_IN_B17_ready(Tile_X03_Y01_SB_T4_NORTH_SB_IN_B17_ready),
		.SB_T4_NORTH_SB_IN_B17_valid(Tile_X03_Y00_io2f_17_valid),
		.SB_T4_NORTH_SB_IN_B1_ready(Tile_X03_Y01_SB_T4_NORTH_SB_IN_B1_ready),
		.SB_T4_NORTH_SB_IN_B1_valid(Tile_X03_Y00_io2f_1_valid),
		.SB_T4_NORTH_SB_OUT_B1(Tile_X03_Y01_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_OUT_B17(Tile_X03_Y01_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T4_NORTH_SB_OUT_B17_valid(Tile_X03_Y01_SB_T4_NORTH_SB_OUT_B17_valid),
		.SB_T4_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T4_NORTH_SB_OUT_B1_valid(Tile_X03_Y01_SB_T4_NORTH_SB_OUT_B1_valid),
		.SB_T4_SOUTH_SB_IN_B1(Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_IN_B17(Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_IN_B17_ready(Tile_X03_Y01_SB_T4_SOUTH_SB_IN_B17_ready),
		.SB_T4_SOUTH_SB_IN_B17_valid(Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B17_valid),
		.SB_T4_SOUTH_SB_IN_B1_ready(Tile_X03_Y01_SB_T4_SOUTH_SB_IN_B1_ready),
		.SB_T4_SOUTH_SB_IN_B1_valid(Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B1_valid),
		.SB_T4_SOUTH_SB_OUT_B1(Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_OUT_B17(Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_OUT_B17_ready(Tile_X03_Y02_SB_T4_NORTH_SB_IN_B17_ready),
		.SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B17_valid),
		.SB_T4_SOUTH_SB_OUT_B1_ready(Tile_X03_Y02_SB_T4_NORTH_SB_IN_B1_ready),
		.SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B1_valid),
		.SB_T4_WEST_SB_IN_B1(Tile_X02_Y01_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_WEST_SB_IN_B17(Tile_X02_Y01_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_WEST_SB_IN_B17_ready(Tile_X03_Y01_SB_T4_WEST_SB_IN_B17_ready),
		.SB_T4_WEST_SB_IN_B17_valid(Tile_X02_Y01_SB_T4_EAST_SB_OUT_B17_valid),
		.SB_T4_WEST_SB_IN_B1_ready(Tile_X03_Y01_SB_T4_WEST_SB_IN_B1_ready),
		.SB_T4_WEST_SB_IN_B1_valid(Tile_X02_Y01_SB_T4_EAST_SB_OUT_B1_valid),
		.SB_T4_WEST_SB_OUT_B1(Tile_X03_Y01_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_WEST_SB_OUT_B17(Tile_X03_Y01_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_WEST_SB_OUT_B17_ready(Tile_X02_Y01_SB_T4_EAST_SB_IN_B17_ready),
		.SB_T4_WEST_SB_OUT_B17_valid(Tile_X03_Y01_SB_T4_WEST_SB_OUT_B17_valid),
		.SB_T4_WEST_SB_OUT_B1_ready(Tile_X02_Y01_SB_T4_EAST_SB_IN_B1_ready),
		.SB_T4_WEST_SB_OUT_B1_valid(Tile_X03_Y01_SB_T4_WEST_SB_OUT_B1_valid),
		.clk(Tile_X02_Y01_clk_pass_through_out_right),
		.clk_out(Tile_X03_Y01_clk_out),
		.config_config_addr(Tile_X03_Y00_config_out_config_addr),
		.config_config_data(Tile_X03_Y00_config_out_config_data),
		.config_out_config_addr(Tile_X03_Y01_config_out_config_addr),
		.config_out_config_data(Tile_X03_Y01_config_out_config_data),
		.config_out_read(Tile_X03_Y01_config_out_read),
		.config_out_write(Tile_X03_Y01_config_out_write),
		.config_read(Tile_X03_Y00_config_out_read),
		.config_write(Tile_X03_Y00_config_out_write),
		.flush(Tile_X03_Y00_flush_out),
		.flush_out(Tile_X03_Y01_flush_out),
		.hi(Tile_X03_Y01_hi),
		.lo(Tile_X03_Y01_lo),
		.read_config_data(Tile_X03_Y01_read_config_data),
		.read_config_data_in(Tile_X03_Y00_read_config_data),
		.reset(Tile_X03_Y00_reset_out),
		.reset_out(Tile_X03_Y01_reset_out),
		.stall(Tile_X03_Y00_stall_out),
		.stall_out(Tile_X03_Y01_stall_out),
		.tile_id(Tile_X03_Y01_tile_id)
	);
	wire [15:0] Tile_X03_Y02_tile_id;
	assign Tile_X03_Y02_tile_id = {Tile_X03_Y02_lo[7], Tile_X03_Y02_lo[7], Tile_X03_Y02_lo[6], Tile_X03_Y02_lo[6], Tile_X03_Y02_lo[5], Tile_X03_Y02_lo[5], Tile_X03_Y02_hi[5], Tile_X03_Y02_hi[4], Tile_X03_Y02_lo[3], Tile_X03_Y02_lo[3], Tile_X03_Y02_lo[2], Tile_X03_Y02_lo[2], Tile_X03_Y02_lo[1], Tile_X03_Y02_lo[1], Tile_X03_Y02_hi[1], Tile_X03_Y02_lo[0]};
	Tile_MemCore Tile_X03_Y02(
		.SB_T0_EAST_SB_IN_B1(const_0_1_out),
		.SB_T0_EAST_SB_IN_B17(const_0_17_out),
		.SB_T0_EAST_SB_IN_B17_ready(Tile_X03_Y02_SB_T0_EAST_SB_IN_B17_ready),
		.SB_T0_EAST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T0_EAST_SB_IN_B1_ready(Tile_X03_Y02_SB_T0_EAST_SB_IN_B1_ready),
		.SB_T0_EAST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T0_EAST_SB_OUT_B1(Tile_X03_Y02_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_EAST_SB_OUT_B17(Tile_X03_Y02_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T0_EAST_SB_OUT_B17_valid(Tile_X03_Y02_SB_T0_EAST_SB_OUT_B17_valid),
		.SB_T0_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T0_EAST_SB_OUT_B1_valid(Tile_X03_Y02_SB_T0_EAST_SB_OUT_B1_valid),
		.SB_T0_NORTH_SB_IN_B1(Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_IN_B17(Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_IN_B17_ready(Tile_X03_Y02_SB_T0_NORTH_SB_IN_B17_ready),
		.SB_T0_NORTH_SB_IN_B17_valid(Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B17_valid),
		.SB_T0_NORTH_SB_IN_B1_ready(Tile_X03_Y02_SB_T0_NORTH_SB_IN_B1_ready),
		.SB_T0_NORTH_SB_IN_B1_valid(Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B1_valid),
		.SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_OUT_B17(Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_OUT_B17_ready(Tile_X03_Y01_SB_T0_SOUTH_SB_IN_B17_ready),
		.SB_T0_NORTH_SB_OUT_B17_valid(Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B17_valid),
		.SB_T0_NORTH_SB_OUT_B1_ready(Tile_X03_Y01_SB_T0_SOUTH_SB_IN_B1_ready),
		.SB_T0_NORTH_SB_OUT_B1_valid(Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B1_valid),
		.SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_IN_B17(Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_IN_B17_ready(Tile_X03_Y02_SB_T0_SOUTH_SB_IN_B17_ready),
		.SB_T0_SOUTH_SB_IN_B17_valid(Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B17_valid),
		.SB_T0_SOUTH_SB_IN_B1_ready(Tile_X03_Y02_SB_T0_SOUTH_SB_IN_B1_ready),
		.SB_T0_SOUTH_SB_IN_B1_valid(Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B1_valid),
		.SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_OUT_B17(Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_OUT_B17_ready(Tile_X03_Y03_SB_T0_NORTH_SB_IN_B17_ready),
		.SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B17_valid),
		.SB_T0_SOUTH_SB_OUT_B1_ready(Tile_X03_Y03_SB_T0_NORTH_SB_IN_B1_ready),
		.SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B1_valid),
		.SB_T0_WEST_SB_IN_B1(Tile_X02_Y02_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_WEST_SB_IN_B17(Tile_X02_Y02_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_WEST_SB_IN_B17_ready(Tile_X03_Y02_SB_T0_WEST_SB_IN_B17_ready),
		.SB_T0_WEST_SB_IN_B17_valid(Tile_X02_Y02_SB_T0_EAST_SB_OUT_B17_valid),
		.SB_T0_WEST_SB_IN_B1_ready(Tile_X03_Y02_SB_T0_WEST_SB_IN_B1_ready),
		.SB_T0_WEST_SB_IN_B1_valid(Tile_X02_Y02_SB_T0_EAST_SB_OUT_B1_valid),
		.SB_T0_WEST_SB_OUT_B1(Tile_X03_Y02_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_WEST_SB_OUT_B17(Tile_X03_Y02_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_WEST_SB_OUT_B17_ready(Tile_X02_Y02_SB_T0_EAST_SB_IN_B17_ready),
		.SB_T0_WEST_SB_OUT_B17_valid(Tile_X03_Y02_SB_T0_WEST_SB_OUT_B17_valid),
		.SB_T0_WEST_SB_OUT_B1_ready(Tile_X02_Y02_SB_T0_EAST_SB_IN_B1_ready),
		.SB_T0_WEST_SB_OUT_B1_valid(Tile_X03_Y02_SB_T0_WEST_SB_OUT_B1_valid),
		.SB_T1_EAST_SB_IN_B1(const_0_1_out),
		.SB_T1_EAST_SB_IN_B17(const_0_17_out),
		.SB_T1_EAST_SB_IN_B17_ready(Tile_X03_Y02_SB_T1_EAST_SB_IN_B17_ready),
		.SB_T1_EAST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T1_EAST_SB_IN_B1_ready(Tile_X03_Y02_SB_T1_EAST_SB_IN_B1_ready),
		.SB_T1_EAST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T1_EAST_SB_OUT_B1(Tile_X03_Y02_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_EAST_SB_OUT_B17(Tile_X03_Y02_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T1_EAST_SB_OUT_B17_valid(Tile_X03_Y02_SB_T1_EAST_SB_OUT_B17_valid),
		.SB_T1_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T1_EAST_SB_OUT_B1_valid(Tile_X03_Y02_SB_T1_EAST_SB_OUT_B1_valid),
		.SB_T1_NORTH_SB_IN_B1(Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_IN_B17(Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_IN_B17_ready(Tile_X03_Y02_SB_T1_NORTH_SB_IN_B17_ready),
		.SB_T1_NORTH_SB_IN_B17_valid(Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B17_valid),
		.SB_T1_NORTH_SB_IN_B1_ready(Tile_X03_Y02_SB_T1_NORTH_SB_IN_B1_ready),
		.SB_T1_NORTH_SB_IN_B1_valid(Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B1_valid),
		.SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_OUT_B17(Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_OUT_B17_ready(Tile_X03_Y01_SB_T1_SOUTH_SB_IN_B17_ready),
		.SB_T1_NORTH_SB_OUT_B17_valid(Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B17_valid),
		.SB_T1_NORTH_SB_OUT_B1_ready(Tile_X03_Y01_SB_T1_SOUTH_SB_IN_B1_ready),
		.SB_T1_NORTH_SB_OUT_B1_valid(Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B1_valid),
		.SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_IN_B17(Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_IN_B17_ready(Tile_X03_Y02_SB_T1_SOUTH_SB_IN_B17_ready),
		.SB_T1_SOUTH_SB_IN_B17_valid(Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B17_valid),
		.SB_T1_SOUTH_SB_IN_B1_ready(Tile_X03_Y02_SB_T1_SOUTH_SB_IN_B1_ready),
		.SB_T1_SOUTH_SB_IN_B1_valid(Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B1_valid),
		.SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_OUT_B17(Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_OUT_B17_ready(Tile_X03_Y03_SB_T1_NORTH_SB_IN_B17_ready),
		.SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B17_valid),
		.SB_T1_SOUTH_SB_OUT_B1_ready(Tile_X03_Y03_SB_T1_NORTH_SB_IN_B1_ready),
		.SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B1_valid),
		.SB_T1_WEST_SB_IN_B1(Tile_X02_Y02_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_WEST_SB_IN_B17(Tile_X02_Y02_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_WEST_SB_IN_B17_ready(Tile_X03_Y02_SB_T1_WEST_SB_IN_B17_ready),
		.SB_T1_WEST_SB_IN_B17_valid(Tile_X02_Y02_SB_T1_EAST_SB_OUT_B17_valid),
		.SB_T1_WEST_SB_IN_B1_ready(Tile_X03_Y02_SB_T1_WEST_SB_IN_B1_ready),
		.SB_T1_WEST_SB_IN_B1_valid(Tile_X02_Y02_SB_T1_EAST_SB_OUT_B1_valid),
		.SB_T1_WEST_SB_OUT_B1(Tile_X03_Y02_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_WEST_SB_OUT_B17(Tile_X03_Y02_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_WEST_SB_OUT_B17_ready(Tile_X02_Y02_SB_T1_EAST_SB_IN_B17_ready),
		.SB_T1_WEST_SB_OUT_B17_valid(Tile_X03_Y02_SB_T1_WEST_SB_OUT_B17_valid),
		.SB_T1_WEST_SB_OUT_B1_ready(Tile_X02_Y02_SB_T1_EAST_SB_IN_B1_ready),
		.SB_T1_WEST_SB_OUT_B1_valid(Tile_X03_Y02_SB_T1_WEST_SB_OUT_B1_valid),
		.SB_T2_EAST_SB_IN_B1(const_0_1_out),
		.SB_T2_EAST_SB_IN_B17(const_0_17_out),
		.SB_T2_EAST_SB_IN_B17_ready(Tile_X03_Y02_SB_T2_EAST_SB_IN_B17_ready),
		.SB_T2_EAST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T2_EAST_SB_IN_B1_ready(Tile_X03_Y02_SB_T2_EAST_SB_IN_B1_ready),
		.SB_T2_EAST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T2_EAST_SB_OUT_B1(Tile_X03_Y02_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_EAST_SB_OUT_B17(Tile_X03_Y02_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T2_EAST_SB_OUT_B17_valid(Tile_X03_Y02_SB_T2_EAST_SB_OUT_B17_valid),
		.SB_T2_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T2_EAST_SB_OUT_B1_valid(Tile_X03_Y02_SB_T2_EAST_SB_OUT_B1_valid),
		.SB_T2_NORTH_SB_IN_B1(Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_IN_B17(Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_IN_B17_ready(Tile_X03_Y02_SB_T2_NORTH_SB_IN_B17_ready),
		.SB_T2_NORTH_SB_IN_B17_valid(Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B17_valid),
		.SB_T2_NORTH_SB_IN_B1_ready(Tile_X03_Y02_SB_T2_NORTH_SB_IN_B1_ready),
		.SB_T2_NORTH_SB_IN_B1_valid(Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B1_valid),
		.SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_OUT_B17(Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_OUT_B17_ready(Tile_X03_Y01_SB_T2_SOUTH_SB_IN_B17_ready),
		.SB_T2_NORTH_SB_OUT_B17_valid(Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B17_valid),
		.SB_T2_NORTH_SB_OUT_B1_ready(Tile_X03_Y01_SB_T2_SOUTH_SB_IN_B1_ready),
		.SB_T2_NORTH_SB_OUT_B1_valid(Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B1_valid),
		.SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_IN_B17(Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_IN_B17_ready(Tile_X03_Y02_SB_T2_SOUTH_SB_IN_B17_ready),
		.SB_T2_SOUTH_SB_IN_B17_valid(Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B17_valid),
		.SB_T2_SOUTH_SB_IN_B1_ready(Tile_X03_Y02_SB_T2_SOUTH_SB_IN_B1_ready),
		.SB_T2_SOUTH_SB_IN_B1_valid(Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B1_valid),
		.SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_OUT_B17(Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_OUT_B17_ready(Tile_X03_Y03_SB_T2_NORTH_SB_IN_B17_ready),
		.SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B17_valid),
		.SB_T2_SOUTH_SB_OUT_B1_ready(Tile_X03_Y03_SB_T2_NORTH_SB_IN_B1_ready),
		.SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B1_valid),
		.SB_T2_WEST_SB_IN_B1(Tile_X02_Y02_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_WEST_SB_IN_B17(Tile_X02_Y02_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_WEST_SB_IN_B17_ready(Tile_X03_Y02_SB_T2_WEST_SB_IN_B17_ready),
		.SB_T2_WEST_SB_IN_B17_valid(Tile_X02_Y02_SB_T2_EAST_SB_OUT_B17_valid),
		.SB_T2_WEST_SB_IN_B1_ready(Tile_X03_Y02_SB_T2_WEST_SB_IN_B1_ready),
		.SB_T2_WEST_SB_IN_B1_valid(Tile_X02_Y02_SB_T2_EAST_SB_OUT_B1_valid),
		.SB_T2_WEST_SB_OUT_B1(Tile_X03_Y02_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_WEST_SB_OUT_B17(Tile_X03_Y02_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_WEST_SB_OUT_B17_ready(Tile_X02_Y02_SB_T2_EAST_SB_IN_B17_ready),
		.SB_T2_WEST_SB_OUT_B17_valid(Tile_X03_Y02_SB_T2_WEST_SB_OUT_B17_valid),
		.SB_T2_WEST_SB_OUT_B1_ready(Tile_X02_Y02_SB_T2_EAST_SB_IN_B1_ready),
		.SB_T2_WEST_SB_OUT_B1_valid(Tile_X03_Y02_SB_T2_WEST_SB_OUT_B1_valid),
		.SB_T3_EAST_SB_IN_B1(const_0_1_out),
		.SB_T3_EAST_SB_IN_B17(const_0_17_out),
		.SB_T3_EAST_SB_IN_B17_ready(Tile_X03_Y02_SB_T3_EAST_SB_IN_B17_ready),
		.SB_T3_EAST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T3_EAST_SB_IN_B1_ready(Tile_X03_Y02_SB_T3_EAST_SB_IN_B1_ready),
		.SB_T3_EAST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T3_EAST_SB_OUT_B1(Tile_X03_Y02_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_EAST_SB_OUT_B17(Tile_X03_Y02_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T3_EAST_SB_OUT_B17_valid(Tile_X03_Y02_SB_T3_EAST_SB_OUT_B17_valid),
		.SB_T3_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T3_EAST_SB_OUT_B1_valid(Tile_X03_Y02_SB_T3_EAST_SB_OUT_B1_valid),
		.SB_T3_NORTH_SB_IN_B1(Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_IN_B17(Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_IN_B17_ready(Tile_X03_Y02_SB_T3_NORTH_SB_IN_B17_ready),
		.SB_T3_NORTH_SB_IN_B17_valid(Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B17_valid),
		.SB_T3_NORTH_SB_IN_B1_ready(Tile_X03_Y02_SB_T3_NORTH_SB_IN_B1_ready),
		.SB_T3_NORTH_SB_IN_B1_valid(Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B1_valid),
		.SB_T3_NORTH_SB_OUT_B1(Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_OUT_B17(Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_OUT_B17_ready(Tile_X03_Y01_SB_T3_SOUTH_SB_IN_B17_ready),
		.SB_T3_NORTH_SB_OUT_B17_valid(Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B17_valid),
		.SB_T3_NORTH_SB_OUT_B1_ready(Tile_X03_Y01_SB_T3_SOUTH_SB_IN_B1_ready),
		.SB_T3_NORTH_SB_OUT_B1_valid(Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B1_valid),
		.SB_T3_SOUTH_SB_IN_B1(Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_IN_B17(Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_IN_B17_ready(Tile_X03_Y02_SB_T3_SOUTH_SB_IN_B17_ready),
		.SB_T3_SOUTH_SB_IN_B17_valid(Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B17_valid),
		.SB_T3_SOUTH_SB_IN_B1_ready(Tile_X03_Y02_SB_T3_SOUTH_SB_IN_B1_ready),
		.SB_T3_SOUTH_SB_IN_B1_valid(Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B1_valid),
		.SB_T3_SOUTH_SB_OUT_B1(Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_OUT_B17(Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_OUT_B17_ready(Tile_X03_Y03_SB_T3_NORTH_SB_IN_B17_ready),
		.SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B17_valid),
		.SB_T3_SOUTH_SB_OUT_B1_ready(Tile_X03_Y03_SB_T3_NORTH_SB_IN_B1_ready),
		.SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B1_valid),
		.SB_T3_WEST_SB_IN_B1(Tile_X02_Y02_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_WEST_SB_IN_B17(Tile_X02_Y02_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_WEST_SB_IN_B17_ready(Tile_X03_Y02_SB_T3_WEST_SB_IN_B17_ready),
		.SB_T3_WEST_SB_IN_B17_valid(Tile_X02_Y02_SB_T3_EAST_SB_OUT_B17_valid),
		.SB_T3_WEST_SB_IN_B1_ready(Tile_X03_Y02_SB_T3_WEST_SB_IN_B1_ready),
		.SB_T3_WEST_SB_IN_B1_valid(Tile_X02_Y02_SB_T3_EAST_SB_OUT_B1_valid),
		.SB_T3_WEST_SB_OUT_B1(Tile_X03_Y02_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_WEST_SB_OUT_B17(Tile_X03_Y02_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_WEST_SB_OUT_B17_ready(Tile_X02_Y02_SB_T3_EAST_SB_IN_B17_ready),
		.SB_T3_WEST_SB_OUT_B17_valid(Tile_X03_Y02_SB_T3_WEST_SB_OUT_B17_valid),
		.SB_T3_WEST_SB_OUT_B1_ready(Tile_X02_Y02_SB_T3_EAST_SB_IN_B1_ready),
		.SB_T3_WEST_SB_OUT_B1_valid(Tile_X03_Y02_SB_T3_WEST_SB_OUT_B1_valid),
		.SB_T4_EAST_SB_IN_B1(const_0_1_out),
		.SB_T4_EAST_SB_IN_B17(const_0_17_out),
		.SB_T4_EAST_SB_IN_B17_ready(Tile_X03_Y02_SB_T4_EAST_SB_IN_B17_ready),
		.SB_T4_EAST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T4_EAST_SB_IN_B1_ready(Tile_X03_Y02_SB_T4_EAST_SB_IN_B1_ready),
		.SB_T4_EAST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T4_EAST_SB_OUT_B1(Tile_X03_Y02_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_EAST_SB_OUT_B17(Tile_X03_Y02_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T4_EAST_SB_OUT_B17_valid(Tile_X03_Y02_SB_T4_EAST_SB_OUT_B17_valid),
		.SB_T4_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T4_EAST_SB_OUT_B1_valid(Tile_X03_Y02_SB_T4_EAST_SB_OUT_B1_valid),
		.SB_T4_NORTH_SB_IN_B1(Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_IN_B17(Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_IN_B17_ready(Tile_X03_Y02_SB_T4_NORTH_SB_IN_B17_ready),
		.SB_T4_NORTH_SB_IN_B17_valid(Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B17_valid),
		.SB_T4_NORTH_SB_IN_B1_ready(Tile_X03_Y02_SB_T4_NORTH_SB_IN_B1_ready),
		.SB_T4_NORTH_SB_IN_B1_valid(Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B1_valid),
		.SB_T4_NORTH_SB_OUT_B1(Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_OUT_B17(Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_OUT_B17_ready(Tile_X03_Y01_SB_T4_SOUTH_SB_IN_B17_ready),
		.SB_T4_NORTH_SB_OUT_B17_valid(Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B17_valid),
		.SB_T4_NORTH_SB_OUT_B1_ready(Tile_X03_Y01_SB_T4_SOUTH_SB_IN_B1_ready),
		.SB_T4_NORTH_SB_OUT_B1_valid(Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B1_valid),
		.SB_T4_SOUTH_SB_IN_B1(Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_IN_B17(Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_IN_B17_ready(Tile_X03_Y02_SB_T4_SOUTH_SB_IN_B17_ready),
		.SB_T4_SOUTH_SB_IN_B17_valid(Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B17_valid),
		.SB_T4_SOUTH_SB_IN_B1_ready(Tile_X03_Y02_SB_T4_SOUTH_SB_IN_B1_ready),
		.SB_T4_SOUTH_SB_IN_B1_valid(Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B1_valid),
		.SB_T4_SOUTH_SB_OUT_B1(Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_OUT_B17(Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_OUT_B17_ready(Tile_X03_Y03_SB_T4_NORTH_SB_IN_B17_ready),
		.SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B17_valid),
		.SB_T4_SOUTH_SB_OUT_B1_ready(Tile_X03_Y03_SB_T4_NORTH_SB_IN_B1_ready),
		.SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B1_valid),
		.SB_T4_WEST_SB_IN_B1(Tile_X02_Y02_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_WEST_SB_IN_B17(Tile_X02_Y02_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_WEST_SB_IN_B17_ready(Tile_X03_Y02_SB_T4_WEST_SB_IN_B17_ready),
		.SB_T4_WEST_SB_IN_B17_valid(Tile_X02_Y02_SB_T4_EAST_SB_OUT_B17_valid),
		.SB_T4_WEST_SB_IN_B1_ready(Tile_X03_Y02_SB_T4_WEST_SB_IN_B1_ready),
		.SB_T4_WEST_SB_IN_B1_valid(Tile_X02_Y02_SB_T4_EAST_SB_OUT_B1_valid),
		.SB_T4_WEST_SB_OUT_B1(Tile_X03_Y02_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_WEST_SB_OUT_B17(Tile_X03_Y02_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_WEST_SB_OUT_B17_ready(Tile_X02_Y02_SB_T4_EAST_SB_IN_B17_ready),
		.SB_T4_WEST_SB_OUT_B17_valid(Tile_X03_Y02_SB_T4_WEST_SB_OUT_B17_valid),
		.SB_T4_WEST_SB_OUT_B1_ready(Tile_X02_Y02_SB_T4_EAST_SB_IN_B1_ready),
		.SB_T4_WEST_SB_OUT_B1_valid(Tile_X03_Y02_SB_T4_WEST_SB_OUT_B1_valid),
		.clk(Tile_X02_Y02_clk_pass_through_out_right),
		.clk_out(Tile_X03_Y02_clk_out),
		.config_config_addr(Tile_X03_Y01_config_out_config_addr),
		.config_config_data(Tile_X03_Y01_config_out_config_data),
		.config_out_config_addr(Tile_X03_Y02_config_out_config_addr),
		.config_out_config_data(Tile_X03_Y02_config_out_config_data),
		.config_out_read(Tile_X03_Y02_config_out_read),
		.config_out_write(Tile_X03_Y02_config_out_write),
		.config_read(Tile_X03_Y01_config_out_read),
		.config_write(Tile_X03_Y01_config_out_write),
		.flush(Tile_X03_Y01_flush_out),
		.flush_out(Tile_X03_Y02_flush_out),
		.hi(Tile_X03_Y02_hi),
		.lo(Tile_X03_Y02_lo),
		.read_config_data(Tile_X03_Y02_read_config_data),
		.read_config_data_in(Tile_X03_Y01_read_config_data),
		.reset(Tile_X03_Y01_reset_out),
		.reset_out(Tile_X03_Y02_reset_out),
		.stall(Tile_X03_Y01_stall_out),
		.stall_out(Tile_X03_Y02_stall_out),
		.tile_id(Tile_X03_Y02_tile_id)
	);
	wire [15:0] Tile_X03_Y03_tile_id;
	assign Tile_X03_Y03_tile_id = {Tile_X03_Y03_lo[7], Tile_X03_Y03_lo[7], Tile_X03_Y03_lo[6], Tile_X03_Y03_lo[6], Tile_X03_Y03_lo[5], Tile_X03_Y03_lo[5], Tile_X03_Y03_hi[5], Tile_X03_Y03_hi[4], Tile_X03_Y03_lo[3], Tile_X03_Y03_lo[3], Tile_X03_Y03_lo[2], Tile_X03_Y03_lo[2], Tile_X03_Y03_lo[1], Tile_X03_Y03_lo[1], Tile_X03_Y03_hi[1], Tile_X03_Y03_hi[0]};
	Tile_MemCore Tile_X03_Y03(
		.SB_T0_EAST_SB_IN_B1(const_0_1_out),
		.SB_T0_EAST_SB_IN_B17(const_0_17_out),
		.SB_T0_EAST_SB_IN_B17_ready(Tile_X03_Y03_SB_T0_EAST_SB_IN_B17_ready),
		.SB_T0_EAST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T0_EAST_SB_IN_B1_ready(Tile_X03_Y03_SB_T0_EAST_SB_IN_B1_ready),
		.SB_T0_EAST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T0_EAST_SB_OUT_B1(Tile_X03_Y03_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_EAST_SB_OUT_B17(Tile_X03_Y03_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T0_EAST_SB_OUT_B17_valid(Tile_X03_Y03_SB_T0_EAST_SB_OUT_B17_valid),
		.SB_T0_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T0_EAST_SB_OUT_B1_valid(Tile_X03_Y03_SB_T0_EAST_SB_OUT_B1_valid),
		.SB_T0_NORTH_SB_IN_B1(Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_IN_B17(Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_IN_B17_ready(Tile_X03_Y03_SB_T0_NORTH_SB_IN_B17_ready),
		.SB_T0_NORTH_SB_IN_B17_valid(Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B17_valid),
		.SB_T0_NORTH_SB_IN_B1_ready(Tile_X03_Y03_SB_T0_NORTH_SB_IN_B1_ready),
		.SB_T0_NORTH_SB_IN_B1_valid(Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B1_valid),
		.SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_OUT_B17(Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_OUT_B17_ready(Tile_X03_Y02_SB_T0_SOUTH_SB_IN_B17_ready),
		.SB_T0_NORTH_SB_OUT_B17_valid(Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B17_valid),
		.SB_T0_NORTH_SB_OUT_B1_ready(Tile_X03_Y02_SB_T0_SOUTH_SB_IN_B1_ready),
		.SB_T0_NORTH_SB_OUT_B1_valid(Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B1_valid),
		.SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_IN_B17(Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_IN_B17_ready(Tile_X03_Y03_SB_T0_SOUTH_SB_IN_B17_ready),
		.SB_T0_SOUTH_SB_IN_B17_valid(Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B17_valid),
		.SB_T0_SOUTH_SB_IN_B1_ready(Tile_X03_Y03_SB_T0_SOUTH_SB_IN_B1_ready),
		.SB_T0_SOUTH_SB_IN_B1_valid(Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B1_valid),
		.SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_OUT_B17(Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_OUT_B17_ready(Tile_X03_Y04_SB_T0_NORTH_SB_IN_B17_ready),
		.SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B17_valid),
		.SB_T0_SOUTH_SB_OUT_B1_ready(Tile_X03_Y04_SB_T0_NORTH_SB_IN_B1_ready),
		.SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B1_valid),
		.SB_T0_WEST_SB_IN_B1(Tile_X02_Y03_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_WEST_SB_IN_B17(Tile_X02_Y03_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_WEST_SB_IN_B17_ready(Tile_X03_Y03_SB_T0_WEST_SB_IN_B17_ready),
		.SB_T0_WEST_SB_IN_B17_valid(Tile_X02_Y03_SB_T0_EAST_SB_OUT_B17_valid),
		.SB_T0_WEST_SB_IN_B1_ready(Tile_X03_Y03_SB_T0_WEST_SB_IN_B1_ready),
		.SB_T0_WEST_SB_IN_B1_valid(Tile_X02_Y03_SB_T0_EAST_SB_OUT_B1_valid),
		.SB_T0_WEST_SB_OUT_B1(Tile_X03_Y03_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_WEST_SB_OUT_B17(Tile_X03_Y03_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_WEST_SB_OUT_B17_ready(Tile_X02_Y03_SB_T0_EAST_SB_IN_B17_ready),
		.SB_T0_WEST_SB_OUT_B17_valid(Tile_X03_Y03_SB_T0_WEST_SB_OUT_B17_valid),
		.SB_T0_WEST_SB_OUT_B1_ready(Tile_X02_Y03_SB_T0_EAST_SB_IN_B1_ready),
		.SB_T0_WEST_SB_OUT_B1_valid(Tile_X03_Y03_SB_T0_WEST_SB_OUT_B1_valid),
		.SB_T1_EAST_SB_IN_B1(const_0_1_out),
		.SB_T1_EAST_SB_IN_B17(const_0_17_out),
		.SB_T1_EAST_SB_IN_B17_ready(Tile_X03_Y03_SB_T1_EAST_SB_IN_B17_ready),
		.SB_T1_EAST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T1_EAST_SB_IN_B1_ready(Tile_X03_Y03_SB_T1_EAST_SB_IN_B1_ready),
		.SB_T1_EAST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T1_EAST_SB_OUT_B1(Tile_X03_Y03_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_EAST_SB_OUT_B17(Tile_X03_Y03_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T1_EAST_SB_OUT_B17_valid(Tile_X03_Y03_SB_T1_EAST_SB_OUT_B17_valid),
		.SB_T1_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T1_EAST_SB_OUT_B1_valid(Tile_X03_Y03_SB_T1_EAST_SB_OUT_B1_valid),
		.SB_T1_NORTH_SB_IN_B1(Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_IN_B17(Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_IN_B17_ready(Tile_X03_Y03_SB_T1_NORTH_SB_IN_B17_ready),
		.SB_T1_NORTH_SB_IN_B17_valid(Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B17_valid),
		.SB_T1_NORTH_SB_IN_B1_ready(Tile_X03_Y03_SB_T1_NORTH_SB_IN_B1_ready),
		.SB_T1_NORTH_SB_IN_B1_valid(Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B1_valid),
		.SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_OUT_B17(Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_OUT_B17_ready(Tile_X03_Y02_SB_T1_SOUTH_SB_IN_B17_ready),
		.SB_T1_NORTH_SB_OUT_B17_valid(Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B17_valid),
		.SB_T1_NORTH_SB_OUT_B1_ready(Tile_X03_Y02_SB_T1_SOUTH_SB_IN_B1_ready),
		.SB_T1_NORTH_SB_OUT_B1_valid(Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B1_valid),
		.SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_IN_B17(Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_IN_B17_ready(Tile_X03_Y03_SB_T1_SOUTH_SB_IN_B17_ready),
		.SB_T1_SOUTH_SB_IN_B17_valid(Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B17_valid),
		.SB_T1_SOUTH_SB_IN_B1_ready(Tile_X03_Y03_SB_T1_SOUTH_SB_IN_B1_ready),
		.SB_T1_SOUTH_SB_IN_B1_valid(Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B1_valid),
		.SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_OUT_B17(Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_OUT_B17_ready(Tile_X03_Y04_SB_T1_NORTH_SB_IN_B17_ready),
		.SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B17_valid),
		.SB_T1_SOUTH_SB_OUT_B1_ready(Tile_X03_Y04_SB_T1_NORTH_SB_IN_B1_ready),
		.SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B1_valid),
		.SB_T1_WEST_SB_IN_B1(Tile_X02_Y03_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_WEST_SB_IN_B17(Tile_X02_Y03_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_WEST_SB_IN_B17_ready(Tile_X03_Y03_SB_T1_WEST_SB_IN_B17_ready),
		.SB_T1_WEST_SB_IN_B17_valid(Tile_X02_Y03_SB_T1_EAST_SB_OUT_B17_valid),
		.SB_T1_WEST_SB_IN_B1_ready(Tile_X03_Y03_SB_T1_WEST_SB_IN_B1_ready),
		.SB_T1_WEST_SB_IN_B1_valid(Tile_X02_Y03_SB_T1_EAST_SB_OUT_B1_valid),
		.SB_T1_WEST_SB_OUT_B1(Tile_X03_Y03_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_WEST_SB_OUT_B17(Tile_X03_Y03_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_WEST_SB_OUT_B17_ready(Tile_X02_Y03_SB_T1_EAST_SB_IN_B17_ready),
		.SB_T1_WEST_SB_OUT_B17_valid(Tile_X03_Y03_SB_T1_WEST_SB_OUT_B17_valid),
		.SB_T1_WEST_SB_OUT_B1_ready(Tile_X02_Y03_SB_T1_EAST_SB_IN_B1_ready),
		.SB_T1_WEST_SB_OUT_B1_valid(Tile_X03_Y03_SB_T1_WEST_SB_OUT_B1_valid),
		.SB_T2_EAST_SB_IN_B1(const_0_1_out),
		.SB_T2_EAST_SB_IN_B17(const_0_17_out),
		.SB_T2_EAST_SB_IN_B17_ready(Tile_X03_Y03_SB_T2_EAST_SB_IN_B17_ready),
		.SB_T2_EAST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T2_EAST_SB_IN_B1_ready(Tile_X03_Y03_SB_T2_EAST_SB_IN_B1_ready),
		.SB_T2_EAST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T2_EAST_SB_OUT_B1(Tile_X03_Y03_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_EAST_SB_OUT_B17(Tile_X03_Y03_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T2_EAST_SB_OUT_B17_valid(Tile_X03_Y03_SB_T2_EAST_SB_OUT_B17_valid),
		.SB_T2_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T2_EAST_SB_OUT_B1_valid(Tile_X03_Y03_SB_T2_EAST_SB_OUT_B1_valid),
		.SB_T2_NORTH_SB_IN_B1(Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_IN_B17(Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_IN_B17_ready(Tile_X03_Y03_SB_T2_NORTH_SB_IN_B17_ready),
		.SB_T2_NORTH_SB_IN_B17_valid(Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B17_valid),
		.SB_T2_NORTH_SB_IN_B1_ready(Tile_X03_Y03_SB_T2_NORTH_SB_IN_B1_ready),
		.SB_T2_NORTH_SB_IN_B1_valid(Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B1_valid),
		.SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_OUT_B17(Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_OUT_B17_ready(Tile_X03_Y02_SB_T2_SOUTH_SB_IN_B17_ready),
		.SB_T2_NORTH_SB_OUT_B17_valid(Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B17_valid),
		.SB_T2_NORTH_SB_OUT_B1_ready(Tile_X03_Y02_SB_T2_SOUTH_SB_IN_B1_ready),
		.SB_T2_NORTH_SB_OUT_B1_valid(Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B1_valid),
		.SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_IN_B17(Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_IN_B17_ready(Tile_X03_Y03_SB_T2_SOUTH_SB_IN_B17_ready),
		.SB_T2_SOUTH_SB_IN_B17_valid(Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B17_valid),
		.SB_T2_SOUTH_SB_IN_B1_ready(Tile_X03_Y03_SB_T2_SOUTH_SB_IN_B1_ready),
		.SB_T2_SOUTH_SB_IN_B1_valid(Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B1_valid),
		.SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_OUT_B17(Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_OUT_B17_ready(Tile_X03_Y04_SB_T2_NORTH_SB_IN_B17_ready),
		.SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B17_valid),
		.SB_T2_SOUTH_SB_OUT_B1_ready(Tile_X03_Y04_SB_T2_NORTH_SB_IN_B1_ready),
		.SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B1_valid),
		.SB_T2_WEST_SB_IN_B1(Tile_X02_Y03_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_WEST_SB_IN_B17(Tile_X02_Y03_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_WEST_SB_IN_B17_ready(Tile_X03_Y03_SB_T2_WEST_SB_IN_B17_ready),
		.SB_T2_WEST_SB_IN_B17_valid(Tile_X02_Y03_SB_T2_EAST_SB_OUT_B17_valid),
		.SB_T2_WEST_SB_IN_B1_ready(Tile_X03_Y03_SB_T2_WEST_SB_IN_B1_ready),
		.SB_T2_WEST_SB_IN_B1_valid(Tile_X02_Y03_SB_T2_EAST_SB_OUT_B1_valid),
		.SB_T2_WEST_SB_OUT_B1(Tile_X03_Y03_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_WEST_SB_OUT_B17(Tile_X03_Y03_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_WEST_SB_OUT_B17_ready(Tile_X02_Y03_SB_T2_EAST_SB_IN_B17_ready),
		.SB_T2_WEST_SB_OUT_B17_valid(Tile_X03_Y03_SB_T2_WEST_SB_OUT_B17_valid),
		.SB_T2_WEST_SB_OUT_B1_ready(Tile_X02_Y03_SB_T2_EAST_SB_IN_B1_ready),
		.SB_T2_WEST_SB_OUT_B1_valid(Tile_X03_Y03_SB_T2_WEST_SB_OUT_B1_valid),
		.SB_T3_EAST_SB_IN_B1(const_0_1_out),
		.SB_T3_EAST_SB_IN_B17(const_0_17_out),
		.SB_T3_EAST_SB_IN_B17_ready(Tile_X03_Y03_SB_T3_EAST_SB_IN_B17_ready),
		.SB_T3_EAST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T3_EAST_SB_IN_B1_ready(Tile_X03_Y03_SB_T3_EAST_SB_IN_B1_ready),
		.SB_T3_EAST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T3_EAST_SB_OUT_B1(Tile_X03_Y03_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_EAST_SB_OUT_B17(Tile_X03_Y03_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T3_EAST_SB_OUT_B17_valid(Tile_X03_Y03_SB_T3_EAST_SB_OUT_B17_valid),
		.SB_T3_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T3_EAST_SB_OUT_B1_valid(Tile_X03_Y03_SB_T3_EAST_SB_OUT_B1_valid),
		.SB_T3_NORTH_SB_IN_B1(Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_IN_B17(Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_IN_B17_ready(Tile_X03_Y03_SB_T3_NORTH_SB_IN_B17_ready),
		.SB_T3_NORTH_SB_IN_B17_valid(Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B17_valid),
		.SB_T3_NORTH_SB_IN_B1_ready(Tile_X03_Y03_SB_T3_NORTH_SB_IN_B1_ready),
		.SB_T3_NORTH_SB_IN_B1_valid(Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B1_valid),
		.SB_T3_NORTH_SB_OUT_B1(Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_OUT_B17(Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_OUT_B17_ready(Tile_X03_Y02_SB_T3_SOUTH_SB_IN_B17_ready),
		.SB_T3_NORTH_SB_OUT_B17_valid(Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B17_valid),
		.SB_T3_NORTH_SB_OUT_B1_ready(Tile_X03_Y02_SB_T3_SOUTH_SB_IN_B1_ready),
		.SB_T3_NORTH_SB_OUT_B1_valid(Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B1_valid),
		.SB_T3_SOUTH_SB_IN_B1(Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_IN_B17(Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_IN_B17_ready(Tile_X03_Y03_SB_T3_SOUTH_SB_IN_B17_ready),
		.SB_T3_SOUTH_SB_IN_B17_valid(Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B17_valid),
		.SB_T3_SOUTH_SB_IN_B1_ready(Tile_X03_Y03_SB_T3_SOUTH_SB_IN_B1_ready),
		.SB_T3_SOUTH_SB_IN_B1_valid(Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B1_valid),
		.SB_T3_SOUTH_SB_OUT_B1(Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_OUT_B17(Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_OUT_B17_ready(Tile_X03_Y04_SB_T3_NORTH_SB_IN_B17_ready),
		.SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B17_valid),
		.SB_T3_SOUTH_SB_OUT_B1_ready(Tile_X03_Y04_SB_T3_NORTH_SB_IN_B1_ready),
		.SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B1_valid),
		.SB_T3_WEST_SB_IN_B1(Tile_X02_Y03_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_WEST_SB_IN_B17(Tile_X02_Y03_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_WEST_SB_IN_B17_ready(Tile_X03_Y03_SB_T3_WEST_SB_IN_B17_ready),
		.SB_T3_WEST_SB_IN_B17_valid(Tile_X02_Y03_SB_T3_EAST_SB_OUT_B17_valid),
		.SB_T3_WEST_SB_IN_B1_ready(Tile_X03_Y03_SB_T3_WEST_SB_IN_B1_ready),
		.SB_T3_WEST_SB_IN_B1_valid(Tile_X02_Y03_SB_T3_EAST_SB_OUT_B1_valid),
		.SB_T3_WEST_SB_OUT_B1(Tile_X03_Y03_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_WEST_SB_OUT_B17(Tile_X03_Y03_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_WEST_SB_OUT_B17_ready(Tile_X02_Y03_SB_T3_EAST_SB_IN_B17_ready),
		.SB_T3_WEST_SB_OUT_B17_valid(Tile_X03_Y03_SB_T3_WEST_SB_OUT_B17_valid),
		.SB_T3_WEST_SB_OUT_B1_ready(Tile_X02_Y03_SB_T3_EAST_SB_IN_B1_ready),
		.SB_T3_WEST_SB_OUT_B1_valid(Tile_X03_Y03_SB_T3_WEST_SB_OUT_B1_valid),
		.SB_T4_EAST_SB_IN_B1(const_0_1_out),
		.SB_T4_EAST_SB_IN_B17(const_0_17_out),
		.SB_T4_EAST_SB_IN_B17_ready(Tile_X03_Y03_SB_T4_EAST_SB_IN_B17_ready),
		.SB_T4_EAST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T4_EAST_SB_IN_B1_ready(Tile_X03_Y03_SB_T4_EAST_SB_IN_B1_ready),
		.SB_T4_EAST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T4_EAST_SB_OUT_B1(Tile_X03_Y03_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_EAST_SB_OUT_B17(Tile_X03_Y03_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T4_EAST_SB_OUT_B17_valid(Tile_X03_Y03_SB_T4_EAST_SB_OUT_B17_valid),
		.SB_T4_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T4_EAST_SB_OUT_B1_valid(Tile_X03_Y03_SB_T4_EAST_SB_OUT_B1_valid),
		.SB_T4_NORTH_SB_IN_B1(Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_IN_B17(Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_IN_B17_ready(Tile_X03_Y03_SB_T4_NORTH_SB_IN_B17_ready),
		.SB_T4_NORTH_SB_IN_B17_valid(Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B17_valid),
		.SB_T4_NORTH_SB_IN_B1_ready(Tile_X03_Y03_SB_T4_NORTH_SB_IN_B1_ready),
		.SB_T4_NORTH_SB_IN_B1_valid(Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B1_valid),
		.SB_T4_NORTH_SB_OUT_B1(Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_OUT_B17(Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_OUT_B17_ready(Tile_X03_Y02_SB_T4_SOUTH_SB_IN_B17_ready),
		.SB_T4_NORTH_SB_OUT_B17_valid(Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B17_valid),
		.SB_T4_NORTH_SB_OUT_B1_ready(Tile_X03_Y02_SB_T4_SOUTH_SB_IN_B1_ready),
		.SB_T4_NORTH_SB_OUT_B1_valid(Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B1_valid),
		.SB_T4_SOUTH_SB_IN_B1(Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_IN_B17(Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_IN_B17_ready(Tile_X03_Y03_SB_T4_SOUTH_SB_IN_B17_ready),
		.SB_T4_SOUTH_SB_IN_B17_valid(Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B17_valid),
		.SB_T4_SOUTH_SB_IN_B1_ready(Tile_X03_Y03_SB_T4_SOUTH_SB_IN_B1_ready),
		.SB_T4_SOUTH_SB_IN_B1_valid(Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B1_valid),
		.SB_T4_SOUTH_SB_OUT_B1(Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_OUT_B17(Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_OUT_B17_ready(Tile_X03_Y04_SB_T4_NORTH_SB_IN_B17_ready),
		.SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B17_valid),
		.SB_T4_SOUTH_SB_OUT_B1_ready(Tile_X03_Y04_SB_T4_NORTH_SB_IN_B1_ready),
		.SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B1_valid),
		.SB_T4_WEST_SB_IN_B1(Tile_X02_Y03_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_WEST_SB_IN_B17(Tile_X02_Y03_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_WEST_SB_IN_B17_ready(Tile_X03_Y03_SB_T4_WEST_SB_IN_B17_ready),
		.SB_T4_WEST_SB_IN_B17_valid(Tile_X02_Y03_SB_T4_EAST_SB_OUT_B17_valid),
		.SB_T4_WEST_SB_IN_B1_ready(Tile_X03_Y03_SB_T4_WEST_SB_IN_B1_ready),
		.SB_T4_WEST_SB_IN_B1_valid(Tile_X02_Y03_SB_T4_EAST_SB_OUT_B1_valid),
		.SB_T4_WEST_SB_OUT_B1(Tile_X03_Y03_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_WEST_SB_OUT_B17(Tile_X03_Y03_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_WEST_SB_OUT_B17_ready(Tile_X02_Y03_SB_T4_EAST_SB_IN_B17_ready),
		.SB_T4_WEST_SB_OUT_B17_valid(Tile_X03_Y03_SB_T4_WEST_SB_OUT_B17_valid),
		.SB_T4_WEST_SB_OUT_B1_ready(Tile_X02_Y03_SB_T4_EAST_SB_IN_B1_ready),
		.SB_T4_WEST_SB_OUT_B1_valid(Tile_X03_Y03_SB_T4_WEST_SB_OUT_B1_valid),
		.clk(Tile_X02_Y03_clk_pass_through_out_right),
		.clk_out(Tile_X03_Y03_clk_out),
		.config_config_addr(Tile_X03_Y02_config_out_config_addr),
		.config_config_data(Tile_X03_Y02_config_out_config_data),
		.config_out_config_addr(Tile_X03_Y03_config_out_config_addr),
		.config_out_config_data(Tile_X03_Y03_config_out_config_data),
		.config_out_read(Tile_X03_Y03_config_out_read),
		.config_out_write(Tile_X03_Y03_config_out_write),
		.config_read(Tile_X03_Y02_config_out_read),
		.config_write(Tile_X03_Y02_config_out_write),
		.flush(Tile_X03_Y02_flush_out),
		.flush_out(Tile_X03_Y03_flush_out),
		.hi(Tile_X03_Y03_hi),
		.lo(Tile_X03_Y03_lo),
		.read_config_data(Tile_X03_Y03_read_config_data),
		.read_config_data_in(Tile_X03_Y02_read_config_data),
		.reset(Tile_X03_Y02_reset_out),
		.reset_out(Tile_X03_Y03_reset_out),
		.stall(Tile_X03_Y02_stall_out),
		.stall_out(Tile_X03_Y03_stall_out),
		.tile_id(Tile_X03_Y03_tile_id)
	);
	wire [15:0] Tile_X03_Y04_tile_id;
	assign Tile_X03_Y04_tile_id = {Tile_X03_Y04_lo[7], Tile_X03_Y04_lo[7], Tile_X03_Y04_lo[6], Tile_X03_Y04_lo[6], Tile_X03_Y04_lo[5], Tile_X03_Y04_lo[5], Tile_X03_Y04_hi[5], Tile_X03_Y04_hi[4], Tile_X03_Y04_lo[3], Tile_X03_Y04_lo[3], Tile_X03_Y04_lo[2], Tile_X03_Y04_lo[2], Tile_X03_Y04_lo[1], Tile_X03_Y04_hi[1], Tile_X03_Y04_lo[0], Tile_X03_Y04_lo[0]};
	Tile_MemCore Tile_X03_Y04(
		.SB_T0_EAST_SB_IN_B1(const_0_1_out),
		.SB_T0_EAST_SB_IN_B17(const_0_17_out),
		.SB_T0_EAST_SB_IN_B17_ready(Tile_X03_Y04_SB_T0_EAST_SB_IN_B17_ready),
		.SB_T0_EAST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T0_EAST_SB_IN_B1_ready(Tile_X03_Y04_SB_T0_EAST_SB_IN_B1_ready),
		.SB_T0_EAST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T0_EAST_SB_OUT_B1(Tile_X03_Y04_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_EAST_SB_OUT_B17(Tile_X03_Y04_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T0_EAST_SB_OUT_B17_valid(Tile_X03_Y04_SB_T0_EAST_SB_OUT_B17_valid),
		.SB_T0_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T0_EAST_SB_OUT_B1_valid(Tile_X03_Y04_SB_T0_EAST_SB_OUT_B1_valid),
		.SB_T0_NORTH_SB_IN_B1(Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_IN_B17(Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_IN_B17_ready(Tile_X03_Y04_SB_T0_NORTH_SB_IN_B17_ready),
		.SB_T0_NORTH_SB_IN_B17_valid(Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B17_valid),
		.SB_T0_NORTH_SB_IN_B1_ready(Tile_X03_Y04_SB_T0_NORTH_SB_IN_B1_ready),
		.SB_T0_NORTH_SB_IN_B1_valid(Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B1_valid),
		.SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_OUT_B17(Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B17),
		.SB_T0_NORTH_SB_OUT_B17_ready(Tile_X03_Y03_SB_T0_SOUTH_SB_IN_B17_ready),
		.SB_T0_NORTH_SB_OUT_B17_valid(Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B17_valid),
		.SB_T0_NORTH_SB_OUT_B1_ready(Tile_X03_Y03_SB_T0_SOUTH_SB_IN_B1_ready),
		.SB_T0_NORTH_SB_OUT_B1_valid(Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B1_valid),
		.SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
		.SB_T0_SOUTH_SB_IN_B17(const_0_17_out),
		.SB_T0_SOUTH_SB_IN_B17_ready(Tile_X03_Y04_SB_T0_SOUTH_SB_IN_B17_ready),
		.SB_T0_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T0_SOUTH_SB_IN_B1_ready(Tile_X03_Y04_SB_T0_SOUTH_SB_IN_B1_ready),
		.SB_T0_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_OUT_B17(Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B17),
		.SB_T0_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B17_valid),
		.SB_T0_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B1_valid),
		.SB_T0_WEST_SB_IN_B1(Tile_X02_Y04_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_WEST_SB_IN_B17(Tile_X02_Y04_SB_T0_EAST_SB_OUT_B17),
		.SB_T0_WEST_SB_IN_B17_ready(Tile_X03_Y04_SB_T0_WEST_SB_IN_B17_ready),
		.SB_T0_WEST_SB_IN_B17_valid(Tile_X02_Y04_SB_T0_EAST_SB_OUT_B17_valid),
		.SB_T0_WEST_SB_IN_B1_ready(Tile_X03_Y04_SB_T0_WEST_SB_IN_B1_ready),
		.SB_T0_WEST_SB_IN_B1_valid(Tile_X02_Y04_SB_T0_EAST_SB_OUT_B1_valid),
		.SB_T0_WEST_SB_OUT_B1(Tile_X03_Y04_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_WEST_SB_OUT_B17(Tile_X03_Y04_SB_T0_WEST_SB_OUT_B17),
		.SB_T0_WEST_SB_OUT_B17_ready(Tile_X02_Y04_SB_T0_EAST_SB_IN_B17_ready),
		.SB_T0_WEST_SB_OUT_B17_valid(Tile_X03_Y04_SB_T0_WEST_SB_OUT_B17_valid),
		.SB_T0_WEST_SB_OUT_B1_ready(Tile_X02_Y04_SB_T0_EAST_SB_IN_B1_ready),
		.SB_T0_WEST_SB_OUT_B1_valid(Tile_X03_Y04_SB_T0_WEST_SB_OUT_B1_valid),
		.SB_T1_EAST_SB_IN_B1(const_0_1_out),
		.SB_T1_EAST_SB_IN_B17(const_0_17_out),
		.SB_T1_EAST_SB_IN_B17_ready(Tile_X03_Y04_SB_T1_EAST_SB_IN_B17_ready),
		.SB_T1_EAST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T1_EAST_SB_IN_B1_ready(Tile_X03_Y04_SB_T1_EAST_SB_IN_B1_ready),
		.SB_T1_EAST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T1_EAST_SB_OUT_B1(Tile_X03_Y04_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_EAST_SB_OUT_B17(Tile_X03_Y04_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T1_EAST_SB_OUT_B17_valid(Tile_X03_Y04_SB_T1_EAST_SB_OUT_B17_valid),
		.SB_T1_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T1_EAST_SB_OUT_B1_valid(Tile_X03_Y04_SB_T1_EAST_SB_OUT_B1_valid),
		.SB_T1_NORTH_SB_IN_B1(Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_IN_B17(Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_IN_B17_ready(Tile_X03_Y04_SB_T1_NORTH_SB_IN_B17_ready),
		.SB_T1_NORTH_SB_IN_B17_valid(Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B17_valid),
		.SB_T1_NORTH_SB_IN_B1_ready(Tile_X03_Y04_SB_T1_NORTH_SB_IN_B1_ready),
		.SB_T1_NORTH_SB_IN_B1_valid(Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B1_valid),
		.SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_OUT_B17(Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B17),
		.SB_T1_NORTH_SB_OUT_B17_ready(Tile_X03_Y03_SB_T1_SOUTH_SB_IN_B17_ready),
		.SB_T1_NORTH_SB_OUT_B17_valid(Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B17_valid),
		.SB_T1_NORTH_SB_OUT_B1_ready(Tile_X03_Y03_SB_T1_SOUTH_SB_IN_B1_ready),
		.SB_T1_NORTH_SB_OUT_B1_valid(Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B1_valid),
		.SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
		.SB_T1_SOUTH_SB_IN_B17(const_0_17_out),
		.SB_T1_SOUTH_SB_IN_B17_ready(Tile_X03_Y04_SB_T1_SOUTH_SB_IN_B17_ready),
		.SB_T1_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T1_SOUTH_SB_IN_B1_ready(Tile_X03_Y04_SB_T1_SOUTH_SB_IN_B1_ready),
		.SB_T1_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_OUT_B17(Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B17),
		.SB_T1_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B17_valid),
		.SB_T1_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B1_valid),
		.SB_T1_WEST_SB_IN_B1(Tile_X02_Y04_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_WEST_SB_IN_B17(Tile_X02_Y04_SB_T1_EAST_SB_OUT_B17),
		.SB_T1_WEST_SB_IN_B17_ready(Tile_X03_Y04_SB_T1_WEST_SB_IN_B17_ready),
		.SB_T1_WEST_SB_IN_B17_valid(Tile_X02_Y04_SB_T1_EAST_SB_OUT_B17_valid),
		.SB_T1_WEST_SB_IN_B1_ready(Tile_X03_Y04_SB_T1_WEST_SB_IN_B1_ready),
		.SB_T1_WEST_SB_IN_B1_valid(Tile_X02_Y04_SB_T1_EAST_SB_OUT_B1_valid),
		.SB_T1_WEST_SB_OUT_B1(Tile_X03_Y04_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_WEST_SB_OUT_B17(Tile_X03_Y04_SB_T1_WEST_SB_OUT_B17),
		.SB_T1_WEST_SB_OUT_B17_ready(Tile_X02_Y04_SB_T1_EAST_SB_IN_B17_ready),
		.SB_T1_WEST_SB_OUT_B17_valid(Tile_X03_Y04_SB_T1_WEST_SB_OUT_B17_valid),
		.SB_T1_WEST_SB_OUT_B1_ready(Tile_X02_Y04_SB_T1_EAST_SB_IN_B1_ready),
		.SB_T1_WEST_SB_OUT_B1_valid(Tile_X03_Y04_SB_T1_WEST_SB_OUT_B1_valid),
		.SB_T2_EAST_SB_IN_B1(const_0_1_out),
		.SB_T2_EAST_SB_IN_B17(const_0_17_out),
		.SB_T2_EAST_SB_IN_B17_ready(Tile_X03_Y04_SB_T2_EAST_SB_IN_B17_ready),
		.SB_T2_EAST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T2_EAST_SB_IN_B1_ready(Tile_X03_Y04_SB_T2_EAST_SB_IN_B1_ready),
		.SB_T2_EAST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T2_EAST_SB_OUT_B1(Tile_X03_Y04_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_EAST_SB_OUT_B17(Tile_X03_Y04_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T2_EAST_SB_OUT_B17_valid(Tile_X03_Y04_SB_T2_EAST_SB_OUT_B17_valid),
		.SB_T2_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T2_EAST_SB_OUT_B1_valid(Tile_X03_Y04_SB_T2_EAST_SB_OUT_B1_valid),
		.SB_T2_NORTH_SB_IN_B1(Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_IN_B17(Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_IN_B17_ready(Tile_X03_Y04_SB_T2_NORTH_SB_IN_B17_ready),
		.SB_T2_NORTH_SB_IN_B17_valid(Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B17_valid),
		.SB_T2_NORTH_SB_IN_B1_ready(Tile_X03_Y04_SB_T2_NORTH_SB_IN_B1_ready),
		.SB_T2_NORTH_SB_IN_B1_valid(Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B1_valid),
		.SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_OUT_B17(Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B17),
		.SB_T2_NORTH_SB_OUT_B17_ready(Tile_X03_Y03_SB_T2_SOUTH_SB_IN_B17_ready),
		.SB_T2_NORTH_SB_OUT_B17_valid(Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B17_valid),
		.SB_T2_NORTH_SB_OUT_B1_ready(Tile_X03_Y03_SB_T2_SOUTH_SB_IN_B1_ready),
		.SB_T2_NORTH_SB_OUT_B1_valid(Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B1_valid),
		.SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
		.SB_T2_SOUTH_SB_IN_B17(const_0_17_out),
		.SB_T2_SOUTH_SB_IN_B17_ready(Tile_X03_Y04_SB_T2_SOUTH_SB_IN_B17_ready),
		.SB_T2_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T2_SOUTH_SB_IN_B1_ready(Tile_X03_Y04_SB_T2_SOUTH_SB_IN_B1_ready),
		.SB_T2_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_OUT_B17(Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B17),
		.SB_T2_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B17_valid),
		.SB_T2_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B1_valid),
		.SB_T2_WEST_SB_IN_B1(Tile_X02_Y04_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_WEST_SB_IN_B17(Tile_X02_Y04_SB_T2_EAST_SB_OUT_B17),
		.SB_T2_WEST_SB_IN_B17_ready(Tile_X03_Y04_SB_T2_WEST_SB_IN_B17_ready),
		.SB_T2_WEST_SB_IN_B17_valid(Tile_X02_Y04_SB_T2_EAST_SB_OUT_B17_valid),
		.SB_T2_WEST_SB_IN_B1_ready(Tile_X03_Y04_SB_T2_WEST_SB_IN_B1_ready),
		.SB_T2_WEST_SB_IN_B1_valid(Tile_X02_Y04_SB_T2_EAST_SB_OUT_B1_valid),
		.SB_T2_WEST_SB_OUT_B1(Tile_X03_Y04_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_WEST_SB_OUT_B17(Tile_X03_Y04_SB_T2_WEST_SB_OUT_B17),
		.SB_T2_WEST_SB_OUT_B17_ready(Tile_X02_Y04_SB_T2_EAST_SB_IN_B17_ready),
		.SB_T2_WEST_SB_OUT_B17_valid(Tile_X03_Y04_SB_T2_WEST_SB_OUT_B17_valid),
		.SB_T2_WEST_SB_OUT_B1_ready(Tile_X02_Y04_SB_T2_EAST_SB_IN_B1_ready),
		.SB_T2_WEST_SB_OUT_B1_valid(Tile_X03_Y04_SB_T2_WEST_SB_OUT_B1_valid),
		.SB_T3_EAST_SB_IN_B1(const_0_1_out),
		.SB_T3_EAST_SB_IN_B17(const_0_17_out),
		.SB_T3_EAST_SB_IN_B17_ready(Tile_X03_Y04_SB_T3_EAST_SB_IN_B17_ready),
		.SB_T3_EAST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T3_EAST_SB_IN_B1_ready(Tile_X03_Y04_SB_T3_EAST_SB_IN_B1_ready),
		.SB_T3_EAST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T3_EAST_SB_OUT_B1(Tile_X03_Y04_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_EAST_SB_OUT_B17(Tile_X03_Y04_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T3_EAST_SB_OUT_B17_valid(Tile_X03_Y04_SB_T3_EAST_SB_OUT_B17_valid),
		.SB_T3_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T3_EAST_SB_OUT_B1_valid(Tile_X03_Y04_SB_T3_EAST_SB_OUT_B1_valid),
		.SB_T3_NORTH_SB_IN_B1(Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_IN_B17(Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_IN_B17_ready(Tile_X03_Y04_SB_T3_NORTH_SB_IN_B17_ready),
		.SB_T3_NORTH_SB_IN_B17_valid(Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B17_valid),
		.SB_T3_NORTH_SB_IN_B1_ready(Tile_X03_Y04_SB_T3_NORTH_SB_IN_B1_ready),
		.SB_T3_NORTH_SB_IN_B1_valid(Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B1_valid),
		.SB_T3_NORTH_SB_OUT_B1(Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B1),
		.SB_T3_NORTH_SB_OUT_B17(Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B17),
		.SB_T3_NORTH_SB_OUT_B17_ready(Tile_X03_Y03_SB_T3_SOUTH_SB_IN_B17_ready),
		.SB_T3_NORTH_SB_OUT_B17_valid(Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B17_valid),
		.SB_T3_NORTH_SB_OUT_B1_ready(Tile_X03_Y03_SB_T3_SOUTH_SB_IN_B1_ready),
		.SB_T3_NORTH_SB_OUT_B1_valid(Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B1_valid),
		.SB_T3_SOUTH_SB_IN_B1(const_0_1_out),
		.SB_T3_SOUTH_SB_IN_B17(const_0_17_out),
		.SB_T3_SOUTH_SB_IN_B17_ready(Tile_X03_Y04_SB_T3_SOUTH_SB_IN_B17_ready),
		.SB_T3_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T3_SOUTH_SB_IN_B1_ready(Tile_X03_Y04_SB_T3_SOUTH_SB_IN_B1_ready),
		.SB_T3_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T3_SOUTH_SB_OUT_B1(Tile_X03_Y04_SB_T3_SOUTH_SB_OUT_B1),
		.SB_T3_SOUTH_SB_OUT_B17(Tile_X03_Y04_SB_T3_SOUTH_SB_OUT_B17),
		.SB_T3_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X03_Y04_SB_T3_SOUTH_SB_OUT_B17_valid),
		.SB_T3_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X03_Y04_SB_T3_SOUTH_SB_OUT_B1_valid),
		.SB_T3_WEST_SB_IN_B1(Tile_X02_Y04_SB_T3_EAST_SB_OUT_B1),
		.SB_T3_WEST_SB_IN_B17(Tile_X02_Y04_SB_T3_EAST_SB_OUT_B17),
		.SB_T3_WEST_SB_IN_B17_ready(Tile_X03_Y04_SB_T3_WEST_SB_IN_B17_ready),
		.SB_T3_WEST_SB_IN_B17_valid(Tile_X02_Y04_SB_T3_EAST_SB_OUT_B17_valid),
		.SB_T3_WEST_SB_IN_B1_ready(Tile_X03_Y04_SB_T3_WEST_SB_IN_B1_ready),
		.SB_T3_WEST_SB_IN_B1_valid(Tile_X02_Y04_SB_T3_EAST_SB_OUT_B1_valid),
		.SB_T3_WEST_SB_OUT_B1(Tile_X03_Y04_SB_T3_WEST_SB_OUT_B1),
		.SB_T3_WEST_SB_OUT_B17(Tile_X03_Y04_SB_T3_WEST_SB_OUT_B17),
		.SB_T3_WEST_SB_OUT_B17_ready(Tile_X02_Y04_SB_T3_EAST_SB_IN_B17_ready),
		.SB_T3_WEST_SB_OUT_B17_valid(Tile_X03_Y04_SB_T3_WEST_SB_OUT_B17_valid),
		.SB_T3_WEST_SB_OUT_B1_ready(Tile_X02_Y04_SB_T3_EAST_SB_IN_B1_ready),
		.SB_T3_WEST_SB_OUT_B1_valid(Tile_X03_Y04_SB_T3_WEST_SB_OUT_B1_valid),
		.SB_T4_EAST_SB_IN_B1(const_0_1_out),
		.SB_T4_EAST_SB_IN_B17(const_0_17_out),
		.SB_T4_EAST_SB_IN_B17_ready(Tile_X03_Y04_SB_T4_EAST_SB_IN_B17_ready),
		.SB_T4_EAST_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T4_EAST_SB_IN_B1_ready(Tile_X03_Y04_SB_T4_EAST_SB_IN_B1_ready),
		.SB_T4_EAST_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T4_EAST_SB_OUT_B1(Tile_X03_Y04_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_EAST_SB_OUT_B17(Tile_X03_Y04_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T4_EAST_SB_OUT_B17_valid(Tile_X03_Y04_SB_T4_EAST_SB_OUT_B17_valid),
		.SB_T4_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T4_EAST_SB_OUT_B1_valid(Tile_X03_Y04_SB_T4_EAST_SB_OUT_B1_valid),
		.SB_T4_NORTH_SB_IN_B1(Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_IN_B17(Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_IN_B17_ready(Tile_X03_Y04_SB_T4_NORTH_SB_IN_B17_ready),
		.SB_T4_NORTH_SB_IN_B17_valid(Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B17_valid),
		.SB_T4_NORTH_SB_IN_B1_ready(Tile_X03_Y04_SB_T4_NORTH_SB_IN_B1_ready),
		.SB_T4_NORTH_SB_IN_B1_valid(Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B1_valid),
		.SB_T4_NORTH_SB_OUT_B1(Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B1),
		.SB_T4_NORTH_SB_OUT_B17(Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B17),
		.SB_T4_NORTH_SB_OUT_B17_ready(Tile_X03_Y03_SB_T4_SOUTH_SB_IN_B17_ready),
		.SB_T4_NORTH_SB_OUT_B17_valid(Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B17_valid),
		.SB_T4_NORTH_SB_OUT_B1_ready(Tile_X03_Y03_SB_T4_SOUTH_SB_IN_B1_ready),
		.SB_T4_NORTH_SB_OUT_B1_valid(Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B1_valid),
		.SB_T4_SOUTH_SB_IN_B1(const_0_1_out),
		.SB_T4_SOUTH_SB_IN_B17(const_0_17_out),
		.SB_T4_SOUTH_SB_IN_B17_ready(Tile_X03_Y04_SB_T4_SOUTH_SB_IN_B17_ready),
		.SB_T4_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
		.SB_T4_SOUTH_SB_IN_B1_ready(Tile_X03_Y04_SB_T4_SOUTH_SB_IN_B1_ready),
		.SB_T4_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
		.SB_T4_SOUTH_SB_OUT_B1(Tile_X03_Y04_SB_T4_SOUTH_SB_OUT_B1),
		.SB_T4_SOUTH_SB_OUT_B17(Tile_X03_Y04_SB_T4_SOUTH_SB_OUT_B17),
		.SB_T4_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
		.SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X03_Y04_SB_T4_SOUTH_SB_OUT_B17_valid),
		.SB_T4_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
		.SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X03_Y04_SB_T4_SOUTH_SB_OUT_B1_valid),
		.SB_T4_WEST_SB_IN_B1(Tile_X02_Y04_SB_T4_EAST_SB_OUT_B1),
		.SB_T4_WEST_SB_IN_B17(Tile_X02_Y04_SB_T4_EAST_SB_OUT_B17),
		.SB_T4_WEST_SB_IN_B17_ready(Tile_X03_Y04_SB_T4_WEST_SB_IN_B17_ready),
		.SB_T4_WEST_SB_IN_B17_valid(Tile_X02_Y04_SB_T4_EAST_SB_OUT_B17_valid),
		.SB_T4_WEST_SB_IN_B1_ready(Tile_X03_Y04_SB_T4_WEST_SB_IN_B1_ready),
		.SB_T4_WEST_SB_IN_B1_valid(Tile_X02_Y04_SB_T4_EAST_SB_OUT_B1_valid),
		.SB_T4_WEST_SB_OUT_B1(Tile_X03_Y04_SB_T4_WEST_SB_OUT_B1),
		.SB_T4_WEST_SB_OUT_B17(Tile_X03_Y04_SB_T4_WEST_SB_OUT_B17),
		.SB_T4_WEST_SB_OUT_B17_ready(Tile_X02_Y04_SB_T4_EAST_SB_IN_B17_ready),
		.SB_T4_WEST_SB_OUT_B17_valid(Tile_X03_Y04_SB_T4_WEST_SB_OUT_B17_valid),
		.SB_T4_WEST_SB_OUT_B1_ready(Tile_X02_Y04_SB_T4_EAST_SB_IN_B1_ready),
		.SB_T4_WEST_SB_OUT_B1_valid(Tile_X03_Y04_SB_T4_WEST_SB_OUT_B1_valid),
		.clk(Tile_X02_Y04_clk_pass_through_out_right),
		.clk_out(Tile_X03_Y04_clk_out),
		.config_config_addr(Tile_X03_Y03_config_out_config_addr),
		.config_config_data(Tile_X03_Y03_config_out_config_data),
		.config_out_config_addr(Tile_X03_Y04_config_out_config_addr),
		.config_out_config_data(Tile_X03_Y04_config_out_config_data),
		.config_out_read(Tile_X03_Y04_config_out_read),
		.config_out_write(Tile_X03_Y04_config_out_write),
		.config_read(Tile_X03_Y03_config_out_read),
		.config_write(Tile_X03_Y03_config_out_write),
		.flush(Tile_X03_Y03_flush_out),
		.flush_out(Tile_X03_Y04_flush_out),
		.hi(Tile_X03_Y04_hi),
		.lo(Tile_X03_Y04_lo),
		.read_config_data(Tile_X03_Y04_read_config_data),
		.read_config_data_in(Tile_X03_Y03_read_config_data),
		.reset(Tile_X03_Y03_reset_out),
		.reset_out(Tile_X03_Y04_reset_out),
		.stall(Tile_X03_Y03_stall_out),
		.stall_out(Tile_X03_Y04_stall_out),
		.tile_id(Tile_X03_Y04_tile_id)
	);
	corebit_const #(.value(1'b0)) bit_const_0_None(.out(bit_const_0_None_out));
	coreir_const #(
		.value(1'h0),
		.width(1)
	) const_0_1(.out(const_0_1_out));
	coreir_const #(
		.value(17'h00000),
		.width(17)
	) const_0_17(.out(const_0_17_out));
	coreir_const #(
		.value(32'h00000000),
		.width(32)
	) const_0_32(.out(const_0_32_out));
	coreir_wrap coreir_wrapInClock_inst0(
		.in(clk),
		.out(coreir_wrapInClock_inst0_out)
	);
	coreir_wrap coreir_wrapInClock_inst1(
		.in(clk),
		.out(coreir_wrapInClock_inst1_out)
	);
	coreir_wrap coreir_wrapInClock_inst2(
		.in(clk),
		.out(coreir_wrapInClock_inst2_out)
	);
	Or4x32 read_config_data_or_final(
		.I0(Tile_X00_Y04_read_config_data),
		.I1(Tile_X01_Y04_read_config_data),
		.I2(Tile_X02_Y04_read_config_data),
		.I3(Tile_X03_Y04_read_config_data),
		.O(read_config_data_or_final_O)
	);
	mantle_wire__typeBit4 self_stall(
		.in(stall),
		.out(self_stall_out)
	);
	assign glb2io_17_X00_Y00_ready = Tile_X00_Y00_glb2io_17_ready;
	assign glb2io_17_X01_Y00_ready = Tile_X01_Y00_glb2io_17_ready;
	assign glb2io_17_X02_Y00_ready = Tile_X02_Y00_glb2io_17_ready;
	assign glb2io_17_X03_Y00_ready = Tile_X03_Y00_glb2io_17_ready;
	assign glb2io_1_X00_Y00_ready = Tile_X00_Y00_glb2io_1_ready;
	assign glb2io_1_X01_Y00_ready = Tile_X01_Y00_glb2io_1_ready;
	assign glb2io_1_X02_Y00_ready = Tile_X02_Y00_glb2io_1_ready;
	assign glb2io_1_X03_Y00_ready = Tile_X03_Y00_glb2io_1_ready;
	assign io2glb_17_X00_Y00 = Tile_X00_Y00_io2glb_17;
	assign io2glb_17_X00_Y00_valid = Tile_X00_Y00_io2glb_17_valid;
	assign io2glb_17_X01_Y00 = Tile_X01_Y00_io2glb_17;
	assign io2glb_17_X01_Y00_valid = Tile_X01_Y00_io2glb_17_valid;
	assign io2glb_17_X02_Y00 = Tile_X02_Y00_io2glb_17;
	assign io2glb_17_X02_Y00_valid = Tile_X02_Y00_io2glb_17_valid;
	assign io2glb_17_X03_Y00 = Tile_X03_Y00_io2glb_17;
	assign io2glb_17_X03_Y00_valid = Tile_X03_Y00_io2glb_17_valid;
	assign io2glb_1_X00_Y00 = Tile_X00_Y00_io2glb_1;
	assign io2glb_1_X00_Y00_valid = Tile_X00_Y00_io2glb_1_valid;
	assign io2glb_1_X01_Y00 = Tile_X01_Y00_io2glb_1;
	assign io2glb_1_X01_Y00_valid = Tile_X01_Y00_io2glb_1_valid;
	assign io2glb_1_X02_Y00 = Tile_X02_Y00_io2glb_1;
	assign io2glb_1_X02_Y00_valid = Tile_X02_Y00_io2glb_1_valid;
	assign io2glb_1_X03_Y00 = Tile_X03_Y00_io2glb_1;
	assign io2glb_1_X03_Y00_valid = Tile_X03_Y00_io2glb_1_valid;
	assign read_config_data = read_config_data_or_final_O;
endmodule
module Garnet (
	axi4_slave_araddr,
	axi4_slave_arready,
	axi4_slave_arvalid,
	axi4_slave_awaddr,
	axi4_slave_awready,
	axi4_slave_awvalid,
	axi4_slave_bready,
	axi4_slave_bresp,
	axi4_slave_bvalid,
	axi4_slave_rdata,
	axi4_slave_rready,
	axi4_slave_rresp,
	axi4_slave_rvalid,
	axi4_slave_wdata,
	axi4_slave_wready,
	axi4_slave_wvalid,
	cgra_running_clk_out,
	clk_in,
	interrupt,
	jtag_tck,
	jtag_tdi,
	jtag_tdo,
	jtag_tms,
	jtag_trst_n,
	proc_packet_rd_addr,
	proc_packet_rd_data,
	proc_packet_rd_data_valid,
	proc_packet_rd_en,
	proc_packet_wr_addr,
	proc_packet_wr_data,
	proc_packet_wr_en,
	proc_packet_wr_strb,
	reset_in
);
	input [12:0] axi4_slave_araddr;
	output wire axi4_slave_arready;
	input axi4_slave_arvalid;
	input [12:0] axi4_slave_awaddr;
	output wire axi4_slave_awready;
	input axi4_slave_awvalid;
	input axi4_slave_bready;
	output wire [1:0] axi4_slave_bresp;
	output wire axi4_slave_bvalid;
	output wire [31:0] axi4_slave_rdata;
	input axi4_slave_rready;
	output wire [1:0] axi4_slave_rresp;
	output wire axi4_slave_rvalid;
	input [31:0] axi4_slave_wdata;
	output wire axi4_slave_wready;
	input axi4_slave_wvalid;
	output wire cgra_running_clk_out;
	input clk_in;
	output wire interrupt;
	input jtag_tck;
	input jtag_tdi;
	output wire jtag_tdo;
	input jtag_tms;
	input jtag_trst_n;
	input [18:0] proc_packet_rd_addr;
	output wire [63:0] proc_packet_rd_data;
	output wire proc_packet_rd_data_valid;
	input proc_packet_rd_en;
	input [18:0] proc_packet_wr_addr;
	input [63:0] proc_packet_wr_data;
	input proc_packet_wr_en;
	input [7:0] proc_packet_wr_strb;
	input reset_in;
	wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_clk_out;
	wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_reset_out;
	wire [3:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_stall;
	wire [1:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_clk_en_master;
	wire [1:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_clk_en_bank_master;
	wire [1:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_pcfg_broadcast_stall;
	wire [0:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_flush_crossbar_sel;
	wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_en;
	wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_clk_en;
	wire [11:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_addr;
	wire [31:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_data;
	wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_rd_en;
	wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_rd_clk_en;
	wire [11:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_rd_addr;
	wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_wr_en;
	wire [18:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_wr_addr;
	wire [31:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_wr_data;
	wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_rd_en;
	wire [18:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_rd_addr;
	wire [1:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_strm_g2f_start_pulse;
	wire [1:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_strm_f2g_start_pulse;
	wire [1:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_pc_start_pulse;
	wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_read;
	wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_write;
	wire [31:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_addr;
	wire [31:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_wr_data;
	wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_awready;
	wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_wready;
	wire [1:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_bresp;
	wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_bvalid;
	wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_arready;
	wire [31:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_rdata;
	wire [1:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_rresp;
	wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_rvalid;
	wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_interrupt;
	wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_tdo;
	wire Interconnect_inst0_glb2io_17_X00_Y00_ready;
	wire Interconnect_inst0_glb2io_17_X01_Y00_ready;
	wire Interconnect_inst0_glb2io_17_X02_Y00_ready;
	wire Interconnect_inst0_glb2io_17_X03_Y00_ready;
	wire Interconnect_inst0_glb2io_1_X00_Y00_ready;
	wire Interconnect_inst0_glb2io_1_X01_Y00_ready;
	wire Interconnect_inst0_glb2io_1_X02_Y00_ready;
	wire Interconnect_inst0_glb2io_1_X03_Y00_ready;
	wire [16:0] Interconnect_inst0_io2glb_17_X00_Y00_unq1;
	wire Interconnect_inst0_io2glb_17_X00_Y00_valid;
	wire [16:0] Interconnect_inst0_io2glb_17_X01_Y00_unq1;
	wire Interconnect_inst0_io2glb_17_X01_Y00_valid;
	wire [16:0] Interconnect_inst0_io2glb_17_X02_Y00_unq1;
	wire Interconnect_inst0_io2glb_17_X02_Y00_valid;
	wire [16:0] Interconnect_inst0_io2glb_17_X03_Y00_unq1;
	wire Interconnect_inst0_io2glb_17_X03_Y00_valid;
	wire [0:0] Interconnect_inst0_io2glb_1_X00_Y00;
	wire Interconnect_inst0_io2glb_1_X00_Y00_valid;
	wire [0:0] Interconnect_inst0_io2glb_1_X01_Y00;
	wire Interconnect_inst0_io2glb_1_X01_Y00_valid;
	wire [0:0] Interconnect_inst0_io2glb_1_X02_Y00;
	wire Interconnect_inst0_io2glb_1_X02_Y00_valid;
	wire [0:0] Interconnect_inst0_io2glb_1_X03_Y00;
	wire Interconnect_inst0_io2glb_1_X03_Y00_valid;
	wire [31:0] Interconnect_inst0_read_config_data;
	wire [16:0] Interconnect_inst0_glb2io_17_X00_Y00_in;
	wire [16:0] Interconnect_inst0_glb2io_17_X01_Y00_in;
	wire [16:0] Interconnect_inst0_glb2io_17_X02_Y00_in;
	wire [16:0] Interconnect_inst0_glb2io_17_X03_Y00_in;
	wire [16:0] Interconnect_inst0_io2glb_17_X00_Y00_out;
	wire [16:0] Interconnect_inst0_io2glb_17_X01_Y00_out;
	wire [16:0] Interconnect_inst0_io2glb_17_X02_Y00_out;
	wire [16:0] Interconnect_inst0_io2glb_17_X03_Y00_out;
	wire bit_const_0_None_out;
	wire bit_const_1_None_out;
	wire [63:0] global_buffer_W_inst0_proc_rd_data;
	wire [0:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_1_0;
	wire [15:0] global_buffer_W_inst0_strm_data_g2f_0_0;
	wire [15:0] global_buffer_W_inst0_strm_data_g2f_1_1;
	wire [0:0] global_buffer_W_inst0_if_sram_cfg_rd_data_valid;
	wire [3:0] global_buffer_W_inst0_cgra_stall;
	wire [1:0] global_buffer_W_inst0_strm_g2f_interrupt_pulse;
	wire [31:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_1_1;
	wire [0:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_1_1;
	wire [0:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_1_0;
	wire [0:0] global_buffer_W_inst0_strm_data_f2g_rdy_0_0;
	wire [0:0] global_buffer_W_inst0_strm_ctrl_g2f_1_1;
	wire [0:0] global_buffer_W_inst0_strm_data_flush_g2f;
	wire [0:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_0_1;
	wire [31:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_1_0;
	wire [0:0] global_buffer_W_inst0_strm_data_g2f_vld_1_0;
	wire [31:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_0_0;
	wire [31:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_0_1;
	wire [31:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_0_0;
	wire [0:0] global_buffer_W_inst0_strm_data_f2g_rdy_0_1;
	wire [1:0] global_buffer_W_inst0_pcfg_g2f_interrupt_pulse;
	wire [0:0] global_buffer_W_inst0_strm_ctrl_g2f_0_0;
	wire [0:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_0_1;
	wire [15:0] global_buffer_W_inst0_strm_data_g2f_1_0;
	wire [0:0] global_buffer_W_inst0_strm_data_g2f_vld_1_1;
	wire [15:0] global_buffer_W_inst0_strm_data_g2f_0_1;
	wire [0:0] global_buffer_W_inst0_strm_data_g2f_vld_0_0;
	wire [0:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_0_0;
	wire [31:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_1_0;
	wire [31:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_1_1;
	wire [0:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_0_0;
	wire [0:0] global_buffer_W_inst0_strm_data_f2g_rdy_1_0;
	wire [0:0] global_buffer_W_inst0_strm_ctrl_g2f_1_0;
	wire [31:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_0_1;
	wire [0:0] global_buffer_W_inst0_if_cfg_rd_data_valid;
	wire [0:0] global_buffer_W_inst0_strm_data_f2g_rdy_1_1;
	wire [0:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_1_1;
	wire [31:0] global_buffer_W_inst0_if_sram_cfg_rd_data;
	wire [1:0] global_buffer_W_inst0_strm_f2g_interrupt_pulse;
	wire [0:0] global_buffer_W_inst0_strm_data_g2f_vld_0_1;
	wire [31:0] global_buffer_W_inst0_if_cfg_rd_data;
	wire [0:0] global_buffer_W_inst0_proc_rd_data_valid;
	wire [0:0] global_buffer_W_inst0_strm_ctrl_g2f_0_1;
	global_controller GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0(
		.clk_in(clk_in),
		.reset_in(reset_in),
		.clk_out(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_clk_out),
		.reset_out(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_reset_out),
		.cgra_stall(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_stall),
		.glb_clk_en_master(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_clk_en_master),
		.glb_clk_en_bank_master(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_clk_en_bank_master),
		.glb_pcfg_broadcast_stall(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_pcfg_broadcast_stall),
		.glb_flush_crossbar_sel(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_flush_crossbar_sel),
		.glb_cfg_wr_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_en),
		.glb_cfg_wr_clk_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_clk_en),
		.glb_cfg_wr_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_addr),
		.glb_cfg_wr_data(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_data),
		.glb_cfg_rd_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_rd_en),
		.glb_cfg_rd_clk_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_rd_clk_en),
		.glb_cfg_rd_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_rd_addr),
		.glb_cfg_rd_data(global_buffer_W_inst0_if_cfg_rd_data),
		.glb_cfg_rd_data_valid(global_buffer_W_inst0_if_cfg_rd_data_valid[0]),
		.sram_cfg_wr_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_wr_en),
		.sram_cfg_wr_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_wr_addr),
		.sram_cfg_wr_data(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_wr_data),
		.sram_cfg_rd_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_rd_en),
		.sram_cfg_rd_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_rd_addr),
		.sram_cfg_rd_data(global_buffer_W_inst0_if_sram_cfg_rd_data),
		.sram_cfg_rd_data_valid(global_buffer_W_inst0_if_sram_cfg_rd_data_valid[0]),
		.strm_g2f_start_pulse(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_strm_g2f_start_pulse),
		.strm_f2g_start_pulse(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_strm_f2g_start_pulse),
		.pc_start_pulse(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_pc_start_pulse),
		.strm_g2f_interrupt_pulse(global_buffer_W_inst0_strm_g2f_interrupt_pulse),
		.strm_f2g_interrupt_pulse(global_buffer_W_inst0_strm_f2g_interrupt_pulse),
		.pcfg_g2f_interrupt_pulse(global_buffer_W_inst0_pcfg_g2f_interrupt_pulse),
		.cgra_cfg_read(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_read),
		.cgra_cfg_write(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_write),
		.cgra_cfg_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_addr),
		.cgra_cfg_wr_data(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_wr_data),
		.cgra_cfg_rd_data(Interconnect_inst0_read_config_data),
		.axi_awaddr(axi4_slave_awaddr),
		.axi_awvalid(axi4_slave_awvalid),
		.axi_awready(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_awready),
		.axi_wdata(axi4_slave_wdata),
		.axi_wvalid(axi4_slave_wvalid),
		.axi_wready(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_wready),
		.axi_bready(axi4_slave_bready),
		.axi_bresp(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_bresp),
		.axi_bvalid(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_bvalid),
		.axi_araddr(axi4_slave_araddr),
		.axi_arvalid(axi4_slave_arvalid),
		.axi_arready(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_arready),
		.axi_rdata(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_rdata),
		.axi_rresp(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_rresp),
		.axi_rvalid(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_rvalid),
		.axi_rready(axi4_slave_rready),
		.interrupt(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_interrupt),
		.tck(jtag_tck),
		.tdi(jtag_tdi),
		.tms(jtag_tms),
		.trst_n(jtag_trst_n),
		.tdo(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_tdo)
	);
	Interconnect Interconnect_inst0(
		.clk(clk_in),
		.config_0_config_addr(global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_0_0),
		.config_0_config_data(global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_0_0),
		.config_0_read(global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_0_0),
		.config_0_write(global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_0_0),
		.config_1_config_addr(global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_0_1),
		.config_1_config_data(global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_0_1),
		.config_1_read(global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_0_1),
		.config_1_write(global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_0_1),
		.config_2_config_addr(global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_1_0),
		.config_2_config_data(global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_1_0),
		.config_2_read(global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_1_0),
		.config_2_write(global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_1_0),
		.config_3_config_addr(global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_1_1),
		.config_3_config_data(global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_1_1),
		.config_3_read(global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_1_1),
		.config_3_write(global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_1_1),
		.flush(global_buffer_W_inst0_strm_data_flush_g2f),
		.glb2io_17_X00_Y00(Interconnect_inst0_glb2io_17_X00_Y00_in),
		.glb2io_17_X00_Y00_ready(Interconnect_inst0_glb2io_17_X00_Y00_ready),
		.glb2io_17_X00_Y00_valid(global_buffer_W_inst0_strm_data_g2f_vld_0_0[0]),
		.glb2io_17_X01_Y00(Interconnect_inst0_glb2io_17_X01_Y00_in),
		.glb2io_17_X01_Y00_ready(Interconnect_inst0_glb2io_17_X01_Y00_ready),
		.glb2io_17_X01_Y00_valid(global_buffer_W_inst0_strm_data_g2f_vld_0_1[0]),
		.glb2io_17_X02_Y00(Interconnect_inst0_glb2io_17_X02_Y00_in),
		.glb2io_17_X02_Y00_ready(Interconnect_inst0_glb2io_17_X02_Y00_ready),
		.glb2io_17_X02_Y00_valid(global_buffer_W_inst0_strm_data_g2f_vld_1_0[0]),
		.glb2io_17_X03_Y00(Interconnect_inst0_glb2io_17_X03_Y00_in),
		.glb2io_17_X03_Y00_ready(Interconnect_inst0_glb2io_17_X03_Y00_ready),
		.glb2io_17_X03_Y00_valid(global_buffer_W_inst0_strm_data_g2f_vld_1_1[0]),
		.glb2io_1_X00_Y00(global_buffer_W_inst0_strm_ctrl_g2f_0_0),
		.glb2io_1_X00_Y00_ready(Interconnect_inst0_glb2io_1_X00_Y00_ready),
		.glb2io_1_X00_Y00_valid(bit_const_1_None_out),
		.glb2io_1_X01_Y00(global_buffer_W_inst0_strm_ctrl_g2f_0_1),
		.glb2io_1_X01_Y00_ready(Interconnect_inst0_glb2io_1_X01_Y00_ready),
		.glb2io_1_X01_Y00_valid(bit_const_1_None_out),
		.glb2io_1_X02_Y00(global_buffer_W_inst0_strm_ctrl_g2f_1_0),
		.glb2io_1_X02_Y00_ready(Interconnect_inst0_glb2io_1_X02_Y00_ready),
		.glb2io_1_X02_Y00_valid(bit_const_1_None_out),
		.glb2io_1_X03_Y00(global_buffer_W_inst0_strm_ctrl_g2f_1_1),
		.glb2io_1_X03_Y00_ready(Interconnect_inst0_glb2io_1_X03_Y00_ready),
		.glb2io_1_X03_Y00_valid(bit_const_1_None_out),
		.io2glb_17_X00_Y00(Interconnect_inst0_io2glb_17_X00_Y00_unq1),
		.io2glb_17_X00_Y00_ready(global_buffer_W_inst0_strm_data_f2g_rdy_0_0[0]),
		.io2glb_17_X00_Y00_valid(Interconnect_inst0_io2glb_17_X00_Y00_valid),
		.io2glb_17_X01_Y00(Interconnect_inst0_io2glb_17_X01_Y00_unq1),
		.io2glb_17_X01_Y00_ready(global_buffer_W_inst0_strm_data_f2g_rdy_0_1[0]),
		.io2glb_17_X01_Y00_valid(Interconnect_inst0_io2glb_17_X01_Y00_valid),
		.io2glb_17_X02_Y00(Interconnect_inst0_io2glb_17_X02_Y00_unq1),
		.io2glb_17_X02_Y00_ready(global_buffer_W_inst0_strm_data_f2g_rdy_1_0[0]),
		.io2glb_17_X02_Y00_valid(Interconnect_inst0_io2glb_17_X02_Y00_valid),
		.io2glb_17_X03_Y00(Interconnect_inst0_io2glb_17_X03_Y00_unq1),
		.io2glb_17_X03_Y00_ready(global_buffer_W_inst0_strm_data_f2g_rdy_1_1[0]),
		.io2glb_17_X03_Y00_valid(Interconnect_inst0_io2glb_17_X03_Y00_valid),
		.io2glb_1_X00_Y00(Interconnect_inst0_io2glb_1_X00_Y00),
		.io2glb_1_X00_Y00_ready(bit_const_1_None_out),
		.io2glb_1_X00_Y00_valid(Interconnect_inst0_io2glb_1_X00_Y00_valid),
		.io2glb_1_X01_Y00(Interconnect_inst0_io2glb_1_X01_Y00),
		.io2glb_1_X01_Y00_ready(bit_const_1_None_out),
		.io2glb_1_X01_Y00_valid(Interconnect_inst0_io2glb_1_X01_Y00_valid),
		.io2glb_1_X02_Y00(Interconnect_inst0_io2glb_1_X02_Y00),
		.io2glb_1_X02_Y00_ready(bit_const_1_None_out),
		.io2glb_1_X02_Y00_valid(Interconnect_inst0_io2glb_1_X02_Y00_valid),
		.io2glb_1_X03_Y00(Interconnect_inst0_io2glb_1_X03_Y00),
		.io2glb_1_X03_Y00_ready(bit_const_1_None_out),
		.io2glb_1_X03_Y00_valid(Interconnect_inst0_io2glb_1_X03_Y00_valid),
		.read_config_data(Interconnect_inst0_read_config_data),
		.reset(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_reset_out),
		.stall(global_buffer_W_inst0_cgra_stall)
	);
	wire [16:0] Interconnect_inst0_glb2io_17_X00_Y00_out;
	assign Interconnect_inst0_glb2io_17_X00_Y00_out = {bit_const_0_None_out, global_buffer_W_inst0_strm_data_g2f_0_0};
	mantle_wire__typeBitIn17 Interconnect_inst0_glb2io_17_X00_Y00(
		.in(Interconnect_inst0_glb2io_17_X00_Y00_in),
		.out(Interconnect_inst0_glb2io_17_X00_Y00_out)
	);
	wire [16:0] Interconnect_inst0_glb2io_17_X01_Y00_out;
	assign Interconnect_inst0_glb2io_17_X01_Y00_out = {bit_const_0_None_out, global_buffer_W_inst0_strm_data_g2f_0_1};
	mantle_wire__typeBitIn17 Interconnect_inst0_glb2io_17_X01_Y00(
		.in(Interconnect_inst0_glb2io_17_X01_Y00_in),
		.out(Interconnect_inst0_glb2io_17_X01_Y00_out)
	);
	wire [16:0] Interconnect_inst0_glb2io_17_X02_Y00_out;
	assign Interconnect_inst0_glb2io_17_X02_Y00_out = {bit_const_0_None_out, global_buffer_W_inst0_strm_data_g2f_1_0};
	mantle_wire__typeBitIn17 Interconnect_inst0_glb2io_17_X02_Y00(
		.in(Interconnect_inst0_glb2io_17_X02_Y00_in),
		.out(Interconnect_inst0_glb2io_17_X02_Y00_out)
	);
	wire [16:0] Interconnect_inst0_glb2io_17_X03_Y00_out;
	assign Interconnect_inst0_glb2io_17_X03_Y00_out = {bit_const_0_None_out, global_buffer_W_inst0_strm_data_g2f_1_1};
	mantle_wire__typeBitIn17 Interconnect_inst0_glb2io_17_X03_Y00(
		.in(Interconnect_inst0_glb2io_17_X03_Y00_in),
		.out(Interconnect_inst0_glb2io_17_X03_Y00_out)
	);
	mantle_wire__typeBit17 Interconnect_inst0_io2glb_17_X00_Y00(
		.in(Interconnect_inst0_io2glb_17_X00_Y00_unq1),
		.out(Interconnect_inst0_io2glb_17_X00_Y00_out)
	);
	mantle_wire__typeBit17 Interconnect_inst0_io2glb_17_X01_Y00(
		.in(Interconnect_inst0_io2glb_17_X01_Y00_unq1),
		.out(Interconnect_inst0_io2glb_17_X01_Y00_out)
	);
	mantle_wire__typeBit17 Interconnect_inst0_io2glb_17_X02_Y00(
		.in(Interconnect_inst0_io2glb_17_X02_Y00_unq1),
		.out(Interconnect_inst0_io2glb_17_X02_Y00_out)
	);
	mantle_wire__typeBit17 Interconnect_inst0_io2glb_17_X03_Y00(
		.in(Interconnect_inst0_io2glb_17_X03_Y00_unq1),
		.out(Interconnect_inst0_io2glb_17_X03_Y00_out)
	);
	corebit_const #(.value(1'b0)) bit_const_0_None(.out(bit_const_0_None_out));
	corebit_const #(.value(1'b1)) bit_const_1_None(.out(bit_const_1_None_out));
	global_buffer_W global_buffer_W_inst0(
		.cgra_cfg_jtag_gc2glb_data(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_wr_data),
		.proc_rd_data(global_buffer_W_inst0_proc_rd_data),
		.if_sram_cfg_wr_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_wr_addr),
		.cgra_cfg_g2f_cfg_wr_en_1_0(global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_1_0),
		.proc_wr_en(proc_packet_wr_en),
		.strm_data_g2f_0_0(global_buffer_W_inst0_strm_data_g2f_0_0),
		.strm_g2f_start_pulse(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_strm_g2f_start_pulse),
		.strm_data_g2f_1_1(global_buffer_W_inst0_strm_data_g2f_1_1),
		.if_sram_cfg_rd_data_valid(global_buffer_W_inst0_if_sram_cfg_rd_data_valid),
		.cgra_stall(global_buffer_W_inst0_cgra_stall),
		.if_cfg_wr_data(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_data),
		.cgra_stall_in(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_stall),
		.strm_g2f_interrupt_pulse(global_buffer_W_inst0_strm_g2f_interrupt_pulse),
		.proc_rd_addr(proc_packet_rd_addr),
		.strm_data_g2f_rdy_1_1(Interconnect_inst0_glb2io_17_X03_Y00_ready),
		.cgra_cfg_g2f_cfg_data_1_1(global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_1_1),
		.cgra_cfg_g2f_cfg_wr_en_1_1(global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_1_1),
		.strm_data_f2g_1_0(Interconnect_inst0_io2glb_17_X02_Y00_out[15:0]),
		.cgra_cfg_g2f_cfg_rd_en_1_0(global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_1_0),
		.strm_data_f2g_rdy_0_0(global_buffer_W_inst0_strm_data_f2g_rdy_0_0),
		.strm_ctrl_g2f_1_1(global_buffer_W_inst0_strm_ctrl_g2f_1_1),
		.strm_data_f2g_1_1(Interconnect_inst0_io2glb_17_X03_Y00_out[15:0]),
		.strm_data_flush_g2f(global_buffer_W_inst0_strm_data_flush_g2f),
		.cgra_cfg_g2f_cfg_rd_en_0_1(global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_0_1),
		.cgra_cfg_g2f_cfg_addr_1_0(global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_1_0),
		.strm_data_f2g_vld_1_1(Interconnect_inst0_io2glb_17_X03_Y00_valid),
		.glb_clk_en_master(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_clk_en_master),
		.if_sram_cfg_wr_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_wr_en),
		.strm_ctrl_f2g_0_0(Interconnect_inst0_io2glb_1_X00_Y00),
		.strm_f2g_start_pulse(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_strm_f2g_start_pulse),
		.strm_data_f2g_vld_0_0(Interconnect_inst0_io2glb_17_X00_Y00_valid),
		.strm_data_g2f_vld_1_0(global_buffer_W_inst0_strm_data_g2f_vld_1_0),
		.strm_data_g2f_rdy_0_0(Interconnect_inst0_glb2io_17_X00_Y00_ready),
		.if_sram_cfg_wr_data(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_wr_data),
		.cgra_cfg_g2f_cfg_data_0_0(global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_0_0),
		.cgra_cfg_g2f_cfg_data_0_1(global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_0_1),
		.clk(clk_in),
		.cgra_cfg_g2f_cfg_addr_0_0(global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_0_0),
		.strm_data_f2g_vld_1_0(Interconnect_inst0_io2glb_17_X02_Y00_valid),
		.strm_data_f2g_vld_0_1(Interconnect_inst0_io2glb_17_X01_Y00_valid),
		.strm_data_f2g_rdy_0_1(global_buffer_W_inst0_strm_data_f2g_rdy_0_1),
		.pcfg_g2f_interrupt_pulse(global_buffer_W_inst0_pcfg_g2f_interrupt_pulse),
		.strm_ctrl_g2f_0_0(global_buffer_W_inst0_strm_ctrl_g2f_0_0),
		.cgra_cfg_g2f_cfg_wr_en_0_1(global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_0_1),
		.strm_data_g2f_rdy_0_1(Interconnect_inst0_glb2io_17_X01_Y00_ready),
		.strm_data_g2f_1_0(global_buffer_W_inst0_strm_data_g2f_1_0),
		.strm_data_g2f_vld_1_1(global_buffer_W_inst0_strm_data_g2f_vld_1_1),
		.if_cfg_wr_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_addr),
		.proc_rd_en(proc_packet_rd_en),
		.strm_data_g2f_0_1(global_buffer_W_inst0_strm_data_g2f_0_1),
		.pcfg_broadcast_stall(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_pcfg_broadcast_stall),
		.if_cfg_rd_clk_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_rd_clk_en),
		.reset(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_reset_out),
		.flush_crossbar_sel(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_flush_crossbar_sel),
		.strm_data_g2f_vld_0_0(global_buffer_W_inst0_strm_data_g2f_vld_0_0),
		.if_cfg_rd_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_rd_en),
		.strm_data_f2g_0_1(Interconnect_inst0_io2glb_17_X01_Y00_out[15:0]),
		.pcfg_start_pulse(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_pc_start_pulse),
		.cgra_cfg_g2f_cfg_rd_en_0_0(global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_0_0),
		.cgra_cfg_g2f_cfg_data_1_0(global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_1_0),
		.if_cfg_wr_clk_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_clk_en),
		.cgra_cfg_g2f_cfg_addr_1_1(global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_1_1),
		.strm_ctrl_f2g_0_1(Interconnect_inst0_io2glb_1_X01_Y00),
		.proc_wr_data(proc_packet_wr_data),
		.cgra_cfg_g2f_cfg_wr_en_0_0(global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_0_0),
		.strm_data_g2f_rdy_1_0(Interconnect_inst0_glb2io_17_X02_Y00_ready),
		.strm_data_f2g_rdy_1_0(global_buffer_W_inst0_strm_data_f2g_rdy_1_0),
		.strm_ctrl_g2f_1_0(global_buffer_W_inst0_strm_ctrl_g2f_1_0),
		.cgra_cfg_jtag_gc2glb_rd_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_read),
		.proc_wr_strb(proc_packet_wr_strb),
		.glb_clk_en_bank_master(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_clk_en_bank_master),
		.if_sram_cfg_rd_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_rd_en),
		.proc_wr_addr(proc_packet_wr_addr),
		.cgra_cfg_g2f_cfg_addr_0_1(global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_0_1),
		.if_cfg_rd_data_valid(global_buffer_W_inst0_if_cfg_rd_data_valid),
		.strm_data_f2g_rdy_1_1(global_buffer_W_inst0_strm_data_f2g_rdy_1_1),
		.cgra_cfg_g2f_cfg_rd_en_1_1(global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_1_1),
		.strm_ctrl_f2g_1_0(Interconnect_inst0_io2glb_1_X02_Y00),
		.if_sram_cfg_rd_data(global_buffer_W_inst0_if_sram_cfg_rd_data),
		.if_cfg_rd_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_rd_addr),
		.cgra_cfg_jtag_gc2glb_wr_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_write),
		.strm_ctrl_f2g_1_1(Interconnect_inst0_io2glb_1_X03_Y00),
		.strm_f2g_interrupt_pulse(global_buffer_W_inst0_strm_f2g_interrupt_pulse),
		.strm_data_g2f_vld_0_1(global_buffer_W_inst0_strm_data_g2f_vld_0_1),
		.cgra_cfg_jtag_gc2glb_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_addr),
		.strm_data_f2g_0_0(Interconnect_inst0_io2glb_17_X00_Y00_out[15:0]),
		.if_cfg_wr_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_en),
		.if_cfg_rd_data(global_buffer_W_inst0_if_cfg_rd_data),
		.if_sram_cfg_rd_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_rd_addr),
		.proc_rd_data_valid(global_buffer_W_inst0_proc_rd_data_valid),
		.strm_ctrl_g2f_0_1(global_buffer_W_inst0_strm_ctrl_g2f_0_1)
	);
	assign axi4_slave_arready = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_arready;
	assign axi4_slave_awready = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_awready;
	assign axi4_slave_bresp = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_bresp;
	assign axi4_slave_bvalid = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_bvalid;
	assign axi4_slave_rdata = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_rdata;
	assign axi4_slave_rresp = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_rresp;
	assign axi4_slave_rvalid = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_rvalid;
	assign axi4_slave_wready = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_wready;
	assign cgra_running_clk_out = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_clk_out;
	assign interrupt = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_interrupt;
	assign jtag_tdo = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_tdo;
	assign proc_packet_rd_data = global_buffer_W_inst0_proc_rd_data;
	assign proc_packet_rd_data_valid = global_buffer_W_inst0_proc_rd_data_valid[0];
endmodule
module AN_CELL (
	A1,
	A2,
	Z
);
	input wire A1;
	input wire A2;
	output wire Z;
	assign Z = A1 & A2;
endmodule
module AO_CELL (
	A1,
	A2,
	B1,
	B2,
	Z
);
	input wire A1;
	input wire A2;
	input wire B1;
	input wire B2;
	output wire Z;
	assign Z = (A1 & A2) | (B1 & B2);
endmodule
module PEGEN_mul_hack (
	a,
	b,
	rnd,
	z,
	status
);
	parameter exp_bits = 1;
	parameter frac_bits = 1;
	parameter ieee_compliance = 1;
	input [exp_bits + frac_bits:0] a;
	input [exp_bits + frac_bits:0] b;
	input [2:0] rnd;
	output wire [exp_bits + frac_bits:0] z;
	output wire [7:0] status;
	wire [exp_bits + frac_bits:0] int_out;
	wire [2:0] results_x;
	reg sign;
	reg [exp_bits - 1:0] exp;
	reg [frac_bits:0] frac;
	CW_fp_mult #(
		.sig_width(frac_bits + 3),
		.exp_width(exp_bits),
		.ieee_compliance(ieee_compliance)
	) mul1(
		.a({a, 3'h0}),
		.b({b, 3'h0}),
		.rnd(rnd),
		.z({int_out, results_x}),
		.status(status)
	);
	always @(*) begin
		sign = int_out[exp_bits + frac_bits];
		exp = int_out[(exp_bits + frac_bits) - 1:frac_bits];
		frac = {1'b0, int_out[frac_bits - 1:0]};
		if ((results_x[2] & (results_x[1] | results_x[0])) | (int_out[0] & results_x[2])) begin
			frac = frac + 1'd1;
			if (~&exp)
				exp = exp + {{exp_bits - 1 {1'b0}}, frac[frac_bits]};
		end
	end
	assign z = {sign, exp, frac[frac_bits - 1:0]};
endmodule
module PEGEN_add (
	a,
	b,
	rnd,
	z,
	status
);
	parameter exp_bits = 1;
	parameter frac_bits = 1;
	parameter ieee_compliance = 1;
	input [exp_bits + frac_bits:0] a;
	input [exp_bits + frac_bits:0] b;
	input [2:0] rnd;
	output wire [exp_bits + frac_bits:0] z;
	output wire [7:0] status;
	CW_fp_add #(
		.sig_width(frac_bits),
		.exp_width(exp_bits),
		.ieee_compliance(ieee_compliance)
	) add_inst(
		.a(a),
		.b(b),
		.rnd(rnd),
		.z(z),
		.status(status)
	);
endmodule
module PEGEN_coreir_xor (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output wire [width - 1:0] out;
	assign out = in0 ^ in1;
endmodule
module PEGEN_coreir_ule (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output wire out;
	assign out = in0 <= in1;
endmodule
module PEGEN_coreir_ugt (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output wire out;
	assign out = in0 > in1;
endmodule
module PEGEN_coreir_uge (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output wire out;
	assign out = in0 >= in1;
endmodule
module PEGEN_coreir_sub (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output wire [width - 1:0] out;
	assign out = in0 - in1;
endmodule
module PEGEN_coreir_slt (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output wire out;
	assign out = $signed(in0) < $signed(in1);
endmodule
module PEGEN_coreir_sle (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output wire out;
	assign out = $signed(in0) <= $signed(in1);
endmodule
module PEGEN_coreir_shl (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output wire [width - 1:0] out;
	assign out = in0 << in1;
endmodule
module PEGEN_coreir_sge (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output wire out;
	assign out = $signed(in0) >= $signed(in1);
endmodule
module PEGEN_coreir_reg_arst (
	clk,
	arst,
	in,
	out
);
	parameter width = 1;
	parameter arst_posedge = 1;
	parameter clk_posedge = 1;
	parameter init = 1;
	input clk;
	input arst;
	input [width - 1:0] in;
	output wire [width - 1:0] out;
	reg [width - 1:0] outReg;
	wire real_rst;
	assign real_rst = (arst_posedge ? arst : ~arst);
	wire real_clk;
	assign real_clk = (clk_posedge ? clk : ~clk);
	always @(posedge real_clk or posedge real_rst)
		if (real_rst)
			outReg <= init;
		else
			outReg <= in;
	assign out = outReg;
endmodule
module PEGEN_coreir_or (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output wire [width - 1:0] out;
	assign out = in0 | in1;
endmodule
module PEGEN_coreir_not (
	in,
	out
);
	parameter width = 1;
	input [width - 1:0] in;
	output wire [width - 1:0] out;
	assign out = ~in;
endmodule
module PEGEN_coreir_neg (
	in,
	out
);
	parameter width = 1;
	input [width - 1:0] in;
	output wire [width - 1:0] out;
	assign out = -in;
endmodule
module PEGEN_coreir_mux (
	in0,
	in1,
	sel,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	input sel;
	output wire [width - 1:0] out;
	assign out = (sel ? in1 : in0);
endmodule
module PEGEN_coreir_mul (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output wire [width - 1:0] out;
	assign out = in0 * in1;
endmodule
module PEGEN_coreir_lshr (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output wire [width - 1:0] out;
	assign out = in0 >> in1;
endmodule
module PEGEN_coreir_eq (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output wire out;
	assign out = in0 == in1;
endmodule
module PEGEN_coreir_const (out);
	parameter width = 1;
	parameter value = 1;
	output wire [width - 1:0] out;
	assign out = value;
endmodule
module PEGEN_float_mul__exp_bits8__frac_bits7 (
	in0,
	in1,
	out
);
	input [15:0] in0;
	input [15:0] in1;
	output wire [15:0] out;
	wire [2:0] _$_U1_out;
	wire [15:0] mi_z;
	wire [7:0] mi_status;
	PEGEN_coreir_const #(
		.value(3'h1),
		.width(3)
	) _$_U1(.out(_$_U1_out));
	PEGEN_mul_hack #(
		.exp_bits(8),
		.frac_bits(7),
		.ieee_compliance(1'b1)
	) mi(
		.a(in0),
		.b(in1),
		.rnd(_$_U1_out),
		.z(mi_z),
		.status(mi_status)
	);
	assign out = mi_z;
endmodule
module PEGEN_float_add__exp_bits8__frac_bits7 (
	in0,
	in1,
	out
);
	input [15:0] in0;
	input [15:0] in1;
	output wire [15:0] out;
	wire [2:0] _$_U0_out;
	wire [15:0] mi_z;
	wire [7:0] mi_status;
	PEGEN_coreir_const #(
		.value(3'h0),
		.width(3)
	) _$_U0(.out(_$_U0_out));
	PEGEN_add #(
		.exp_bits(8),
		.frac_bits(7),
		.ieee_compliance(1'b1)
	) mi(
		.a(in0),
		.b(in1),
		.rnd(_$_U0_out),
		.z(mi_z),
		.status(mi_status)
	);
	assign out = mi_z;
endmodule
module PEGEN_coreir_ashr (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output wire [width - 1:0] out;
	assign out = $signed(in0) >>> in1;
endmodule
module PEGEN_coreir_and (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output wire [width - 1:0] out;
	assign out = in0 & in1;
endmodule
module PEGEN_coreir_add (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output wire [width - 1:0] out;
	assign out = in0 + in1;
endmodule
module PEGEN_corebit_xor (
	in0,
	in1,
	out
);
	input in0;
	input in1;
	output wire out;
	assign out = in0 ^ in1;
endmodule
module PEGEN_corebit_or (
	in0,
	in1,
	out
);
	input in0;
	input in1;
	output wire out;
	assign out = in0 | in1;
endmodule
module PEGEN_corebit_not (
	in,
	out
);
	input in;
	output wire out;
	assign out = ~in;
endmodule
module PEGEN_corebit_const (out);
	parameter value = 1;
	output wire out;
	assign out = value;
endmodule
module PEGEN_corebit_and (
	in0,
	in1,
	out
);
	input in0;
	input in1;
	output wire out;
	assign out = in0 & in1;
endmodule
module PEGEN_commonlib_muxn__N2__width9 (
	in_data,
	in_sel,
	out
);
	input [17:0] in_data;
	input [0:0] in_sel;
	output wire [8:0] out;
	wire [8:0] _join_out;
	PEGEN_coreir_mux #(.width(9)) _join(
		.in0(in_data[0+:9]),
		.in1(in_data[9+:9]),
		.sel(in_sel[0]),
		.out(_join_out)
	);
	assign out = _join_out;
endmodule
module PEGEN_commonlib_muxn__N2__width8 (
	in_data,
	in_sel,
	out
);
	input [15:0] in_data;
	input [0:0] in_sel;
	output wire [7:0] out;
	wire [7:0] _join_out;
	PEGEN_coreir_mux #(.width(8)) _join(
		.in0(in_data[0+:8]),
		.in1(in_data[8+:8]),
		.sel(in_sel[0]),
		.out(_join_out)
	);
	assign out = _join_out;
endmodule
module PEGEN_commonlib_muxn__N2__width5 (
	in_data,
	in_sel,
	out
);
	input [9:0] in_data;
	input [0:0] in_sel;
	output wire [4:0] out;
	wire [4:0] _join_out;
	PEGEN_coreir_mux #(.width(5)) _join(
		.in0(in_data[0+:5]),
		.in1(in_data[5+:5]),
		.sel(in_sel[0]),
		.out(_join_out)
	);
	assign out = _join_out;
endmodule
module PEGEN_commonlib_muxn__N2__width32 (
	in_data,
	in_sel,
	out
);
	input [63:0] in_data;
	input [0:0] in_sel;
	output wire [31:0] out;
	wire [31:0] _join_out;
	PEGEN_coreir_mux #(.width(32)) _join(
		.in0(in_data[0+:32]),
		.in1(in_data[32+:32]),
		.sel(in_sel[0]),
		.out(_join_out)
	);
	assign out = _join_out;
endmodule
module PEGEN_commonlib_muxn__N2__width3 (
	in_data,
	in_sel,
	out
);
	input [5:0] in_data;
	input [0:0] in_sel;
	output wire [2:0] out;
	wire [2:0] _join_out;
	PEGEN_coreir_mux #(.width(3)) _join(
		.in0(in_data[0+:3]),
		.in1(in_data[3+:3]),
		.sel(in_sel[0]),
		.out(_join_out)
	);
	assign out = _join_out;
endmodule
module PEGEN_commonlib_muxn__N2__width23 (
	in_data,
	in_sel,
	out
);
	input [45:0] in_data;
	input [0:0] in_sel;
	output wire [22:0] out;
	wire [22:0] _join_out;
	PEGEN_coreir_mux #(.width(23)) _join(
		.in0(in_data[0+:23]),
		.in1(in_data[23+:23]),
		.sel(in_sel[0]),
		.out(_join_out)
	);
	assign out = _join_out;
endmodule
module PEGEN_commonlib_muxn__N2__width2 (
	in_data,
	in_sel,
	out
);
	input [3:0] in_data;
	input [0:0] in_sel;
	output wire [1:0] out;
	wire [1:0] _join_out;
	PEGEN_coreir_mux #(.width(2)) _join(
		.in0(in_data[0+:2]),
		.in1(in_data[2+:2]),
		.sel(in_sel[0]),
		.out(_join_out)
	);
	assign out = _join_out;
endmodule
module PEGEN_commonlib_muxn__N2__width16 (
	in_data,
	in_sel,
	out
);
	input [31:0] in_data;
	input [0:0] in_sel;
	output wire [15:0] out;
	wire [15:0] _join_out;
	PEGEN_coreir_mux #(.width(16)) _join(
		.in0(in_data[0+:16]),
		.in1(in_data[16+:16]),
		.sel(in_sel[0]),
		.out(_join_out)
	);
	assign out = _join_out;
endmodule
module PEGEN_commonlib_muxn__N2__width1 (
	in_data,
	in_sel,
	out
);
	input [1:0] in_data;
	input [0:0] in_sel;
	output wire [0:0] out;
	wire [0:0] _join_out;
	PEGEN_coreir_mux #(.width(1)) _join(
		.in0(in_data[0+:1]),
		.in1(in_data[1+:1]),
		.sel(in_sel[0]),
		.out(_join_out)
	);
	assign out = _join_out;
endmodule
module PEGEN_Op_unq1 (
	in0,
	in1,
	O,
	CLK,
	ASYNCRESET
);
	input [15:0] in0;
	input [15:0] in1;
	output wire [15:0] O;
	input CLK;
	input ASYNCRESET;
	wire [15:0] magma_BFloat_16_mul_inst0_out;
	PEGEN_float_mul__exp_bits8__frac_bits7 magma_BFloat_16_mul_inst0(
		.in0(in0),
		.in1(in1),
		.out(magma_BFloat_16_mul_inst0_out)
	);
	assign O = magma_BFloat_16_mul_inst0_out;
endmodule
module PEGEN_Op (
	in0,
	in1,
	O,
	CLK,
	ASYNCRESET
);
	input [15:0] in0;
	input [15:0] in1;
	output wire [15:0] O;
	input CLK;
	input ASYNCRESET;
	wire [15:0] magma_BFloat_16_add_inst0_out;
	PEGEN_float_add__exp_bits8__frac_bits7 magma_BFloat_16_add_inst0(
		.in0(in0),
		.in1(in1),
		.out(magma_BFloat_16_add_inst0_out)
	);
	assign O = magma_BFloat_16_add_inst0_out;
endmodule
module PEGEN_Mux2xUInt32 (
	I0,
	I1,
	S,
	O
);
	input [31:0] I0;
	input [31:0] I1;
	input S;
	output wire [31:0] O;
	wire [31:0] coreir_commonlib_mux2x32_inst0_out;
	wire [63:0] coreir_commonlib_mux2x32_inst0_in_data;
	assign coreir_commonlib_mux2x32_inst0_in_data[32+:32] = I1;
	assign coreir_commonlib_mux2x32_inst0_in_data[0+:32] = I0;
	PEGEN_commonlib_muxn__N2__width32 coreir_commonlib_mux2x32_inst0(
		.in_data(coreir_commonlib_mux2x32_inst0_in_data),
		.in_sel(S),
		.out(coreir_commonlib_mux2x32_inst0_out)
	);
	assign O = coreir_commonlib_mux2x32_inst0_out;
endmodule
module PEGEN_Mux2xUInt16 (
	I0,
	I1,
	S,
	O
);
	input [15:0] I0;
	input [15:0] I1;
	input S;
	output wire [15:0] O;
	wire [15:0] coreir_commonlib_mux2x16_inst0_out;
	wire [31:0] coreir_commonlib_mux2x16_inst0_in_data;
	assign coreir_commonlib_mux2x16_inst0_in_data[16+:16] = I1;
	assign coreir_commonlib_mux2x16_inst0_in_data[0+:16] = I0;
	PEGEN_commonlib_muxn__N2__width16 coreir_commonlib_mux2x16_inst0(
		.in_data(coreir_commonlib_mux2x16_inst0_in_data),
		.in_sel(S),
		.out(coreir_commonlib_mux2x16_inst0_out)
	);
	assign O = coreir_commonlib_mux2x16_inst0_out;
endmodule
module PEGEN_Mux2xSInt9 (
	I0,
	I1,
	S,
	O
);
	input [8:0] I0;
	input [8:0] I1;
	input S;
	output wire [8:0] O;
	wire [8:0] coreir_commonlib_mux2x9_inst0_out;
	wire [17:0] coreir_commonlib_mux2x9_inst0_in_data;
	assign coreir_commonlib_mux2x9_inst0_in_data[9+:9] = I1;
	assign coreir_commonlib_mux2x9_inst0_in_data[0+:9] = I0;
	PEGEN_commonlib_muxn__N2__width9 coreir_commonlib_mux2x9_inst0(
		.in_data(coreir_commonlib_mux2x9_inst0_in_data),
		.in_sel(S),
		.out(coreir_commonlib_mux2x9_inst0_out)
	);
	assign O = coreir_commonlib_mux2x9_inst0_out;
endmodule
module PEGEN_Mux2xSInt16 (
	I0,
	I1,
	S,
	O
);
	input [15:0] I0;
	input [15:0] I1;
	input S;
	output wire [15:0] O;
	wire [15:0] coreir_commonlib_mux2x16_inst0_out;
	wire [31:0] coreir_commonlib_mux2x16_inst0_in_data;
	assign coreir_commonlib_mux2x16_inst0_in_data[16+:16] = I1;
	assign coreir_commonlib_mux2x16_inst0_in_data[0+:16] = I0;
	PEGEN_commonlib_muxn__N2__width16 coreir_commonlib_mux2x16_inst0(
		.in_data(coreir_commonlib_mux2x16_inst0_in_data),
		.in_sel(S),
		.out(coreir_commonlib_mux2x16_inst0_out)
	);
	assign O = coreir_commonlib_mux2x16_inst0_out;
endmodule
module PEGEN_Mux2xMagmaADTFPU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3 (
	I0,
	I1,
	S,
	O
);
	input [1:0] I0;
	input [1:0] I1;
	input S;
	output wire [1:0] O;
	wire [1:0] coreir_commonlib_mux2x2_inst0_out;
	wire [3:0] coreir_commonlib_mux2x2_inst0_in_data;
	assign coreir_commonlib_mux2x2_inst0_in_data[2+:2] = I1;
	assign coreir_commonlib_mux2x2_inst0_in_data[0+:2] = I0;
	PEGEN_commonlib_muxn__N2__width2 coreir_commonlib_mux2x2_inst0(
		.in_data(coreir_commonlib_mux2x2_inst0_in_data),
		.in_sel(S),
		.out(coreir_commonlib_mux2x2_inst0_out)
	);
	assign O = coreir_commonlib_mux2x2_inst0_out;
endmodule
module PEGEN_Mux2xMagmaADTFPCustom_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3 (
	I0,
	I1,
	S,
	O
);
	input [2:0] I0;
	input [2:0] I1;
	input S;
	output wire [2:0] O;
	wire [2:0] coreir_commonlib_mux2x3_inst0_out;
	wire [5:0] coreir_commonlib_mux2x3_inst0_in_data;
	assign coreir_commonlib_mux2x3_inst0_in_data[3+:3] = I1;
	assign coreir_commonlib_mux2x3_inst0_in_data[0+:3] = I0;
	PEGEN_commonlib_muxn__N2__width3 coreir_commonlib_mux2x3_inst0(
		.in_data(coreir_commonlib_mux2x3_inst0_in_data),
		.in_sel(S),
		.out(coreir_commonlib_mux2x3_inst0_out)
	);
	assign O = coreir_commonlib_mux2x3_inst0_out;
endmodule
module PEGEN_Mux2xMagmaADTALU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3 (
	I0,
	I1,
	S,
	O
);
	input [4:0] I0;
	input [4:0] I1;
	input S;
	output wire [4:0] O;
	wire [4:0] coreir_commonlib_mux2x5_inst0_out;
	wire [9:0] coreir_commonlib_mux2x5_inst0_in_data;
	assign coreir_commonlib_mux2x5_inst0_in_data[5+:5] = I1;
	assign coreir_commonlib_mux2x5_inst0_in_data[0+:5] = I0;
	PEGEN_commonlib_muxn__N2__width5 coreir_commonlib_mux2x5_inst0(
		.in_data(coreir_commonlib_mux2x5_inst0_in_data),
		.in_sel(S),
		.out(coreir_commonlib_mux2x5_inst0_out)
	);
	assign O = coreir_commonlib_mux2x5_inst0_out;
endmodule
module PEGEN_Mux2xBits8 (
	I0,
	I1,
	S,
	O
);
	input [7:0] I0;
	input [7:0] I1;
	input S;
	output wire [7:0] O;
	wire [7:0] coreir_commonlib_mux2x8_inst0_out;
	wire [15:0] coreir_commonlib_mux2x8_inst0_in_data;
	assign coreir_commonlib_mux2x8_inst0_in_data[8+:8] = I1;
	assign coreir_commonlib_mux2x8_inst0_in_data[0+:8] = I0;
	PEGEN_commonlib_muxn__N2__width8 coreir_commonlib_mux2x8_inst0(
		.in_data(coreir_commonlib_mux2x8_inst0_in_data),
		.in_sel(S),
		.out(coreir_commonlib_mux2x8_inst0_out)
	);
	assign O = coreir_commonlib_mux2x8_inst0_out;
endmodule
module PEGEN_Mux2xBits23 (
	I0,
	I1,
	S,
	O
);
	input [22:0] I0;
	input [22:0] I1;
	input S;
	output wire [22:0] O;
	wire [22:0] coreir_commonlib_mux2x23_inst0_out;
	wire [45:0] coreir_commonlib_mux2x23_inst0_in_data;
	assign coreir_commonlib_mux2x23_inst0_in_data[23+:23] = I1;
	assign coreir_commonlib_mux2x23_inst0_in_data[0+:23] = I0;
	PEGEN_commonlib_muxn__N2__width23 coreir_commonlib_mux2x23_inst0(
		.in_data(coreir_commonlib_mux2x23_inst0_in_data),
		.in_sel(S),
		.out(coreir_commonlib_mux2x23_inst0_out)
	);
	assign O = coreir_commonlib_mux2x23_inst0_out;
endmodule
module PEGEN_Mux2xBits16 (
	I0,
	I1,
	S,
	O
);
	input [15:0] I0;
	input [15:0] I1;
	input S;
	output wire [15:0] O;
	wire [15:0] coreir_commonlib_mux2x16_inst0_out;
	wire [31:0] coreir_commonlib_mux2x16_inst0_in_data;
	assign coreir_commonlib_mux2x16_inst0_in_data[16+:16] = I1;
	assign coreir_commonlib_mux2x16_inst0_in_data[0+:16] = I0;
	PEGEN_commonlib_muxn__N2__width16 coreir_commonlib_mux2x16_inst0(
		.in_data(coreir_commonlib_mux2x16_inst0_in_data),
		.in_sel(S),
		.out(coreir_commonlib_mux2x16_inst0_out)
	);
	assign O = coreir_commonlib_mux2x16_inst0_out;
endmodule
module PEGEN_Register (
	value,
	O,
	en,
	CLK,
	ASYNCRESET
);
	input [15:0] value;
	output wire [15:0] O;
	input en;
	input CLK;
	input ASYNCRESET;
	wire [15:0] enable_mux_O;
	wire [15:0] reg_PR16_inst0_out;
	PEGEN_Mux2xBits16 enable_mux(
		.I0(reg_PR16_inst0_out),
		.I1(value),
		.S(en),
		.O(enable_mux_O)
	);
	PEGEN_coreir_reg_arst #(
		.arst_posedge(1'b1),
		.clk_posedge(1'b1),
		.init(16'h0000),
		.width(16)
	) reg_PR16_inst0(
		.clk(CLK),
		.arst(ASYNCRESET),
		.in(enable_mux_O),
		.out(reg_PR16_inst0_out)
	);
	assign O = reg_PR16_inst0_out;
endmodule
module PEGEN_Mux2xBit (
	I0,
	I1,
	S,
	O
);
	input I0;
	input I1;
	input S;
	output wire O;
	wire [0:0] coreir_commonlib_mux2x1_inst0_out;
	wire [1:0] coreir_commonlib_mux2x1_inst0_in_data;
	assign coreir_commonlib_mux2x1_inst0_in_data[1+:1] = I1;
	assign coreir_commonlib_mux2x1_inst0_in_data[0+:1] = I0;
	PEGEN_commonlib_muxn__N2__width1 coreir_commonlib_mux2x1_inst0(
		.in_data(coreir_commonlib_mux2x1_inst0_in_data),
		.in_sel(S),
		.out(coreir_commonlib_mux2x1_inst0_out)
	);
	assign O = coreir_commonlib_mux2x1_inst0_out[0];
endmodule
module PEGEN_Register_unq1 (
	value,
	O,
	en,
	CLK,
	ASYNCRESET
);
	input value;
	output wire O;
	input en;
	input CLK;
	input ASYNCRESET;
	wire enable_mux_O;
	wire [0:0] reg_PR1_inst0_out;
	PEGEN_Mux2xBit enable_mux(
		.I0(reg_PR1_inst0_out[0]),
		.I1(value),
		.S(en),
		.O(enable_mux_O)
	);
	PEGEN_coreir_reg_arst #(
		.arst_posedge(1'b1),
		.clk_posedge(1'b1),
		.init(1'h0),
		.width(1)
	) reg_PR1_inst0(
		.clk(CLK),
		.arst(ASYNCRESET),
		.in(enable_mux_O),
		.out(reg_PR1_inst0_out)
	);
	assign O = reg_PR1_inst0_out[0];
endmodule
module PEGEN_RegisterMode_unq1 (
	mode,
	const_,
	value,
	clk_en,
	O0,
	O1,
	CLK,
	ASYNCRESET
);
	input [1:0] mode;
	input const_;
	input value;
	input clk_en;
	output wire O0;
	output wire O1;
	input CLK;
	input ASYNCRESET;
	wire Mux2xBit_inst0_O;
	wire Mux2xBit_inst1_O;
	wire Mux2xBit_inst2_O;
	wire Mux2xBit_inst3_O;
	wire Mux2xBit_inst4_O;
	wire Mux2xBit_inst5_O;
	wire Register_inst0_O;
	wire bit_const_0_None_out;
	wire [1:0] const_0_2_out;
	wire [1:0] const_2_2_out;
	wire [1:0] const_3_2_out;
	wire magma_Bits_2_eq_inst0_out;
	wire magma_Bits_2_eq_inst1_out;
	wire magma_Bits_2_eq_inst2_out;
	PEGEN_Mux2xBit Mux2xBit_inst0(
		.I0(value),
		.I1(value),
		.S(magma_Bits_2_eq_inst0_out),
		.O(Mux2xBit_inst0_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst1(
		.I0(bit_const_0_None_out),
		.I1(clk_en),
		.S(magma_Bits_2_eq_inst0_out),
		.O(Mux2xBit_inst1_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst2(
		.I0(Register_inst0_O),
		.I1(value),
		.S(magma_Bits_2_eq_inst2_out),
		.O(Mux2xBit_inst2_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst3(
		.I0(Register_inst0_O),
		.I1(Register_inst0_O),
		.S(magma_Bits_2_eq_inst2_out),
		.O(Mux2xBit_inst3_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst4(
		.I0(Mux2xBit_inst2_O),
		.I1(const_),
		.S(magma_Bits_2_eq_inst1_out),
		.O(Mux2xBit_inst4_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst5(
		.I0(Mux2xBit_inst3_O),
		.I1(Register_inst0_O),
		.S(magma_Bits_2_eq_inst1_out),
		.O(Mux2xBit_inst5_O)
	);
	PEGEN_Register_unq1 Register_inst0(
		.value(Mux2xBit_inst0_O),
		.O(Register_inst0_O),
		.en(Mux2xBit_inst1_O),
		.CLK(CLK),
		.ASYNCRESET(ASYNCRESET)
	);
	PEGEN_corebit_const #(.value(1'b0)) bit_const_0_None(.out(bit_const_0_None_out));
	PEGEN_coreir_const #(
		.value(2'h0),
		.width(2)
	) const_0_2(.out(const_0_2_out));
	PEGEN_coreir_const #(
		.value(2'h2),
		.width(2)
	) const_2_2(.out(const_2_2_out));
	PEGEN_coreir_const #(
		.value(2'h3),
		.width(2)
	) const_3_2(.out(const_3_2_out));
	PEGEN_coreir_eq #(.width(2)) magma_Bits_2_eq_inst0(
		.in0(mode),
		.in1(const_3_2_out),
		.out(magma_Bits_2_eq_inst0_out)
	);
	PEGEN_coreir_eq #(.width(2)) magma_Bits_2_eq_inst1(
		.in0(mode),
		.in1(const_0_2_out),
		.out(magma_Bits_2_eq_inst1_out)
	);
	PEGEN_coreir_eq #(.width(2)) magma_Bits_2_eq_inst2(
		.in0(mode),
		.in1(const_2_2_out),
		.out(magma_Bits_2_eq_inst2_out)
	);
	assign O0 = Mux2xBit_inst4_O;
	assign O1 = Mux2xBit_inst5_O;
endmodule
module PEGEN_RegisterMode (
	mode,
	const_,
	value,
	clk_en,
	O0,
	O1,
	CLK,
	ASYNCRESET
);
	input [1:0] mode;
	input [15:0] const_;
	input [15:0] value;
	input clk_en;
	output wire [15:0] O0;
	output wire [15:0] O1;
	input CLK;
	input ASYNCRESET;
	wire Mux2xBit_inst0_O;
	wire [15:0] Mux2xBits16_inst0_O;
	wire [15:0] Mux2xBits16_inst1_O;
	wire [15:0] Mux2xBits16_inst2_O;
	wire [15:0] Mux2xBits16_inst3_O;
	wire [15:0] Mux2xBits16_inst4_O;
	wire [15:0] Register_inst0_O;
	wire bit_const_0_None_out;
	wire [1:0] const_0_2_out;
	wire [1:0] const_2_2_out;
	wire [1:0] const_3_2_out;
	wire magma_Bits_2_eq_inst0_out;
	wire magma_Bits_2_eq_inst1_out;
	wire magma_Bits_2_eq_inst2_out;
	PEGEN_Mux2xBit Mux2xBit_inst0(
		.I0(bit_const_0_None_out),
		.I1(clk_en),
		.S(magma_Bits_2_eq_inst0_out),
		.O(Mux2xBit_inst0_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst0(
		.I0(value),
		.I1(value),
		.S(magma_Bits_2_eq_inst0_out),
		.O(Mux2xBits16_inst0_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst1(
		.I0(Register_inst0_O),
		.I1(value),
		.S(magma_Bits_2_eq_inst2_out),
		.O(Mux2xBits16_inst1_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst2(
		.I0(Register_inst0_O),
		.I1(Register_inst0_O),
		.S(magma_Bits_2_eq_inst2_out),
		.O(Mux2xBits16_inst2_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst3(
		.I0(Mux2xBits16_inst1_O),
		.I1(const_),
		.S(magma_Bits_2_eq_inst1_out),
		.O(Mux2xBits16_inst3_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst4(
		.I0(Mux2xBits16_inst2_O),
		.I1(Register_inst0_O),
		.S(magma_Bits_2_eq_inst1_out),
		.O(Mux2xBits16_inst4_O)
	);
	PEGEN_Register Register_inst0(
		.value(Mux2xBits16_inst0_O),
		.O(Register_inst0_O),
		.en(Mux2xBit_inst0_O),
		.CLK(CLK),
		.ASYNCRESET(ASYNCRESET)
	);
	PEGEN_corebit_const #(.value(1'b0)) bit_const_0_None(.out(bit_const_0_None_out));
	PEGEN_coreir_const #(
		.value(2'h0),
		.width(2)
	) const_0_2(.out(const_0_2_out));
	PEGEN_coreir_const #(
		.value(2'h2),
		.width(2)
	) const_2_2(.out(const_2_2_out));
	PEGEN_coreir_const #(
		.value(2'h3),
		.width(2)
	) const_3_2(.out(const_3_2_out));
	PEGEN_coreir_eq #(.width(2)) magma_Bits_2_eq_inst0(
		.in0(mode),
		.in1(const_3_2_out),
		.out(magma_Bits_2_eq_inst0_out)
	);
	PEGEN_coreir_eq #(.width(2)) magma_Bits_2_eq_inst1(
		.in0(mode),
		.in1(const_0_2_out),
		.out(magma_Bits_2_eq_inst1_out)
	);
	PEGEN_coreir_eq #(.width(2)) magma_Bits_2_eq_inst2(
		.in0(mode),
		.in1(const_2_2_out),
		.out(magma_Bits_2_eq_inst2_out)
	);
	assign O0 = Mux2xBits16_inst3_O;
	assign O1 = Mux2xBits16_inst4_O;
endmodule
module PEGEN_LUT (
	lut,
	bit0,
	bit1,
	bit2,
	O,
	CLK,
	ASYNCRESET
);
	input [7:0] lut;
	input bit0;
	input bit1;
	input bit2;
	output wire O;
	input CLK;
	input ASYNCRESET;
	wire bit_const_0_None_out;
	wire [7:0] const_1_8_out;
	wire [7:0] magma_Bits_8_and_inst0_out;
	wire [7:0] magma_Bits_8_lshr_inst0_out;
	PEGEN_corebit_const #(.value(1'b0)) bit_const_0_None(.out(bit_const_0_None_out));
	PEGEN_coreir_const #(
		.value(8'h01),
		.width(8)
	) const_1_8(.out(const_1_8_out));
	PEGEN_coreir_and #(.width(8)) magma_Bits_8_and_inst0(
		.in0(magma_Bits_8_lshr_inst0_out),
		.in1(const_1_8_out),
		.out(magma_Bits_8_and_inst0_out)
	);
	wire [7:0] magma_Bits_8_lshr_inst0_in1;
	assign magma_Bits_8_lshr_inst0_in1 = {bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit2, bit1, bit0};
	PEGEN_coreir_lshr #(.width(8)) magma_Bits_8_lshr_inst0(
		.in0(lut),
		.in1(magma_Bits_8_lshr_inst0_in1),
		.out(magma_Bits_8_lshr_inst0_out)
	);
	assign O = magma_Bits_8_and_inst0_out[0];
endmodule
module PEGEN_FPU (
	fpu_op,
	a,
	b,
	res,
	N,
	Z,
	CLK,
	ASYNCRESET
);
	input [1:0] fpu_op;
	input [15:0] a;
	input [15:0] b;
	output wire [15:0] res;
	output wire N;
	output wire Z;
	input CLK;
	input ASYNCRESET;
	wire Mux2xBit_inst0_O;
	wire Mux2xBit_inst1_O;
	wire [15:0] Mux2xBits16_inst0_O;
	wire [15:0] Mux2xBits16_inst1_O;
	wire [15:0] Op_inst0_O;
	wire [15:0] Op_inst1_O;
	wire bit_const_1_None_out;
	wire [1:0] const_0_2_out;
	wire [6:0] const_0_7_out;
	wire [7:0] const_0_8_out;
	wire [1:0] const_1_2_out;
	wire [7:0] const_255_8_out;
	wire [1:0] const_2_2_out;
	wire [15:0] const_32768_16_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bit_and_inst1_out;
	wire magma_Bit_and_inst2_out;
	wire magma_Bit_and_inst3_out;
	wire magma_Bit_and_inst4_out;
	wire magma_Bit_not_inst0_out;
	wire magma_Bit_or_inst0_out;
	wire magma_Bit_or_inst1_out;
	wire magma_Bit_or_inst2_out;
	wire magma_Bit_xor_inst0_out;
	wire [15:0] magma_Bits_16_xor_inst0_out;
	wire magma_Bits_2_eq_inst0_out;
	wire magma_Bits_2_eq_inst1_out;
	wire magma_Bits_2_eq_inst2_out;
	wire magma_Bits_2_eq_inst3_out;
	wire magma_Bits_2_eq_inst4_out;
	wire magma_Bits_2_eq_inst5_out;
	wire magma_Bits_7_eq_inst0_out;
	wire magma_Bits_7_eq_inst1_out;
	wire magma_Bits_7_eq_inst2_out;
	wire magma_Bits_8_eq_inst0_out;
	wire magma_Bits_8_eq_inst1_out;
	wire magma_Bits_8_eq_inst2_out;
	PEGEN_Mux2xBit Mux2xBit_inst0(
		.I0(magma_Bit_and_inst2_out),
		.I1(bit_const_1_None_out),
		.S(magma_Bit_and_inst4_out),
		.O(Mux2xBit_inst0_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst1(
		.I0(magma_Bit_and_inst2_out),
		.I1(Mux2xBit_inst0_O),
		.S(magma_Bits_2_eq_inst5_out),
		.O(Mux2xBit_inst1_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst0(
		.I0(b),
		.I1(magma_Bits_16_xor_inst0_out),
		.S(magma_Bit_or_inst0_out),
		.O(Mux2xBits16_inst0_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst1(
		.I0(Op_inst1_O),
		.I1(Op_inst0_O),
		.S(magma_Bit_or_inst2_out),
		.O(Mux2xBits16_inst1_O)
	);
	PEGEN_Op Op_inst0(
		.in0(a),
		.in1(Mux2xBits16_inst0_O),
		.O(Op_inst0_O),
		.CLK(CLK),
		.ASYNCRESET(ASYNCRESET)
	);
	PEGEN_Op_unq1 Op_inst1(
		.in0(a),
		.in1(Mux2xBits16_inst0_O),
		.O(Op_inst1_O),
		.CLK(CLK),
		.ASYNCRESET(ASYNCRESET)
	);
	PEGEN_corebit_const #(.value(1'b1)) bit_const_1_None(.out(bit_const_1_None_out));
	PEGEN_coreir_const #(
		.value(2'h0),
		.width(2)
	) const_0_2(.out(const_0_2_out));
	PEGEN_coreir_const #(
		.value(7'h00),
		.width(7)
	) const_0_7(.out(const_0_7_out));
	PEGEN_coreir_const #(
		.value(8'h00),
		.width(8)
	) const_0_8(.out(const_0_8_out));
	PEGEN_coreir_const #(
		.value(2'h1),
		.width(2)
	) const_1_2(.out(const_1_2_out));
	PEGEN_coreir_const #(
		.value(8'hff),
		.width(8)
	) const_255_8(.out(const_255_8_out));
	PEGEN_coreir_const #(
		.value(2'h2),
		.width(2)
	) const_2_2(.out(const_2_2_out));
	PEGEN_coreir_const #(
		.value(16'h8000),
		.width(16)
	) const_32768_16(.out(const_32768_16_out));
	PEGEN_corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(magma_Bits_7_eq_inst0_out),
		.out(magma_Bit_and_inst0_out)
	);
	PEGEN_corebit_and magma_Bit_and_inst1(
		.in0(magma_Bits_8_eq_inst1_out),
		.in1(magma_Bits_7_eq_inst1_out),
		.out(magma_Bit_and_inst1_out)
	);
	PEGEN_corebit_and magma_Bit_and_inst2(
		.in0(magma_Bits_8_eq_inst2_out),
		.in1(magma_Bits_7_eq_inst2_out),
		.out(magma_Bit_and_inst2_out)
	);
	PEGEN_corebit_and magma_Bit_and_inst3(
		.in0(magma_Bit_and_inst0_out),
		.in1(magma_Bit_and_inst1_out),
		.out(magma_Bit_and_inst3_out)
	);
	PEGEN_corebit_and magma_Bit_and_inst4(
		.in0(magma_Bit_and_inst3_out),
		.in1(magma_Bit_not_inst0_out),
		.out(magma_Bit_and_inst4_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst0(
		.in(magma_Bit_xor_inst0_out),
		.out(magma_Bit_not_inst0_out)
	);
	PEGEN_corebit_or magma_Bit_or_inst0(
		.in0(magma_Bits_2_eq_inst0_out),
		.in1(magma_Bits_2_eq_inst1_out),
		.out(magma_Bit_or_inst0_out)
	);
	PEGEN_corebit_or magma_Bit_or_inst1(
		.in0(magma_Bits_2_eq_inst2_out),
		.in1(magma_Bits_2_eq_inst3_out),
		.out(magma_Bit_or_inst1_out)
	);
	PEGEN_corebit_or magma_Bit_or_inst2(
		.in0(magma_Bit_or_inst1_out),
		.in1(magma_Bits_2_eq_inst4_out),
		.out(magma_Bit_or_inst2_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst0(
		.in0(a[15]),
		.in1(b[15]),
		.out(magma_Bit_xor_inst0_out)
	);
	PEGEN_coreir_xor #(.width(16)) magma_Bits_16_xor_inst0(
		.in0(b),
		.in1(const_32768_16_out),
		.out(magma_Bits_16_xor_inst0_out)
	);
	PEGEN_coreir_eq #(.width(2)) magma_Bits_2_eq_inst0(
		.in0(fpu_op),
		.in1(const_1_2_out),
		.out(magma_Bits_2_eq_inst0_out)
	);
	PEGEN_coreir_eq #(.width(2)) magma_Bits_2_eq_inst1(
		.in0(fpu_op),
		.in1(const_2_2_out),
		.out(magma_Bits_2_eq_inst1_out)
	);
	PEGEN_coreir_eq #(.width(2)) magma_Bits_2_eq_inst2(
		.in0(fpu_op),
		.in1(const_0_2_out),
		.out(magma_Bits_2_eq_inst2_out)
	);
	PEGEN_coreir_eq #(.width(2)) magma_Bits_2_eq_inst3(
		.in0(fpu_op),
		.in1(const_1_2_out),
		.out(magma_Bits_2_eq_inst3_out)
	);
	PEGEN_coreir_eq #(.width(2)) magma_Bits_2_eq_inst4(
		.in0(fpu_op),
		.in1(const_2_2_out),
		.out(magma_Bits_2_eq_inst4_out)
	);
	PEGEN_coreir_eq #(.width(2)) magma_Bits_2_eq_inst5(
		.in0(fpu_op),
		.in1(const_2_2_out),
		.out(magma_Bits_2_eq_inst5_out)
	);
	PEGEN_coreir_eq #(.width(7)) magma_Bits_7_eq_inst0(
		.in0(a[6:0]),
		.in1(const_0_7_out),
		.out(magma_Bits_7_eq_inst0_out)
	);
	PEGEN_coreir_eq #(.width(7)) magma_Bits_7_eq_inst1(
		.in0(b[6:0]),
		.in1(const_0_7_out),
		.out(magma_Bits_7_eq_inst1_out)
	);
	PEGEN_coreir_eq #(.width(7)) magma_Bits_7_eq_inst2(
		.in0(Mux2xBits16_inst1_O[6:0]),
		.in1(const_0_7_out),
		.out(magma_Bits_7_eq_inst2_out)
	);
	PEGEN_coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(a[14:7]),
		.in1(const_255_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	PEGEN_coreir_eq #(.width(8)) magma_Bits_8_eq_inst1(
		.in0(b[14:7]),
		.in1(const_255_8_out),
		.out(magma_Bits_8_eq_inst1_out)
	);
	PEGEN_coreir_eq #(.width(8)) magma_Bits_8_eq_inst2(
		.in0(Mux2xBits16_inst1_O[14:7]),
		.in1(const_0_8_out),
		.out(magma_Bits_8_eq_inst2_out)
	);
	assign res = Mux2xBits16_inst1_O;
	assign N = Mux2xBits16_inst1_O[15];
	assign Z = Mux2xBit_inst1_O;
endmodule
module PEGEN_FPCustom (
	op,
	signed_,
	a,
	b,
	res,
	res_p,
	V,
	CLK,
	ASYNCRESET
);
	input [2:0] op;
	input [0:0] signed_;
	input [15:0] a;
	input [15:0] b;
	output wire [15:0] res;
	output wire res_p;
	output wire V;
	input CLK;
	input ASYNCRESET;
	wire Mux2xBit_inst0_O;
	wire Mux2xBit_inst1_O;
	wire Mux2xBit_inst10_O;
	wire Mux2xBit_inst2_O;
	wire Mux2xBit_inst3_O;
	wire Mux2xBit_inst4_O;
	wire Mux2xBit_inst5_O;
	wire Mux2xBit_inst6_O;
	wire Mux2xBit_inst7_O;
	wire Mux2xBit_inst8_O;
	wire Mux2xBit_inst9_O;
	wire [15:0] Mux2xBits16_inst0_O;
	wire [15:0] Mux2xBits16_inst1_O;
	wire [15:0] Mux2xBits16_inst10_O;
	wire [15:0] Mux2xBits16_inst11_O;
	wire [15:0] Mux2xBits16_inst12_O;
	wire [15:0] Mux2xBits16_inst13_O;
	wire [15:0] Mux2xBits16_inst14_O;
	wire [15:0] Mux2xBits16_inst15_O;
	wire [15:0] Mux2xBits16_inst16_O;
	wire [15:0] Mux2xBits16_inst17_O;
	wire [15:0] Mux2xBits16_inst18_O;
	wire [15:0] Mux2xBits16_inst19_O;
	wire [15:0] Mux2xBits16_inst2_O;
	wire [15:0] Mux2xBits16_inst20_O;
	wire [15:0] Mux2xBits16_inst3_O;
	wire [15:0] Mux2xBits16_inst4_O;
	wire [15:0] Mux2xBits16_inst5_O;
	wire [15:0] Mux2xBits16_inst6_O;
	wire [15:0] Mux2xBits16_inst7_O;
	wire [15:0] Mux2xBits16_inst8_O;
	wire [15:0] Mux2xBits16_inst9_O;
	wire [22:0] Mux2xBits23_inst0_O;
	wire [7:0] Mux2xBits8_inst0_O;
	wire [7:0] Mux2xBits8_inst1_O;
	wire [7:0] Mux2xBits8_inst2_O;
	wire [7:0] Mux2xBits8_inst3_O;
	wire [7:0] Mux2xBits8_inst4_O;
	wire [7:0] Mux2xBits8_inst5_O;
	wire [15:0] Mux2xSInt16_inst0_O;
	wire [15:0] Mux2xSInt16_inst1_O;
	wire [15:0] Mux2xSInt16_inst10_O;
	wire [15:0] Mux2xSInt16_inst11_O;
	wire [15:0] Mux2xSInt16_inst12_O;
	wire [15:0] Mux2xSInt16_inst13_O;
	wire [15:0] Mux2xSInt16_inst14_O;
	wire [15:0] Mux2xSInt16_inst15_O;
	wire [15:0] Mux2xSInt16_inst16_O;
	wire [15:0] Mux2xSInt16_inst17_O;
	wire [15:0] Mux2xSInt16_inst18_O;
	wire [15:0] Mux2xSInt16_inst19_O;
	wire [15:0] Mux2xSInt16_inst2_O;
	wire [15:0] Mux2xSInt16_inst20_O;
	wire [15:0] Mux2xSInt16_inst21_O;
	wire [15:0] Mux2xSInt16_inst22_O;
	wire [15:0] Mux2xSInt16_inst23_O;
	wire [15:0] Mux2xSInt16_inst24_O;
	wire [15:0] Mux2xSInt16_inst25_O;
	wire [15:0] Mux2xSInt16_inst26_O;
	wire [15:0] Mux2xSInt16_inst27_O;
	wire [15:0] Mux2xSInt16_inst28_O;
	wire [15:0] Mux2xSInt16_inst29_O;
	wire [15:0] Mux2xSInt16_inst3_O;
	wire [15:0] Mux2xSInt16_inst30_O;
	wire [15:0] Mux2xSInt16_inst4_O;
	wire [15:0] Mux2xSInt16_inst5_O;
	wire [15:0] Mux2xSInt16_inst6_O;
	wire [15:0] Mux2xSInt16_inst7_O;
	wire [15:0] Mux2xSInt16_inst8_O;
	wire [15:0] Mux2xSInt16_inst9_O;
	wire [8:0] Mux2xSInt9_inst0_O;
	wire [8:0] Mux2xSInt9_inst1_O;
	wire [8:0] Mux2xSInt9_inst10_O;
	wire [8:0] Mux2xSInt9_inst11_O;
	wire [8:0] Mux2xSInt9_inst12_O;
	wire [8:0] Mux2xSInt9_inst2_O;
	wire [8:0] Mux2xSInt9_inst3_O;
	wire [8:0] Mux2xSInt9_inst4_O;
	wire [8:0] Mux2xSInt9_inst5_O;
	wire [8:0] Mux2xSInt9_inst6_O;
	wire [8:0] Mux2xSInt9_inst7_O;
	wire [8:0] Mux2xSInt9_inst8_O;
	wire [8:0] Mux2xSInt9_inst9_O;
	wire bit_const_0_None_out;
	wire bit_const_1_None_out;
	wire [15:0] const_0_16_out;
	wire [22:0] const_0_23_out;
	wire [2:0] const_0_3_out;
	wire [8:0] const_0_9_out;
	wire [15:0] const_10_16_out;
	wire [15:0] const_11_16_out;
	wire [15:0] const_127_16_out;
	wire [7:0] const_127_8_out;
	wire [8:0] const_127_9_out;
	wire [15:0] const_128_16_out;
	wire [15:0] const_12_16_out;
	wire [15:0] const_13_16_out;
	wire [7:0] const_142_8_out;
	wire [15:0] const_14_16_out;
	wire [15:0] const_15_16_out;
	wire [0:0] const_1_1_out;
	wire [15:0] const_1_16_out;
	wire [2:0] const_1_3_out;
	wire [8:0] const_255_9_out;
	wire [15:0] const_2_16_out;
	wire [2:0] const_2_3_out;
	wire [15:0] const_32512_16_out;
	wire [15:0] const_32640_16_out;
	wire [15:0] const_32768_16_out;
	wire [15:0] const_3_16_out;
	wire [2:0] const_3_3_out;
	wire [15:0] const_4_16_out;
	wire [2:0] const_4_3_out;
	wire [15:0] const_5_16_out;
	wire [2:0] const_5_3_out;
	wire [15:0] const_65409_16_out;
	wire [15:0] const_6_16_out;
	wire [2:0] const_6_3_out;
	wire [15:0] const_7_16_out;
	wire [22:0] const_7_23_out;
	wire [15:0] const_8_16_out;
	wire [15:0] const_9_16_out;
	wire magma_Bit_not_inst0_out;
	wire magma_Bit_not_inst1_out;
	wire magma_Bit_not_inst10_out;
	wire magma_Bit_not_inst11_out;
	wire magma_Bit_not_inst12_out;
	wire magma_Bit_not_inst13_out;
	wire magma_Bit_not_inst14_out;
	wire magma_Bit_not_inst15_out;
	wire magma_Bit_not_inst16_out;
	wire magma_Bit_not_inst17_out;
	wire magma_Bit_not_inst18_out;
	wire magma_Bit_not_inst19_out;
	wire magma_Bit_not_inst2_out;
	wire magma_Bit_not_inst20_out;
	wire magma_Bit_not_inst21_out;
	wire magma_Bit_not_inst22_out;
	wire magma_Bit_not_inst23_out;
	wire magma_Bit_not_inst24_out;
	wire magma_Bit_not_inst3_out;
	wire magma_Bit_not_inst4_out;
	wire magma_Bit_not_inst5_out;
	wire magma_Bit_not_inst6_out;
	wire magma_Bit_not_inst7_out;
	wire magma_Bit_not_inst8_out;
	wire magma_Bit_not_inst9_out;
	wire magma_Bit_xor_inst0_out;
	wire magma_Bit_xor_inst1_out;
	wire magma_Bit_xor_inst10_out;
	wire magma_Bit_xor_inst11_out;
	wire magma_Bit_xor_inst12_out;
	wire magma_Bit_xor_inst13_out;
	wire magma_Bit_xor_inst14_out;
	wire magma_Bit_xor_inst15_out;
	wire magma_Bit_xor_inst16_out;
	wire magma_Bit_xor_inst17_out;
	wire magma_Bit_xor_inst18_out;
	wire magma_Bit_xor_inst19_out;
	wire magma_Bit_xor_inst2_out;
	wire magma_Bit_xor_inst20_out;
	wire magma_Bit_xor_inst21_out;
	wire magma_Bit_xor_inst22_out;
	wire magma_Bit_xor_inst23_out;
	wire magma_Bit_xor_inst24_out;
	wire magma_Bit_xor_inst3_out;
	wire magma_Bit_xor_inst4_out;
	wire magma_Bit_xor_inst5_out;
	wire magma_Bit_xor_inst6_out;
	wire magma_Bit_xor_inst7_out;
	wire magma_Bit_xor_inst8_out;
	wire magma_Bit_xor_inst9_out;
	wire [15:0] magma_Bits_16_and_inst0_out;
	wire [15:0] magma_Bits_16_and_inst1_out;
	wire [15:0] magma_Bits_16_and_inst10_out;
	wire [15:0] magma_Bits_16_and_inst11_out;
	wire [15:0] magma_Bits_16_and_inst12_out;
	wire [15:0] magma_Bits_16_and_inst2_out;
	wire [15:0] magma_Bits_16_and_inst3_out;
	wire [15:0] magma_Bits_16_and_inst4_out;
	wire [15:0] magma_Bits_16_and_inst5_out;
	wire [15:0] magma_Bits_16_and_inst6_out;
	wire [15:0] magma_Bits_16_and_inst7_out;
	wire [15:0] magma_Bits_16_and_inst8_out;
	wire [15:0] magma_Bits_16_and_inst9_out;
	wire magma_Bits_16_eq_inst0_out;
	wire magma_Bits_16_eq_inst1_out;
	wire [15:0] magma_Bits_16_lshr_inst0_out;
	wire [15:0] magma_Bits_16_lshr_inst1_out;
	wire [15:0] magma_Bits_16_or_inst0_out;
	wire [15:0] magma_Bits_16_or_inst1_out;
	wire [15:0] magma_Bits_16_or_inst2_out;
	wire [15:0] magma_Bits_16_or_inst3_out;
	wire [15:0] magma_Bits_16_or_inst4_out;
	wire [15:0] magma_Bits_16_or_inst5_out;
	wire [15:0] magma_Bits_16_or_inst6_out;
	wire [15:0] magma_Bits_16_or_inst7_out;
	wire [15:0] magma_Bits_16_or_inst8_out;
	wire [15:0] magma_Bits_16_shl_inst0_out;
	wire [15:0] magma_Bits_16_shl_inst1_out;
	wire [15:0] magma_Bits_16_shl_inst2_out;
	wire [15:0] magma_Bits_16_shl_inst3_out;
	wire magma_Bits_1_eq_inst0_out;
	wire [22:0] magma_Bits_23_lshr_inst0_out;
	wire [22:0] magma_Bits_23_shl_inst0_out;
	wire magma_Bits_3_eq_inst0_out;
	wire magma_Bits_3_eq_inst1_out;
	wire magma_Bits_3_eq_inst2_out;
	wire magma_Bits_3_eq_inst3_out;
	wire magma_Bits_3_eq_inst4_out;
	wire magma_Bits_3_eq_inst5_out;
	wire magma_Bits_3_eq_inst6_out;
	wire magma_Bits_3_eq_inst7_out;
	wire [15:0] magma_SInt_16_add_inst0_out;
	wire [15:0] magma_SInt_16_and_inst0_out;
	wire [15:0] magma_SInt_16_neg_inst0_out;
	wire [15:0] magma_SInt_16_neg_inst1_out;
	wire [15:0] magma_SInt_16_neg_inst2_out;
	wire magma_SInt_16_sge_inst0_out;
	wire [15:0] magma_SInt_16_shl_inst0_out;
	wire [15:0] magma_SInt_16_sub_inst0_out;
	wire [15:0] magma_SInt_16_sub_inst1_out;
	wire [8:0] magma_SInt_9_neg_inst0_out;
	wire [8:0] magma_SInt_9_neg_inst1_out;
	wire magma_SInt_9_slt_inst0_out;
	wire magma_SInt_9_slt_inst1_out;
	wire magma_SInt_9_slt_inst2_out;
	wire [8:0] magma_SInt_9_sub_inst0_out;
	wire [8:0] magma_SInt_9_sub_inst1_out;
	wire [8:0] magma_SInt_9_sub_inst2_out;
	wire [7:0] magma_UInt_8_add_inst0_out;
	wire [7:0] magma_UInt_8_add_inst1_out;
	wire [7:0] magma_UInt_8_sub_inst0_out;
	wire magma_UInt_8_ugt_inst0_out;
	wire [8:0] magma_UInt_9_add_inst0_out;
	wire magma_UInt_9_ugt_inst0_out;
	PEGEN_Mux2xBit Mux2xBit_inst0(
		.I0(bit_const_0_None_out),
		.I1(bit_const_0_None_out),
		.S(magma_Bits_3_eq_inst7_out),
		.O(Mux2xBit_inst0_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst1(
		.I0(bit_const_0_None_out),
		.I1(magma_UInt_8_ugt_inst0_out),
		.S(magma_Bits_3_eq_inst6_out),
		.O(Mux2xBit_inst1_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst10(
		.I0(Mux2xBit_inst8_O),
		.I1(bit_const_0_None_out),
		.S(magma_Bits_3_eq_inst2_out),
		.O(Mux2xBit_inst10_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst2(
		.I0(Mux2xBit_inst0_O),
		.I1(bit_const_0_None_out),
		.S(magma_Bits_3_eq_inst6_out),
		.O(Mux2xBit_inst2_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst3(
		.I0(Mux2xBit_inst1_O),
		.I1(bit_const_0_None_out),
		.S(magma_Bits_3_eq_inst5_out),
		.O(Mux2xBit_inst3_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst4(
		.I0(Mux2xBit_inst2_O),
		.I1(bit_const_0_None_out),
		.S(magma_Bits_3_eq_inst5_out),
		.O(Mux2xBit_inst4_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst5(
		.I0(Mux2xBit_inst3_O),
		.I1(bit_const_0_None_out),
		.S(magma_Bits_3_eq_inst4_out),
		.O(Mux2xBit_inst5_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst6(
		.I0(Mux2xBit_inst4_O),
		.I1(bit_const_0_None_out),
		.S(magma_Bits_3_eq_inst4_out),
		.O(Mux2xBit_inst6_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst7(
		.I0(Mux2xBit_inst5_O),
		.I1(bit_const_0_None_out),
		.S(magma_Bits_3_eq_inst3_out),
		.O(Mux2xBit_inst7_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst8(
		.I0(Mux2xBit_inst6_O),
		.I1(magma_UInt_9_ugt_inst0_out),
		.S(magma_Bits_3_eq_inst3_out),
		.O(Mux2xBit_inst8_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst9(
		.I0(Mux2xBit_inst7_O),
		.I1(bit_const_0_None_out),
		.S(magma_Bits_3_eq_inst2_out),
		.O(Mux2xBit_inst9_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst0(
		.I0(const_0_16_out),
		.I1(const_32768_16_out),
		.S(magma_SInt_9_slt_inst0_out),
		.O(Mux2xBits16_inst0_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst1(
		.I0(const_0_16_out),
		.I1(magma_Bits_16_and_inst0_out),
		.S(magma_Bits_1_eq_inst0_out),
		.O(Mux2xBits16_inst1_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst10(
		.I0(magma_Bits_16_and_inst10_out),
		.I1(magma_Bits_16_and_inst8_out),
		.S(magma_Bits_3_eq_inst6_out),
		.O(Mux2xBits16_inst10_O)
	);
	wire [15:0] Mux2xBits16_inst11_I1;
	assign Mux2xBits16_inst11_I1 = {magma_Bits_23_lshr_inst0_out[15], magma_Bits_23_lshr_inst0_out[14], magma_Bits_23_lshr_inst0_out[13], magma_Bits_23_lshr_inst0_out[12], magma_Bits_23_lshr_inst0_out[11], magma_Bits_23_lshr_inst0_out[10], magma_Bits_23_lshr_inst0_out[9], magma_Bits_23_lshr_inst0_out[8], magma_Bits_23_lshr_inst0_out[7], magma_Bits_23_lshr_inst0_out[6], magma_Bits_23_lshr_inst0_out[5], magma_Bits_23_lshr_inst0_out[4], magma_Bits_23_lshr_inst0_out[3], magma_Bits_23_lshr_inst0_out[2], magma_Bits_23_lshr_inst0_out[1], magma_Bits_23_lshr_inst0_out[0]};
	PEGEN_Mux2xBits16 Mux2xBits16_inst11(
		.I0(magma_Bits_16_and_inst12_out),
		.I1(Mux2xBits16_inst11_I1),
		.S(magma_Bits_3_eq_inst6_out),
		.O(Mux2xBits16_inst11_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst12(
		.I0(Mux2xBits16_inst9_O),
		.I1(magma_Bits_16_or_inst1_out),
		.S(magma_Bits_3_eq_inst5_out),
		.O(Mux2xBits16_inst12_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst13(
		.I0(Mux2xBits16_inst8_O),
		.I1(magma_Bits_16_and_inst7_out),
		.S(magma_Bits_3_eq_inst4_out),
		.O(Mux2xBits16_inst13_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst14(
		.I0(Mux2xBits16_inst12_O),
		.I1(magma_Bits_16_or_inst6_out),
		.S(magma_Bits_3_eq_inst4_out),
		.O(Mux2xBits16_inst14_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst15(
		.I0(Mux2xBits16_inst10_O),
		.I1(magma_Bits_16_and_inst5_out),
		.S(magma_Bits_3_eq_inst4_out),
		.O(Mux2xBits16_inst15_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst16(
		.I0(magma_Bits_16_shl_inst2_out),
		.I1(magma_Bits_16_shl_inst1_out),
		.S(magma_Bits_3_eq_inst3_out),
		.O(Mux2xBits16_inst16_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst17(
		.I0(Mux2xBits16_inst14_O),
		.I1(magma_Bits_16_or_inst3_out),
		.S(magma_Bits_3_eq_inst3_out),
		.O(Mux2xBits16_inst17_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst18(
		.I0(Mux2xBits16_inst3_O),
		.I1(magma_Bits_16_and_inst3_out),
		.S(magma_Bits_3_eq_inst3_out),
		.O(Mux2xBits16_inst18_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst19(
		.I0(Mux2xBits16_inst17_O),
		.I1(magma_Bits_16_and_inst2_out),
		.S(magma_Bits_3_eq_inst2_out),
		.O(Mux2xBits16_inst19_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst2(
		.I0(a),
		.I1(magma_SInt_16_neg_inst0_out),
		.S(magma_Bit_not_inst8_out),
		.O(Mux2xBits16_inst2_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst20(
		.I0(Mux2xBits16_inst18_O),
		.I1(Mux2xBits16_inst3_O),
		.S(magma_Bits_3_eq_inst2_out),
		.O(Mux2xBits16_inst20_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst3(
		.I0(Mux2xBits16_inst1_O),
		.I1(Mux2xBits16_inst0_O),
		.S(magma_Bits_3_eq_inst0_out),
		.O(Mux2xBits16_inst3_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst4(
		.I0(const_0_16_out),
		.I1(magma_SInt_16_and_inst0_out),
		.S(magma_SInt_16_sge_inst0_out),
		.O(Mux2xBits16_inst4_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst5(
		.I0(Mux2xBits16_inst4_O),
		.I1(magma_Bits_16_lshr_inst0_out),
		.S(magma_Bits_3_eq_inst1_out),
		.O(Mux2xBits16_inst5_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst6(
		.I0(magma_Bits_16_shl_inst3_out),
		.I1(magma_Bits_16_lshr_inst1_out),
		.S(magma_SInt_9_slt_inst2_out),
		.O(Mux2xBits16_inst6_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst7(
		.I0(magma_Bits_16_or_inst1_out),
		.I1(Mux2xSInt16_inst29_O),
		.S(magma_Bits_3_eq_inst7_out),
		.O(Mux2xBits16_inst7_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst8(
		.I0(magma_Bits_16_or_inst8_out),
		.I1(magma_Bits_16_or_inst7_out),
		.S(magma_Bits_3_eq_inst6_out),
		.O(Mux2xBits16_inst8_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst9(
		.I0(Mux2xBits16_inst7_O),
		.I1(Mux2xSInt16_inst28_O),
		.S(magma_Bits_3_eq_inst6_out),
		.O(Mux2xBits16_inst9_O)
	);
	PEGEN_Mux2xBits23 Mux2xBits23_inst0(
		.I0(magma_Bits_23_shl_inst0_out),
		.I1(const_0_23_out),
		.S(magma_SInt_9_slt_inst1_out),
		.O(Mux2xBits23_inst0_O)
	);
	wire [7:0] Mux2xBits8_inst0_I0;
	assign Mux2xBits8_inst0_I0 = {a[14], a[13], a[12], a[11], a[10], a[9], a[8], a[7]};
	wire [7:0] Mux2xBits8_inst0_I1;
	assign Mux2xBits8_inst0_I1 = {a[14], a[13], a[12], a[11], a[10], a[9], a[8], a[7]};
	PEGEN_Mux2xBits8 Mux2xBits8_inst0(
		.I0(Mux2xBits8_inst0_I0),
		.I1(Mux2xBits8_inst0_I1),
		.S(magma_Bits_3_eq_inst7_out),
		.O(Mux2xBits8_inst0_O)
	);
	wire [7:0] Mux2xBits8_inst1_I1;
	assign Mux2xBits8_inst1_I1 = {a[14], a[13], a[12], a[11], a[10], a[9], a[8], a[7]};
	PEGEN_Mux2xBits8 Mux2xBits8_inst1(
		.I0(Mux2xBits8_inst0_O),
		.I1(Mux2xBits8_inst1_I1),
		.S(magma_Bits_3_eq_inst6_out),
		.O(Mux2xBits8_inst1_O)
	);
	wire [7:0] Mux2xBits8_inst2_I1;
	assign Mux2xBits8_inst2_I1 = {a[14], a[13], a[12], a[11], a[10], a[9], a[8], a[7]};
	PEGEN_Mux2xBits8 Mux2xBits8_inst2(
		.I0(Mux2xBits8_inst1_O),
		.I1(Mux2xBits8_inst2_I1),
		.S(magma_Bits_3_eq_inst5_out),
		.O(Mux2xBits8_inst2_O)
	);
	wire [7:0] Mux2xBits8_inst3_I1;
	assign Mux2xBits8_inst3_I1 = {a[14], a[13], a[12], a[11], a[10], a[9], a[8], a[7]};
	PEGEN_Mux2xBits8 Mux2xBits8_inst3(
		.I0(Mux2xBits8_inst2_O),
		.I1(Mux2xBits8_inst3_I1),
		.S(magma_Bits_3_eq_inst4_out),
		.O(Mux2xBits8_inst3_O)
	);
	wire [7:0] Mux2xBits8_inst4_I1;
	assign Mux2xBits8_inst4_I1 = {a[14], a[13], a[12], a[11], a[10], a[9], a[8], a[7]};
	PEGEN_Mux2xBits8 Mux2xBits8_inst4(
		.I0(Mux2xBits8_inst3_O),
		.I1(Mux2xBits8_inst4_I1),
		.S(magma_Bits_3_eq_inst3_out),
		.O(Mux2xBits8_inst4_O)
	);
	wire [7:0] Mux2xBits8_inst5_I1;
	assign Mux2xBits8_inst5_I1 = {a[14], a[13], a[12], a[11], a[10], a[9], a[8], a[7]};
	PEGEN_Mux2xBits8 Mux2xBits8_inst5(
		.I0(Mux2xBits8_inst4_O),
		.I1(Mux2xBits8_inst5_I1),
		.S(magma_Bits_3_eq_inst2_out),
		.O(Mux2xBits8_inst5_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst0(
		.I0(const_65409_16_out),
		.I1(const_0_16_out),
		.S(magma_Bit_not_inst0_out),
		.O(Mux2xSInt16_inst0_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst1(
		.I0(Mux2xSInt16_inst0_O),
		.I1(const_1_16_out),
		.S(magma_Bit_not_inst1_out),
		.O(Mux2xSInt16_inst1_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst10(
		.I0(Mux2xSInt16_inst9_O),
		.I1(const_2_16_out),
		.S(magma_Bit_not_inst11_out),
		.O(Mux2xSInt16_inst10_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst11(
		.I0(Mux2xSInt16_inst10_O),
		.I1(const_3_16_out),
		.S(magma_Bit_not_inst12_out),
		.O(Mux2xSInt16_inst11_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst12(
		.I0(Mux2xSInt16_inst11_O),
		.I1(const_4_16_out),
		.S(magma_Bit_not_inst13_out),
		.O(Mux2xSInt16_inst12_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst13(
		.I0(Mux2xSInt16_inst12_O),
		.I1(const_5_16_out),
		.S(magma_Bit_not_inst14_out),
		.O(Mux2xSInt16_inst13_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst14(
		.I0(Mux2xSInt16_inst13_O),
		.I1(const_6_16_out),
		.S(magma_Bit_not_inst15_out),
		.O(Mux2xSInt16_inst14_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst15(
		.I0(Mux2xSInt16_inst14_O),
		.I1(const_7_16_out),
		.S(magma_Bit_not_inst16_out),
		.O(Mux2xSInt16_inst15_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst16(
		.I0(Mux2xSInt16_inst15_O),
		.I1(const_8_16_out),
		.S(magma_Bit_not_inst17_out),
		.O(Mux2xSInt16_inst16_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst17(
		.I0(Mux2xSInt16_inst16_O),
		.I1(const_9_16_out),
		.S(magma_Bit_not_inst18_out),
		.O(Mux2xSInt16_inst17_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst18(
		.I0(Mux2xSInt16_inst17_O),
		.I1(const_10_16_out),
		.S(magma_Bit_not_inst19_out),
		.O(Mux2xSInt16_inst18_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst19(
		.I0(Mux2xSInt16_inst18_O),
		.I1(const_11_16_out),
		.S(magma_Bit_not_inst20_out),
		.O(Mux2xSInt16_inst19_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst2(
		.I0(Mux2xSInt16_inst1_O),
		.I1(const_2_16_out),
		.S(magma_Bit_not_inst2_out),
		.O(Mux2xSInt16_inst2_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst20(
		.I0(Mux2xSInt16_inst19_O),
		.I1(const_12_16_out),
		.S(magma_Bit_not_inst21_out),
		.O(Mux2xSInt16_inst20_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst21(
		.I0(Mux2xSInt16_inst20_O),
		.I1(const_13_16_out),
		.S(magma_Bit_not_inst22_out),
		.O(Mux2xSInt16_inst21_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst22(
		.I0(Mux2xSInt16_inst21_O),
		.I1(const_14_16_out),
		.S(magma_Bit_not_inst23_out),
		.O(Mux2xSInt16_inst22_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst23(
		.I0(Mux2xSInt16_inst22_O),
		.I1(const_15_16_out),
		.S(magma_Bit_not_inst24_out),
		.O(Mux2xSInt16_inst23_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst24(
		.I0(const_32512_16_out),
		.I1(const_127_16_out),
		.S(magma_Bits_3_eq_inst0_out),
		.O(Mux2xSInt16_inst24_O)
	);
	wire [15:0] Mux2xSInt16_inst25_I1;
	assign Mux2xSInt16_inst25_I1 = {Mux2xSInt9_inst0_O[7], Mux2xSInt9_inst0_O[7], Mux2xSInt9_inst0_O[7], Mux2xSInt9_inst0_O[7], Mux2xSInt9_inst0_O[7], Mux2xSInt9_inst0_O[7], Mux2xSInt9_inst0_O[7], Mux2xSInt9_inst0_O[7], Mux2xSInt9_inst0_O[7], Mux2xSInt9_inst0_O[6], Mux2xSInt9_inst0_O[5], Mux2xSInt9_inst0_O[4], Mux2xSInt9_inst0_O[3], Mux2xSInt9_inst0_O[2], Mux2xSInt9_inst0_O[1], Mux2xSInt9_inst0_O[0]};
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst25(
		.I0(Mux2xBits16_inst2_O),
		.I1(Mux2xSInt16_inst25_I1),
		.S(magma_Bits_3_eq_inst0_out),
		.O(Mux2xSInt16_inst25_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst26(
		.I0(magma_SInt_16_sub_inst1_out),
		.I1(magma_SInt_16_sub_inst0_out),
		.S(magma_Bits_3_eq_inst0_out),
		.O(Mux2xSInt16_inst26_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst27(
		.I0(Mux2xSInt16_inst23_O),
		.I1(Mux2xSInt16_inst7_O),
		.S(magma_Bits_3_eq_inst0_out),
		.O(Mux2xSInt16_inst27_O)
	);
	wire [15:0] Mux2xSInt16_inst28_I0;
	assign Mux2xSInt16_inst28_I0 = {magma_Bits_23_lshr_inst0_out[15], magma_Bits_23_lshr_inst0_out[14], magma_Bits_23_lshr_inst0_out[13], magma_Bits_23_lshr_inst0_out[12], magma_Bits_23_lshr_inst0_out[11], magma_Bits_23_lshr_inst0_out[10], magma_Bits_23_lshr_inst0_out[9], magma_Bits_23_lshr_inst0_out[8], magma_Bits_23_lshr_inst0_out[7], magma_Bits_23_lshr_inst0_out[6], magma_Bits_23_lshr_inst0_out[5], magma_Bits_23_lshr_inst0_out[4], magma_Bits_23_lshr_inst0_out[3], magma_Bits_23_lshr_inst0_out[2], magma_Bits_23_lshr_inst0_out[1], magma_Bits_23_lshr_inst0_out[0]};
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst28(
		.I0(Mux2xSInt16_inst28_I0),
		.I1(magma_SInt_16_neg_inst1_out),
		.S(magma_Bits_16_eq_inst0_out),
		.O(Mux2xSInt16_inst28_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst29(
		.I0(magma_Bits_16_and_inst12_out),
		.I1(magma_SInt_16_neg_inst2_out),
		.S(magma_Bits_16_eq_inst1_out),
		.O(Mux2xSInt16_inst29_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst3(
		.I0(Mux2xSInt16_inst2_O),
		.I1(const_3_16_out),
		.S(magma_Bit_not_inst3_out),
		.O(Mux2xSInt16_inst3_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst30(
		.I0(Mux2xSInt16_inst29_O),
		.I1(Mux2xSInt16_inst28_O),
		.S(magma_Bits_3_eq_inst6_out),
		.O(Mux2xSInt16_inst30_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst4(
		.I0(Mux2xSInt16_inst3_O),
		.I1(const_4_16_out),
		.S(magma_Bit_not_inst4_out),
		.O(Mux2xSInt16_inst4_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst5(
		.I0(Mux2xSInt16_inst4_O),
		.I1(const_5_16_out),
		.S(magma_Bit_not_inst5_out),
		.O(Mux2xSInt16_inst5_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst6(
		.I0(Mux2xSInt16_inst5_O),
		.I1(const_6_16_out),
		.S(magma_Bit_not_inst6_out),
		.O(Mux2xSInt16_inst6_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst7(
		.I0(Mux2xSInt16_inst6_O),
		.I1(const_7_16_out),
		.S(magma_Bit_not_inst7_out),
		.O(Mux2xSInt16_inst7_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst8(
		.I0(const_65409_16_out),
		.I1(const_0_16_out),
		.S(magma_Bit_not_inst9_out),
		.O(Mux2xSInt16_inst8_O)
	);
	PEGEN_Mux2xSInt16 Mux2xSInt16_inst9(
		.I0(Mux2xSInt16_inst8_O),
		.I1(const_1_16_out),
		.S(magma_Bit_not_inst10_out),
		.O(Mux2xSInt16_inst9_O)
	);
	PEGEN_Mux2xSInt9 Mux2xSInt9_inst0(
		.I0(magma_SInt_9_sub_inst0_out),
		.I1(magma_SInt_9_neg_inst0_out),
		.S(magma_SInt_9_slt_inst0_out),
		.O(Mux2xSInt9_inst0_O)
	);
	wire [8:0] Mux2xSInt9_inst1_I0;
	assign Mux2xSInt9_inst1_I0 = {bit_const_0_None_out, a[14], a[13], a[12], a[11], a[10], a[9], a[8], a[7]};
	wire [8:0] Mux2xSInt9_inst1_I1;
	assign Mux2xSInt9_inst1_I1 = {bit_const_0_None_out, a[14], a[13], a[12], a[11], a[10], a[9], a[8], a[7]};
	PEGEN_Mux2xSInt9 Mux2xSInt9_inst1(
		.I0(Mux2xSInt9_inst1_I0),
		.I1(Mux2xSInt9_inst1_I1),
		.S(magma_Bits_3_eq_inst7_out),
		.O(Mux2xSInt9_inst1_O)
	);
	PEGEN_Mux2xSInt9 Mux2xSInt9_inst10(
		.I0(Mux2xSInt9_inst8_O),
		.I1(magma_SInt_9_sub_inst0_out),
		.S(magma_Bits_3_eq_inst3_out),
		.O(Mux2xSInt9_inst10_O)
	);
	wire [8:0] Mux2xSInt9_inst11_I1;
	assign Mux2xSInt9_inst11_I1 = {bit_const_0_None_out, a[14], a[13], a[12], a[11], a[10], a[9], a[8], a[7]};
	PEGEN_Mux2xSInt9 Mux2xSInt9_inst11(
		.I0(Mux2xSInt9_inst9_O),
		.I1(Mux2xSInt9_inst11_I1),
		.S(magma_Bits_3_eq_inst2_out),
		.O(Mux2xSInt9_inst11_O)
	);
	PEGEN_Mux2xSInt9 Mux2xSInt9_inst12(
		.I0(Mux2xSInt9_inst10_O),
		.I1(magma_SInt_9_sub_inst0_out),
		.S(magma_Bits_3_eq_inst2_out),
		.O(Mux2xSInt9_inst12_O)
	);
	PEGEN_Mux2xSInt9 Mux2xSInt9_inst2(
		.I0(magma_SInt_9_sub_inst0_out),
		.I1(magma_SInt_9_sub_inst2_out),
		.S(magma_Bits_3_eq_inst7_out),
		.O(Mux2xSInt9_inst2_O)
	);
	wire [8:0] Mux2xSInt9_inst3_I1;
	assign Mux2xSInt9_inst3_I1 = {bit_const_0_None_out, a[14], a[13], a[12], a[11], a[10], a[9], a[8], a[7]};
	PEGEN_Mux2xSInt9 Mux2xSInt9_inst3(
		.I0(Mux2xSInt9_inst1_O),
		.I1(Mux2xSInt9_inst3_I1),
		.S(magma_Bits_3_eq_inst6_out),
		.O(Mux2xSInt9_inst3_O)
	);
	PEGEN_Mux2xSInt9 Mux2xSInt9_inst4(
		.I0(Mux2xSInt9_inst2_O),
		.I1(magma_SInt_9_sub_inst1_out),
		.S(magma_Bits_3_eq_inst6_out),
		.O(Mux2xSInt9_inst4_O)
	);
	wire [8:0] Mux2xSInt9_inst5_I1;
	assign Mux2xSInt9_inst5_I1 = {bit_const_0_None_out, a[14], a[13], a[12], a[11], a[10], a[9], a[8], a[7]};
	PEGEN_Mux2xSInt9 Mux2xSInt9_inst5(
		.I0(Mux2xSInt9_inst3_O),
		.I1(Mux2xSInt9_inst5_I1),
		.S(magma_Bits_3_eq_inst5_out),
		.O(Mux2xSInt9_inst5_O)
	);
	PEGEN_Mux2xSInt9 Mux2xSInt9_inst6(
		.I0(Mux2xSInt9_inst4_O),
		.I1(magma_SInt_9_sub_inst0_out),
		.S(magma_Bits_3_eq_inst5_out),
		.O(Mux2xSInt9_inst6_O)
	);
	wire [8:0] Mux2xSInt9_inst7_I1;
	assign Mux2xSInt9_inst7_I1 = {bit_const_0_None_out, a[14], a[13], a[12], a[11], a[10], a[9], a[8], a[7]};
	PEGEN_Mux2xSInt9 Mux2xSInt9_inst7(
		.I0(Mux2xSInt9_inst5_O),
		.I1(Mux2xSInt9_inst7_I1),
		.S(magma_Bits_3_eq_inst4_out),
		.O(Mux2xSInt9_inst7_O)
	);
	PEGEN_Mux2xSInt9 Mux2xSInt9_inst8(
		.I0(Mux2xSInt9_inst6_O),
		.I1(magma_SInt_9_sub_inst0_out),
		.S(magma_Bits_3_eq_inst4_out),
		.O(Mux2xSInt9_inst8_O)
	);
	wire [8:0] Mux2xSInt9_inst9_I1;
	assign Mux2xSInt9_inst9_I1 = {bit_const_0_None_out, a[14], a[13], a[12], a[11], a[10], a[9], a[8], a[7]};
	PEGEN_Mux2xSInt9 Mux2xSInt9_inst9(
		.I0(Mux2xSInt9_inst7_O),
		.I1(Mux2xSInt9_inst9_I1),
		.S(magma_Bits_3_eq_inst3_out),
		.O(Mux2xSInt9_inst9_O)
	);
	PEGEN_corebit_const #(.value(1'b0)) bit_const_0_None(.out(bit_const_0_None_out));
	PEGEN_corebit_const #(.value(1'b1)) bit_const_1_None(.out(bit_const_1_None_out));
	PEGEN_coreir_const #(
		.value(16'h0000),
		.width(16)
	) const_0_16(.out(const_0_16_out));
	PEGEN_coreir_const #(
		.value(23'h000000),
		.width(23)
	) const_0_23(.out(const_0_23_out));
	PEGEN_coreir_const #(
		.value(3'h0),
		.width(3)
	) const_0_3(.out(const_0_3_out));
	PEGEN_coreir_const #(
		.value(9'h000),
		.width(9)
	) const_0_9(.out(const_0_9_out));
	PEGEN_coreir_const #(
		.value(16'h000a),
		.width(16)
	) const_10_16(.out(const_10_16_out));
	PEGEN_coreir_const #(
		.value(16'h000b),
		.width(16)
	) const_11_16(.out(const_11_16_out));
	PEGEN_coreir_const #(
		.value(16'h007f),
		.width(16)
	) const_127_16(.out(const_127_16_out));
	PEGEN_coreir_const #(
		.value(8'h7f),
		.width(8)
	) const_127_8(.out(const_127_8_out));
	PEGEN_coreir_const #(
		.value(9'h07f),
		.width(9)
	) const_127_9(.out(const_127_9_out));
	PEGEN_coreir_const #(
		.value(16'h0080),
		.width(16)
	) const_128_16(.out(const_128_16_out));
	PEGEN_coreir_const #(
		.value(16'h000c),
		.width(16)
	) const_12_16(.out(const_12_16_out));
	PEGEN_coreir_const #(
		.value(16'h000d),
		.width(16)
	) const_13_16(.out(const_13_16_out));
	PEGEN_coreir_const #(
		.value(8'h8e),
		.width(8)
	) const_142_8(.out(const_142_8_out));
	PEGEN_coreir_const #(
		.value(16'h000e),
		.width(16)
	) const_14_16(.out(const_14_16_out));
	PEGEN_coreir_const #(
		.value(16'h000f),
		.width(16)
	) const_15_16(.out(const_15_16_out));
	PEGEN_coreir_const #(
		.value(1'h1),
		.width(1)
	) const_1_1(.out(const_1_1_out));
	PEGEN_coreir_const #(
		.value(16'h0001),
		.width(16)
	) const_1_16(.out(const_1_16_out));
	PEGEN_coreir_const #(
		.value(3'h1),
		.width(3)
	) const_1_3(.out(const_1_3_out));
	PEGEN_coreir_const #(
		.value(9'h0ff),
		.width(9)
	) const_255_9(.out(const_255_9_out));
	PEGEN_coreir_const #(
		.value(16'h0002),
		.width(16)
	) const_2_16(.out(const_2_16_out));
	PEGEN_coreir_const #(
		.value(3'h2),
		.width(3)
	) const_2_3(.out(const_2_3_out));
	PEGEN_coreir_const #(
		.value(16'h7f00),
		.width(16)
	) const_32512_16(.out(const_32512_16_out));
	PEGEN_coreir_const #(
		.value(16'h7f80),
		.width(16)
	) const_32640_16(.out(const_32640_16_out));
	PEGEN_coreir_const #(
		.value(16'h8000),
		.width(16)
	) const_32768_16(.out(const_32768_16_out));
	PEGEN_coreir_const #(
		.value(16'h0003),
		.width(16)
	) const_3_16(.out(const_3_16_out));
	PEGEN_coreir_const #(
		.value(3'h3),
		.width(3)
	) const_3_3(.out(const_3_3_out));
	PEGEN_coreir_const #(
		.value(16'h0004),
		.width(16)
	) const_4_16(.out(const_4_16_out));
	PEGEN_coreir_const #(
		.value(3'h4),
		.width(3)
	) const_4_3(.out(const_4_3_out));
	PEGEN_coreir_const #(
		.value(16'h0005),
		.width(16)
	) const_5_16(.out(const_5_16_out));
	PEGEN_coreir_const #(
		.value(3'h5),
		.width(3)
	) const_5_3(.out(const_5_3_out));
	PEGEN_coreir_const #(
		.value(16'hff81),
		.width(16)
	) const_65409_16(.out(const_65409_16_out));
	PEGEN_coreir_const #(
		.value(16'h0006),
		.width(16)
	) const_6_16(.out(const_6_16_out));
	PEGEN_coreir_const #(
		.value(3'h6),
		.width(3)
	) const_6_3(.out(const_6_3_out));
	PEGEN_coreir_const #(
		.value(16'h0007),
		.width(16)
	) const_7_16(.out(const_7_16_out));
	PEGEN_coreir_const #(
		.value(23'h000007),
		.width(23)
	) const_7_23(.out(const_7_23_out));
	PEGEN_coreir_const #(
		.value(16'h0008),
		.width(16)
	) const_8_16(.out(const_8_16_out));
	PEGEN_coreir_const #(
		.value(16'h0009),
		.width(16)
	) const_9_16(.out(const_9_16_out));
	PEGEN_corebit_not magma_Bit_not_inst0(
		.in(magma_Bit_xor_inst0_out),
		.out(magma_Bit_not_inst0_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst1(
		.in(magma_Bit_xor_inst1_out),
		.out(magma_Bit_not_inst1_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst10(
		.in(magma_Bit_xor_inst10_out),
		.out(magma_Bit_not_inst10_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst11(
		.in(magma_Bit_xor_inst11_out),
		.out(magma_Bit_not_inst11_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst12(
		.in(magma_Bit_xor_inst12_out),
		.out(magma_Bit_not_inst12_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst13(
		.in(magma_Bit_xor_inst13_out),
		.out(magma_Bit_not_inst13_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst14(
		.in(magma_Bit_xor_inst14_out),
		.out(magma_Bit_not_inst14_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst15(
		.in(magma_Bit_xor_inst15_out),
		.out(magma_Bit_not_inst15_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst16(
		.in(magma_Bit_xor_inst16_out),
		.out(magma_Bit_not_inst16_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst17(
		.in(magma_Bit_xor_inst17_out),
		.out(magma_Bit_not_inst17_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst18(
		.in(magma_Bit_xor_inst18_out),
		.out(magma_Bit_not_inst18_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst19(
		.in(magma_Bit_xor_inst19_out),
		.out(magma_Bit_not_inst19_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst2(
		.in(magma_Bit_xor_inst2_out),
		.out(magma_Bit_not_inst2_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst20(
		.in(magma_Bit_xor_inst20_out),
		.out(magma_Bit_not_inst20_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst21(
		.in(magma_Bit_xor_inst21_out),
		.out(magma_Bit_not_inst21_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst22(
		.in(magma_Bit_xor_inst22_out),
		.out(magma_Bit_not_inst22_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst23(
		.in(magma_Bit_xor_inst23_out),
		.out(magma_Bit_not_inst23_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst24(
		.in(magma_Bit_xor_inst24_out),
		.out(magma_Bit_not_inst24_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst3(
		.in(magma_Bit_xor_inst3_out),
		.out(magma_Bit_not_inst3_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst4(
		.in(magma_Bit_xor_inst4_out),
		.out(magma_Bit_not_inst4_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst5(
		.in(magma_Bit_xor_inst5_out),
		.out(magma_Bit_not_inst5_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst6(
		.in(magma_Bit_xor_inst6_out),
		.out(magma_Bit_not_inst6_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst7(
		.in(magma_Bit_xor_inst7_out),
		.out(magma_Bit_not_inst7_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst8(
		.in(magma_Bit_xor_inst8_out),
		.out(magma_Bit_not_inst8_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst9(
		.in(magma_Bit_xor_inst9_out),
		.out(magma_Bit_not_inst9_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst0(
		.in0(Mux2xSInt9_inst0_O[0]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst0_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst1(
		.in0(Mux2xSInt9_inst0_O[1]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst1_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst10(
		.in0(Mux2xBits16_inst2_O[1]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst10_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst11(
		.in0(Mux2xBits16_inst2_O[2]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst11_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst12(
		.in0(Mux2xBits16_inst2_O[3]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst12_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst13(
		.in0(Mux2xBits16_inst2_O[4]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst13_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst14(
		.in0(Mux2xBits16_inst2_O[5]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst14_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst15(
		.in0(Mux2xBits16_inst2_O[6]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst15_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst16(
		.in0(Mux2xBits16_inst2_O[7]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst16_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst17(
		.in0(Mux2xBits16_inst2_O[8]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst17_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst18(
		.in0(Mux2xBits16_inst2_O[9]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst18_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst19(
		.in0(Mux2xBits16_inst2_O[10]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst19_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst2(
		.in0(Mux2xSInt9_inst0_O[2]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst2_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst20(
		.in0(Mux2xBits16_inst2_O[11]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst20_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst21(
		.in0(Mux2xBits16_inst2_O[12]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst21_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst22(
		.in0(Mux2xBits16_inst2_O[13]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst22_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst23(
		.in0(Mux2xBits16_inst2_O[14]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst23_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst24(
		.in0(Mux2xBits16_inst2_O[15]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst24_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst3(
		.in0(Mux2xSInt9_inst0_O[3]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst3_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst4(
		.in0(Mux2xSInt9_inst0_O[4]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst4_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst5(
		.in0(Mux2xSInt9_inst0_O[5]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst5_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst6(
		.in0(Mux2xSInt9_inst0_O[6]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst6_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst7(
		.in0(Mux2xSInt9_inst0_O[7]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst7_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst8(
		.in0(Mux2xBits16_inst1_O[15]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst8_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst9(
		.in0(Mux2xBits16_inst2_O[0]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst9_out)
	);
	PEGEN_coreir_and #(.width(16)) magma_Bits_16_and_inst0(
		.in0(a),
		.in1(const_32768_16_out),
		.out(magma_Bits_16_and_inst0_out)
	);
	PEGEN_coreir_and #(.width(16)) magma_Bits_16_and_inst1(
		.in0(magma_Bits_16_shl_inst0_out),
		.in1(const_32640_16_out),
		.out(magma_Bits_16_and_inst1_out)
	);
	PEGEN_coreir_and #(.width(16)) magma_Bits_16_and_inst10(
		.in0(a),
		.in1(const_32768_16_out),
		.out(magma_Bits_16_and_inst10_out)
	);
	PEGEN_coreir_and #(.width(16)) magma_Bits_16_and_inst11(
		.in0(a),
		.in1(const_127_16_out),
		.out(magma_Bits_16_and_inst11_out)
	);
	PEGEN_coreir_and #(.width(16)) magma_Bits_16_and_inst12(
		.in0(Mux2xBits16_inst6_O),
		.in1(const_127_16_out),
		.out(magma_Bits_16_and_inst12_out)
	);
	PEGEN_coreir_and #(.width(16)) magma_Bits_16_and_inst2(
		.in0(a),
		.in1(const_127_16_out),
		.out(magma_Bits_16_and_inst2_out)
	);
	PEGEN_coreir_and #(.width(16)) magma_Bits_16_and_inst3(
		.in0(a),
		.in1(const_32768_16_out),
		.out(magma_Bits_16_and_inst3_out)
	);
	PEGEN_coreir_and #(.width(16)) magma_Bits_16_and_inst4(
		.in0(a),
		.in1(const_127_16_out),
		.out(magma_Bits_16_and_inst4_out)
	);
	PEGEN_coreir_and #(.width(16)) magma_Bits_16_and_inst5(
		.in0(a),
		.in1(const_32768_16_out),
		.out(magma_Bits_16_and_inst5_out)
	);
	PEGEN_coreir_and #(.width(16)) magma_Bits_16_and_inst6(
		.in0(b),
		.in1(const_32768_16_out),
		.out(magma_Bits_16_and_inst6_out)
	);
	PEGEN_coreir_and #(.width(16)) magma_Bits_16_and_inst7(
		.in0(a),
		.in1(const_127_16_out),
		.out(magma_Bits_16_and_inst7_out)
	);
	PEGEN_coreir_and #(.width(16)) magma_Bits_16_and_inst8(
		.in0(a),
		.in1(const_32768_16_out),
		.out(magma_Bits_16_and_inst8_out)
	);
	PEGEN_coreir_and #(.width(16)) magma_Bits_16_and_inst9(
		.in0(a),
		.in1(const_127_16_out),
		.out(magma_Bits_16_and_inst9_out)
	);
	PEGEN_coreir_eq #(.width(16)) magma_Bits_16_eq_inst0(
		.in0(magma_Bits_16_and_inst8_out),
		.in1(const_32768_16_out),
		.out(magma_Bits_16_eq_inst0_out)
	);
	PEGEN_coreir_eq #(.width(16)) magma_Bits_16_eq_inst1(
		.in0(magma_Bits_16_and_inst10_out),
		.in1(const_32768_16_out),
		.out(magma_Bits_16_eq_inst1_out)
	);
	PEGEN_coreir_lshr #(.width(16)) magma_Bits_16_lshr_inst0(
		.in0(Mux2xBits16_inst4_O),
		.in1(const_8_16_out),
		.out(magma_Bits_16_lshr_inst0_out)
	);
	wire [15:0] magma_Bits_16_lshr_inst1_in1;
	assign magma_Bits_16_lshr_inst1_in1 = {bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, magma_SInt_9_neg_inst1_out};
	PEGEN_coreir_lshr #(.width(16)) magma_Bits_16_lshr_inst1(
		.in0(magma_Bits_16_or_inst8_out),
		.in1(magma_Bits_16_lshr_inst1_in1),
		.out(magma_Bits_16_lshr_inst1_out)
	);
	PEGEN_coreir_or #(.width(16)) magma_Bits_16_or_inst0(
		.in0(Mux2xBits16_inst3_O),
		.in1(magma_Bits_16_and_inst1_out),
		.out(magma_Bits_16_or_inst0_out)
	);
	PEGEN_coreir_or #(.width(16)) magma_Bits_16_or_inst1(
		.in0(magma_Bits_16_or_inst0_out),
		.in1(Mux2xBits16_inst5_O),
		.out(magma_Bits_16_or_inst1_out)
	);
	PEGEN_coreir_or #(.width(16)) magma_Bits_16_or_inst2(
		.in0(magma_Bits_16_and_inst3_out),
		.in1(magma_Bits_16_shl_inst1_out),
		.out(magma_Bits_16_or_inst2_out)
	);
	PEGEN_coreir_or #(.width(16)) magma_Bits_16_or_inst3(
		.in0(magma_Bits_16_or_inst2_out),
		.in1(magma_Bits_16_and_inst4_out),
		.out(magma_Bits_16_or_inst3_out)
	);
	PEGEN_coreir_or #(.width(16)) magma_Bits_16_or_inst4(
		.in0(magma_Bits_16_and_inst5_out),
		.in1(magma_Bits_16_and_inst6_out),
		.out(magma_Bits_16_or_inst4_out)
	);
	PEGEN_coreir_or #(.width(16)) magma_Bits_16_or_inst5(
		.in0(magma_Bits_16_or_inst4_out),
		.in1(magma_Bits_16_shl_inst2_out),
		.out(magma_Bits_16_or_inst5_out)
	);
	PEGEN_coreir_or #(.width(16)) magma_Bits_16_or_inst6(
		.in0(magma_Bits_16_or_inst5_out),
		.in1(magma_Bits_16_and_inst7_out),
		.out(magma_Bits_16_or_inst6_out)
	);
	PEGEN_coreir_or #(.width(16)) magma_Bits_16_or_inst7(
		.in0(magma_Bits_16_and_inst9_out),
		.in1(const_128_16_out),
		.out(magma_Bits_16_or_inst7_out)
	);
	PEGEN_coreir_or #(.width(16)) magma_Bits_16_or_inst8(
		.in0(magma_Bits_16_and_inst11_out),
		.in1(const_128_16_out),
		.out(magma_Bits_16_or_inst8_out)
	);
	PEGEN_coreir_shl #(.width(16)) magma_Bits_16_shl_inst0(
		.in0(magma_SInt_16_add_inst0_out),
		.in1(const_7_16_out),
		.out(magma_Bits_16_shl_inst0_out)
	);
	wire [15:0] magma_Bits_16_shl_inst1_in0;
	assign magma_Bits_16_shl_inst1_in0 = {bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, magma_UInt_8_add_inst0_out};
	PEGEN_coreir_shl #(.width(16)) magma_Bits_16_shl_inst1(
		.in0(magma_Bits_16_shl_inst1_in0),
		.in1(const_7_16_out),
		.out(magma_Bits_16_shl_inst1_out)
	);
	wire [15:0] magma_Bits_16_shl_inst2_in0;
	assign magma_Bits_16_shl_inst2_in0 = {bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, magma_UInt_8_add_inst1_out};
	PEGEN_coreir_shl #(.width(16)) magma_Bits_16_shl_inst2(
		.in0(magma_Bits_16_shl_inst2_in0),
		.in1(const_7_16_out),
		.out(magma_Bits_16_shl_inst2_out)
	);
	wire [15:0] magma_Bits_16_shl_inst3_in1;
	assign magma_Bits_16_shl_inst3_in1 = {bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, magma_SInt_9_sub_inst2_out};
	PEGEN_coreir_shl #(.width(16)) magma_Bits_16_shl_inst3(
		.in0(magma_Bits_16_or_inst8_out),
		.in1(magma_Bits_16_shl_inst3_in1),
		.out(magma_Bits_16_shl_inst3_out)
	);
	PEGEN_coreir_eq #(.width(1)) magma_Bits_1_eq_inst0(
		.in0(signed_),
		.in1(const_1_1_out),
		.out(magma_Bits_1_eq_inst0_out)
	);
	PEGEN_coreir_lshr #(.width(23)) magma_Bits_23_lshr_inst0(
		.in0(Mux2xBits23_inst0_O),
		.in1(const_7_23_out),
		.out(magma_Bits_23_lshr_inst0_out)
	);
	wire [22:0] magma_Bits_23_shl_inst0_in0;
	assign magma_Bits_23_shl_inst0_in0 = {bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, magma_Bits_16_or_inst7_out};
	wire [22:0] magma_Bits_23_shl_inst0_in1;
	assign magma_Bits_23_shl_inst0_in1 = {bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, magma_SInt_9_sub_inst1_out};
	PEGEN_coreir_shl #(.width(23)) magma_Bits_23_shl_inst0(
		.in0(magma_Bits_23_shl_inst0_in0),
		.in1(magma_Bits_23_shl_inst0_in1),
		.out(magma_Bits_23_shl_inst0_out)
	);
	PEGEN_coreir_eq #(.width(3)) magma_Bits_3_eq_inst0(
		.in0(op),
		.in1(const_3_3_out),
		.out(magma_Bits_3_eq_inst0_out)
	);
	PEGEN_coreir_eq #(.width(3)) magma_Bits_3_eq_inst1(
		.in0(op),
		.in1(const_6_3_out),
		.out(magma_Bits_3_eq_inst1_out)
	);
	PEGEN_coreir_eq #(.width(3)) magma_Bits_3_eq_inst2(
		.in0(op),
		.in1(const_0_3_out),
		.out(magma_Bits_3_eq_inst2_out)
	);
	PEGEN_coreir_eq #(.width(3)) magma_Bits_3_eq_inst3(
		.in0(op),
		.in1(const_1_3_out),
		.out(magma_Bits_3_eq_inst3_out)
	);
	PEGEN_coreir_eq #(.width(3)) magma_Bits_3_eq_inst4(
		.in0(op),
		.in1(const_2_3_out),
		.out(magma_Bits_3_eq_inst4_out)
	);
	PEGEN_coreir_eq #(.width(3)) magma_Bits_3_eq_inst5(
		.in0(op),
		.in1(const_3_3_out),
		.out(magma_Bits_3_eq_inst5_out)
	);
	PEGEN_coreir_eq #(.width(3)) magma_Bits_3_eq_inst6(
		.in0(op),
		.in1(const_4_3_out),
		.out(magma_Bits_3_eq_inst6_out)
	);
	PEGEN_coreir_eq #(.width(3)) magma_Bits_3_eq_inst7(
		.in0(op),
		.in1(const_5_3_out),
		.out(magma_Bits_3_eq_inst7_out)
	);
	PEGEN_coreir_add #(.width(16)) magma_SInt_16_add_inst0(
		.in0(Mux2xSInt16_inst27_O),
		.in1(const_127_16_out),
		.out(magma_SInt_16_add_inst0_out)
	);
	PEGEN_coreir_and #(.width(16)) magma_SInt_16_and_inst0(
		.in0(magma_SInt_16_shl_inst0_out),
		.in1(Mux2xSInt16_inst24_O),
		.out(magma_SInt_16_and_inst0_out)
	);
	PEGEN_coreir_neg #(.width(16)) magma_SInt_16_neg_inst0(
		.in(a),
		.out(magma_SInt_16_neg_inst0_out)
	);
	wire [15:0] magma_SInt_16_neg_inst1_in;
	assign magma_SInt_16_neg_inst1_in = {magma_Bits_23_lshr_inst0_out[15], magma_Bits_23_lshr_inst0_out[14], magma_Bits_23_lshr_inst0_out[13], magma_Bits_23_lshr_inst0_out[12], magma_Bits_23_lshr_inst0_out[11], magma_Bits_23_lshr_inst0_out[10], magma_Bits_23_lshr_inst0_out[9], magma_Bits_23_lshr_inst0_out[8], magma_Bits_23_lshr_inst0_out[7], magma_Bits_23_lshr_inst0_out[6], magma_Bits_23_lshr_inst0_out[5], magma_Bits_23_lshr_inst0_out[4], magma_Bits_23_lshr_inst0_out[3], magma_Bits_23_lshr_inst0_out[2], magma_Bits_23_lshr_inst0_out[1], magma_Bits_23_lshr_inst0_out[0]};
	PEGEN_coreir_neg #(.width(16)) magma_SInt_16_neg_inst1(
		.in(magma_SInt_16_neg_inst1_in),
		.out(magma_SInt_16_neg_inst1_out)
	);
	PEGEN_coreir_neg #(.width(16)) magma_SInt_16_neg_inst2(
		.in(magma_Bits_16_and_inst12_out),
		.out(magma_SInt_16_neg_inst2_out)
	);
	PEGEN_coreir_sge #(.width(16)) magma_SInt_16_sge_inst0(
		.in0(Mux2xSInt16_inst27_O),
		.in1(const_0_16_out),
		.out(magma_SInt_16_sge_inst0_out)
	);
	PEGEN_coreir_shl #(.width(16)) magma_SInt_16_shl_inst0(
		.in0(Mux2xSInt16_inst25_O),
		.in1(Mux2xSInt16_inst26_O),
		.out(magma_SInt_16_shl_inst0_out)
	);
	PEGEN_coreir_sub #(.width(16)) magma_SInt_16_sub_inst0(
		.in0(const_7_16_out),
		.in1(Mux2xSInt16_inst7_O),
		.out(magma_SInt_16_sub_inst0_out)
	);
	PEGEN_coreir_sub #(.width(16)) magma_SInt_16_sub_inst1(
		.in0(const_15_16_out),
		.in1(Mux2xSInt16_inst23_O),
		.out(magma_SInt_16_sub_inst1_out)
	);
	PEGEN_coreir_neg #(.width(9)) magma_SInt_9_neg_inst0(
		.in(magma_SInt_9_sub_inst0_out),
		.out(magma_SInt_9_neg_inst0_out)
	);
	PEGEN_coreir_neg #(.width(9)) magma_SInt_9_neg_inst1(
		.in(magma_SInt_9_sub_inst2_out),
		.out(magma_SInt_9_neg_inst1_out)
	);
	PEGEN_coreir_slt #(.width(9)) magma_SInt_9_slt_inst0(
		.in0(magma_SInt_9_sub_inst0_out),
		.in1(const_0_9_out),
		.out(magma_SInt_9_slt_inst0_out)
	);
	PEGEN_coreir_slt #(.width(9)) magma_SInt_9_slt_inst1(
		.in0(magma_SInt_9_sub_inst1_out),
		.in1(const_0_9_out),
		.out(magma_SInt_9_slt_inst1_out)
	);
	PEGEN_coreir_slt #(.width(9)) magma_SInt_9_slt_inst2(
		.in0(magma_SInt_9_sub_inst2_out),
		.in1(const_0_9_out),
		.out(magma_SInt_9_slt_inst2_out)
	);
	wire [8:0] magma_SInt_9_sub_inst0_in0;
	assign magma_SInt_9_sub_inst0_in0 = {bit_const_0_None_out, a[14], a[13], a[12], a[11], a[10], a[9], a[8], a[7]};
	PEGEN_coreir_sub #(.width(9)) magma_SInt_9_sub_inst0(
		.in0(magma_SInt_9_sub_inst0_in0),
		.in1(const_127_9_out),
		.out(magma_SInt_9_sub_inst0_out)
	);
	wire [8:0] magma_SInt_9_sub_inst1_in0;
	assign magma_SInt_9_sub_inst1_in0 = {bit_const_0_None_out, a[14], a[13], a[12], a[11], a[10], a[9], a[8], a[7]};
	PEGEN_coreir_sub #(.width(9)) magma_SInt_9_sub_inst1(
		.in0(magma_SInt_9_sub_inst1_in0),
		.in1(const_127_9_out),
		.out(magma_SInt_9_sub_inst1_out)
	);
	wire [8:0] magma_SInt_9_sub_inst2_in0;
	assign magma_SInt_9_sub_inst2_in0 = {bit_const_0_None_out, a[14], a[13], a[12], a[11], a[10], a[9], a[8], a[7]};
	PEGEN_coreir_sub #(.width(9)) magma_SInt_9_sub_inst2(
		.in0(magma_SInt_9_sub_inst2_in0),
		.in1(const_127_9_out),
		.out(magma_SInt_9_sub_inst2_out)
	);
	wire [7:0] magma_UInt_8_add_inst0_in0;
	assign magma_UInt_8_add_inst0_in0 = {a[14], a[13], a[12], a[11], a[10], a[9], a[8], a[7]};
	wire [7:0] magma_UInt_8_add_inst0_in1;
	assign magma_UInt_8_add_inst0_in1 = {b[7], b[6], b[5], b[4], b[3], b[2], b[1], b[0]};
	PEGEN_coreir_add #(.width(8)) magma_UInt_8_add_inst0(
		.in0(magma_UInt_8_add_inst0_in0),
		.in1(magma_UInt_8_add_inst0_in1),
		.out(magma_UInt_8_add_inst0_out)
	);
	PEGEN_coreir_add #(.width(8)) magma_UInt_8_add_inst1(
		.in0(magma_UInt_8_sub_inst0_out),
		.in1(const_127_8_out),
		.out(magma_UInt_8_add_inst1_out)
	);
	wire [7:0] magma_UInt_8_sub_inst0_in0;
	assign magma_UInt_8_sub_inst0_in0 = {a[14], a[13], a[12], a[11], a[10], a[9], a[8], a[7]};
	wire [7:0] magma_UInt_8_sub_inst0_in1;
	assign magma_UInt_8_sub_inst0_in1 = {b[14], b[13], b[12], b[11], b[10], b[9], b[8], b[7]};
	PEGEN_coreir_sub #(.width(8)) magma_UInt_8_sub_inst0(
		.in0(magma_UInt_8_sub_inst0_in0),
		.in1(magma_UInt_8_sub_inst0_in1),
		.out(magma_UInt_8_sub_inst0_out)
	);
	wire [7:0] magma_UInt_8_ugt_inst0_in0;
	assign magma_UInt_8_ugt_inst0_in0 = {a[14], a[13], a[12], a[11], a[10], a[9], a[8], a[7]};
	PEGEN_coreir_ugt #(.width(8)) magma_UInt_8_ugt_inst0(
		.in0(magma_UInt_8_ugt_inst0_in0),
		.in1(const_142_8_out),
		.out(magma_UInt_8_ugt_inst0_out)
	);
	wire [8:0] magma_UInt_9_add_inst0_in0;
	assign magma_UInt_9_add_inst0_in0 = {bit_const_0_None_out, a[14], a[13], a[12], a[11], a[10], a[9], a[8], a[7]};
	wire [8:0] magma_UInt_9_add_inst0_in1;
	assign magma_UInt_9_add_inst0_in1 = {b[8], b[7], b[6], b[5], b[4], b[3], b[2], b[1], b[0]};
	PEGEN_coreir_add #(.width(9)) magma_UInt_9_add_inst0(
		.in0(magma_UInt_9_add_inst0_in0),
		.in1(magma_UInt_9_add_inst0_in1),
		.out(magma_UInt_9_add_inst0_out)
	);
	PEGEN_coreir_ugt #(.width(9)) magma_UInt_9_ugt_inst0(
		.in0(magma_UInt_9_add_inst0_out),
		.in1(const_255_9_out),
		.out(magma_UInt_9_ugt_inst0_out)
	);
	assign res = Mux2xBits16_inst19_O;
	assign res_p = Mux2xBit_inst10_O;
	assign V = Mux2xBit_inst9_O;
endmodule
module PEGEN_Cond (
	code,
	alu,
	lut,
	Z,
	N,
	C,
	V,
	O,
	CLK,
	ASYNCRESET
);
	input [4:0] code;
	input alu;
	input lut;
	input Z;
	input N;
	input C;
	input V;
	output wire O;
	input CLK;
	input ASYNCRESET;
	wire Mux2xBit_inst0_O;
	wire Mux2xBit_inst1_O;
	wire Mux2xBit_inst10_O;
	wire Mux2xBit_inst11_O;
	wire Mux2xBit_inst12_O;
	wire Mux2xBit_inst13_O;
	wire Mux2xBit_inst14_O;
	wire Mux2xBit_inst15_O;
	wire Mux2xBit_inst16_O;
	wire Mux2xBit_inst17_O;
	wire Mux2xBit_inst18_O;
	wire Mux2xBit_inst2_O;
	wire Mux2xBit_inst3_O;
	wire Mux2xBit_inst4_O;
	wire Mux2xBit_inst5_O;
	wire Mux2xBit_inst6_O;
	wire Mux2xBit_inst7_O;
	wire Mux2xBit_inst8_O;
	wire Mux2xBit_inst9_O;
	wire [4:0] const_0_5_out;
	wire [4:0] const_10_5_out;
	wire [4:0] const_11_5_out;
	wire [4:0] const_12_5_out;
	wire [4:0] const_13_5_out;
	wire [4:0] const_14_5_out;
	wire [4:0] const_15_5_out;
	wire [4:0] const_16_5_out;
	wire [4:0] const_17_5_out;
	wire [4:0] const_18_5_out;
	wire [4:0] const_1_5_out;
	wire [4:0] const_2_5_out;
	wire [4:0] const_3_5_out;
	wire [4:0] const_4_5_out;
	wire [4:0] const_5_5_out;
	wire [4:0] const_6_5_out;
	wire [4:0] const_7_5_out;
	wire [4:0] const_8_5_out;
	wire [4:0] const_9_5_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bit_and_inst1_out;
	wire magma_Bit_and_inst2_out;
	wire magma_Bit_and_inst3_out;
	wire magma_Bit_not_inst0_out;
	wire magma_Bit_not_inst1_out;
	wire magma_Bit_not_inst10_out;
	wire magma_Bit_not_inst11_out;
	wire magma_Bit_not_inst12_out;
	wire magma_Bit_not_inst2_out;
	wire magma_Bit_not_inst3_out;
	wire magma_Bit_not_inst4_out;
	wire magma_Bit_not_inst5_out;
	wire magma_Bit_not_inst6_out;
	wire magma_Bit_not_inst7_out;
	wire magma_Bit_not_inst8_out;
	wire magma_Bit_not_inst9_out;
	wire magma_Bit_or_inst0_out;
	wire magma_Bit_or_inst1_out;
	wire magma_Bit_or_inst2_out;
	wire magma_Bit_or_inst3_out;
	wire magma_Bit_or_inst4_out;
	wire magma_Bit_or_inst5_out;
	wire magma_Bit_xor_inst0_out;
	wire magma_Bit_xor_inst1_out;
	wire magma_Bit_xor_inst2_out;
	wire magma_Bit_xor_inst3_out;
	wire magma_Bits_5_eq_inst0_out;
	wire magma_Bits_5_eq_inst1_out;
	wire magma_Bits_5_eq_inst10_out;
	wire magma_Bits_5_eq_inst11_out;
	wire magma_Bits_5_eq_inst12_out;
	wire magma_Bits_5_eq_inst13_out;
	wire magma_Bits_5_eq_inst14_out;
	wire magma_Bits_5_eq_inst15_out;
	wire magma_Bits_5_eq_inst16_out;
	wire magma_Bits_5_eq_inst17_out;
	wire magma_Bits_5_eq_inst18_out;
	wire magma_Bits_5_eq_inst19_out;
	wire magma_Bits_5_eq_inst2_out;
	wire magma_Bits_5_eq_inst20_out;
	wire magma_Bits_5_eq_inst3_out;
	wire magma_Bits_5_eq_inst4_out;
	wire magma_Bits_5_eq_inst5_out;
	wire magma_Bits_5_eq_inst6_out;
	wire magma_Bits_5_eq_inst7_out;
	wire magma_Bits_5_eq_inst8_out;
	wire magma_Bits_5_eq_inst9_out;
	PEGEN_Mux2xBit Mux2xBit_inst0(
		.I0(magma_Bit_and_inst3_out),
		.I1(magma_Bit_or_inst5_out),
		.S(magma_Bits_5_eq_inst20_out),
		.O(Mux2xBit_inst0_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst1(
		.I0(Mux2xBit_inst0_O),
		.I1(magma_Bit_and_inst2_out),
		.S(magma_Bits_5_eq_inst19_out),
		.O(Mux2xBit_inst1_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst10(
		.I0(Mux2xBit_inst9_O),
		.I1(magma_Bit_and_inst0_out),
		.S(magma_Bits_5_eq_inst10_out),
		.O(Mux2xBit_inst10_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst11(
		.I0(Mux2xBit_inst10_O),
		.I1(magma_Bit_not_inst3_out),
		.S(magma_Bits_5_eq_inst9_out),
		.O(Mux2xBit_inst11_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst12(
		.I0(Mux2xBit_inst11_O),
		.I1(V),
		.S(magma_Bits_5_eq_inst8_out),
		.O(Mux2xBit_inst12_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst13(
		.I0(Mux2xBit_inst12_O),
		.I1(magma_Bit_not_inst2_out),
		.S(magma_Bits_5_eq_inst7_out),
		.O(Mux2xBit_inst13_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst14(
		.I0(Mux2xBit_inst13_O),
		.I1(N),
		.S(magma_Bits_5_eq_inst6_out),
		.O(Mux2xBit_inst14_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst15(
		.I0(Mux2xBit_inst14_O),
		.I1(magma_Bit_not_inst1_out),
		.S(magma_Bit_or_inst1_out),
		.O(Mux2xBit_inst15_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst16(
		.I0(Mux2xBit_inst15_O),
		.I1(C),
		.S(magma_Bit_or_inst0_out),
		.O(Mux2xBit_inst16_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst17(
		.I0(Mux2xBit_inst16_O),
		.I1(magma_Bit_not_inst0_out),
		.S(magma_Bits_5_eq_inst1_out),
		.O(Mux2xBit_inst17_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst18(
		.I0(Mux2xBit_inst17_O),
		.I1(Z),
		.S(magma_Bits_5_eq_inst0_out),
		.O(Mux2xBit_inst18_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst2(
		.I0(Mux2xBit_inst1_O),
		.I1(magma_Bit_or_inst4_out),
		.S(magma_Bits_5_eq_inst18_out),
		.O(Mux2xBit_inst2_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst3(
		.I0(Mux2xBit_inst2_O),
		.I1(lut),
		.S(magma_Bits_5_eq_inst17_out),
		.O(Mux2xBit_inst3_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst4(
		.I0(Mux2xBit_inst3_O),
		.I1(alu),
		.S(magma_Bits_5_eq_inst16_out),
		.O(Mux2xBit_inst4_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst5(
		.I0(Mux2xBit_inst4_O),
		.I1(magma_Bit_or_inst3_out),
		.S(magma_Bits_5_eq_inst15_out),
		.O(Mux2xBit_inst5_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst6(
		.I0(Mux2xBit_inst5_O),
		.I1(magma_Bit_and_inst1_out),
		.S(magma_Bits_5_eq_inst14_out),
		.O(Mux2xBit_inst6_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst7(
		.I0(Mux2xBit_inst6_O),
		.I1(magma_Bit_xor_inst1_out),
		.S(magma_Bits_5_eq_inst13_out),
		.O(Mux2xBit_inst7_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst8(
		.I0(Mux2xBit_inst7_O),
		.I1(magma_Bit_not_inst6_out),
		.S(magma_Bits_5_eq_inst12_out),
		.O(Mux2xBit_inst8_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst9(
		.I0(Mux2xBit_inst8_O),
		.I1(magma_Bit_or_inst2_out),
		.S(magma_Bits_5_eq_inst11_out),
		.O(Mux2xBit_inst9_O)
	);
	PEGEN_coreir_const #(
		.value(5'h00),
		.width(5)
	) const_0_5(.out(const_0_5_out));
	PEGEN_coreir_const #(
		.value(5'h0a),
		.width(5)
	) const_10_5(.out(const_10_5_out));
	PEGEN_coreir_const #(
		.value(5'h0b),
		.width(5)
	) const_11_5(.out(const_11_5_out));
	PEGEN_coreir_const #(
		.value(5'h0c),
		.width(5)
	) const_12_5(.out(const_12_5_out));
	PEGEN_coreir_const #(
		.value(5'h0d),
		.width(5)
	) const_13_5(.out(const_13_5_out));
	PEGEN_coreir_const #(
		.value(5'h0e),
		.width(5)
	) const_14_5(.out(const_14_5_out));
	PEGEN_coreir_const #(
		.value(5'h0f),
		.width(5)
	) const_15_5(.out(const_15_5_out));
	PEGEN_coreir_const #(
		.value(5'h10),
		.width(5)
	) const_16_5(.out(const_16_5_out));
	PEGEN_coreir_const #(
		.value(5'h11),
		.width(5)
	) const_17_5(.out(const_17_5_out));
	PEGEN_coreir_const #(
		.value(5'h12),
		.width(5)
	) const_18_5(.out(const_18_5_out));
	PEGEN_coreir_const #(
		.value(5'h01),
		.width(5)
	) const_1_5(.out(const_1_5_out));
	PEGEN_coreir_const #(
		.value(5'h02),
		.width(5)
	) const_2_5(.out(const_2_5_out));
	PEGEN_coreir_const #(
		.value(5'h03),
		.width(5)
	) const_3_5(.out(const_3_5_out));
	PEGEN_coreir_const #(
		.value(5'h04),
		.width(5)
	) const_4_5(.out(const_4_5_out));
	PEGEN_coreir_const #(
		.value(5'h05),
		.width(5)
	) const_5_5(.out(const_5_5_out));
	PEGEN_coreir_const #(
		.value(5'h06),
		.width(5)
	) const_6_5(.out(const_6_5_out));
	PEGEN_coreir_const #(
		.value(5'h07),
		.width(5)
	) const_7_5(.out(const_7_5_out));
	PEGEN_coreir_const #(
		.value(5'h08),
		.width(5)
	) const_8_5(.out(const_8_5_out));
	PEGEN_coreir_const #(
		.value(5'h09),
		.width(5)
	) const_9_5(.out(const_9_5_out));
	PEGEN_corebit_and magma_Bit_and_inst0(
		.in0(C),
		.in1(magma_Bit_not_inst4_out),
		.out(magma_Bit_and_inst0_out)
	);
	PEGEN_corebit_and magma_Bit_and_inst1(
		.in0(magma_Bit_not_inst7_out),
		.in1(magma_Bit_not_inst8_out),
		.out(magma_Bit_and_inst1_out)
	);
	PEGEN_corebit_and magma_Bit_and_inst2(
		.in0(magma_Bit_not_inst10_out),
		.in1(magma_Bit_not_inst11_out),
		.out(magma_Bit_and_inst2_out)
	);
	PEGEN_corebit_and magma_Bit_and_inst3(
		.in0(N),
		.in1(magma_Bit_not_inst12_out),
		.out(magma_Bit_and_inst3_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst0(
		.in(Z),
		.out(magma_Bit_not_inst0_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst1(
		.in(C),
		.out(magma_Bit_not_inst1_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst10(
		.in(N),
		.out(magma_Bit_not_inst10_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst11(
		.in(Z),
		.out(magma_Bit_not_inst11_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst12(
		.in(Z),
		.out(magma_Bit_not_inst12_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst2(
		.in(N),
		.out(magma_Bit_not_inst2_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst3(
		.in(V),
		.out(magma_Bit_not_inst3_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst4(
		.in(Z),
		.out(magma_Bit_not_inst4_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst5(
		.in(C),
		.out(magma_Bit_not_inst5_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst6(
		.in(magma_Bit_xor_inst0_out),
		.out(magma_Bit_not_inst6_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst7(
		.in(Z),
		.out(magma_Bit_not_inst7_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst8(
		.in(magma_Bit_xor_inst2_out),
		.out(magma_Bit_not_inst8_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst9(
		.in(N),
		.out(magma_Bit_not_inst9_out)
	);
	PEGEN_corebit_or magma_Bit_or_inst0(
		.in0(magma_Bits_5_eq_inst2_out),
		.in1(magma_Bits_5_eq_inst3_out),
		.out(magma_Bit_or_inst0_out)
	);
	PEGEN_corebit_or magma_Bit_or_inst1(
		.in0(magma_Bits_5_eq_inst4_out),
		.in1(magma_Bits_5_eq_inst5_out),
		.out(magma_Bit_or_inst1_out)
	);
	PEGEN_corebit_or magma_Bit_or_inst2(
		.in0(magma_Bit_not_inst5_out),
		.in1(Z),
		.out(magma_Bit_or_inst2_out)
	);
	PEGEN_corebit_or magma_Bit_or_inst3(
		.in0(Z),
		.in1(magma_Bit_xor_inst3_out),
		.out(magma_Bit_or_inst3_out)
	);
	PEGEN_corebit_or magma_Bit_or_inst4(
		.in0(magma_Bit_not_inst9_out),
		.in1(Z),
		.out(magma_Bit_or_inst4_out)
	);
	PEGEN_corebit_or magma_Bit_or_inst5(
		.in0(N),
		.in1(Z),
		.out(magma_Bit_or_inst5_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst0(
		.in0(N),
		.in1(V),
		.out(magma_Bit_xor_inst0_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst1(
		.in0(N),
		.in1(V),
		.out(magma_Bit_xor_inst1_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst2(
		.in0(N),
		.in1(V),
		.out(magma_Bit_xor_inst2_out)
	);
	PEGEN_corebit_xor magma_Bit_xor_inst3(
		.in0(N),
		.in1(V),
		.out(magma_Bit_xor_inst3_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst0(
		.in0(code),
		.in1(const_0_5_out),
		.out(magma_Bits_5_eq_inst0_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst1(
		.in0(code),
		.in1(const_1_5_out),
		.out(magma_Bits_5_eq_inst1_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst10(
		.in0(code),
		.in1(const_8_5_out),
		.out(magma_Bits_5_eq_inst10_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst11(
		.in0(code),
		.in1(const_9_5_out),
		.out(magma_Bits_5_eq_inst11_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst12(
		.in0(code),
		.in1(const_10_5_out),
		.out(magma_Bits_5_eq_inst12_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst13(
		.in0(code),
		.in1(const_11_5_out),
		.out(magma_Bits_5_eq_inst13_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst14(
		.in0(code),
		.in1(const_12_5_out),
		.out(magma_Bits_5_eq_inst14_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst15(
		.in0(code),
		.in1(const_13_5_out),
		.out(magma_Bits_5_eq_inst15_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst16(
		.in0(code),
		.in1(const_15_5_out),
		.out(magma_Bits_5_eq_inst16_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst17(
		.in0(code),
		.in1(const_14_5_out),
		.out(magma_Bits_5_eq_inst17_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst18(
		.in0(code),
		.in1(const_16_5_out),
		.out(magma_Bits_5_eq_inst18_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst19(
		.in0(code),
		.in1(const_17_5_out),
		.out(magma_Bits_5_eq_inst19_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst2(
		.in0(code),
		.in1(const_2_5_out),
		.out(magma_Bits_5_eq_inst2_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst20(
		.in0(code),
		.in1(const_18_5_out),
		.out(magma_Bits_5_eq_inst20_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst3(
		.in0(code),
		.in1(const_2_5_out),
		.out(magma_Bits_5_eq_inst3_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst4(
		.in0(code),
		.in1(const_3_5_out),
		.out(magma_Bits_5_eq_inst4_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst5(
		.in0(code),
		.in1(const_3_5_out),
		.out(magma_Bits_5_eq_inst5_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst6(
		.in0(code),
		.in1(const_4_5_out),
		.out(magma_Bits_5_eq_inst6_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst7(
		.in0(code),
		.in1(const_5_5_out),
		.out(magma_Bits_5_eq_inst7_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst8(
		.in0(code),
		.in1(const_6_5_out),
		.out(magma_Bits_5_eq_inst8_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst9(
		.in0(code),
		.in1(const_7_5_out),
		.out(magma_Bits_5_eq_inst9_out)
	);
	assign O = Mux2xBit_inst18_O;
endmodule
module PEGEN_ALU (
	alu,
	signed_,
	a,
	b,
	c,
	d,
	res,
	res_p,
	Z,
	N,
	C,
	V,
	CLK,
	ASYNCRESET
);
	input [4:0] alu;
	input [0:0] signed_;
	input [15:0] a;
	input [15:0] b;
	input [15:0] c;
	input d;
	output wire [15:0] res;
	output wire res_p;
	output wire Z;
	output wire N;
	output wire C;
	output wire V;
	input CLK;
	input ASYNCRESET;
	wire Mux2xBit_inst0_O;
	wire Mux2xBit_inst1_O;
	wire Mux2xBit_inst10_O;
	wire Mux2xBit_inst11_O;
	wire Mux2xBit_inst12_O;
	wire Mux2xBit_inst13_O;
	wire Mux2xBit_inst14_O;
	wire Mux2xBit_inst15_O;
	wire Mux2xBit_inst16_O;
	wire Mux2xBit_inst17_O;
	wire Mux2xBit_inst18_O;
	wire Mux2xBit_inst19_O;
	wire Mux2xBit_inst2_O;
	wire Mux2xBit_inst20_O;
	wire Mux2xBit_inst21_O;
	wire Mux2xBit_inst22_O;
	wire Mux2xBit_inst23_O;
	wire Mux2xBit_inst3_O;
	wire Mux2xBit_inst4_O;
	wire Mux2xBit_inst5_O;
	wire Mux2xBit_inst6_O;
	wire Mux2xBit_inst7_O;
	wire Mux2xBit_inst8_O;
	wire Mux2xBit_inst9_O;
	wire [15:0] Mux2xBits16_inst0_O;
	wire [15:0] Mux2xBits16_inst1_O;
	wire [15:0] Mux2xBits16_inst10_O;
	wire [15:0] Mux2xBits16_inst11_O;
	wire [15:0] Mux2xBits16_inst12_O;
	wire [15:0] Mux2xBits16_inst13_O;
	wire [15:0] Mux2xBits16_inst14_O;
	wire [15:0] Mux2xBits16_inst15_O;
	wire [15:0] Mux2xBits16_inst16_O;
	wire [15:0] Mux2xBits16_inst17_O;
	wire [15:0] Mux2xBits16_inst18_O;
	wire [15:0] Mux2xBits16_inst19_O;
	wire [15:0] Mux2xBits16_inst2_O;
	wire [15:0] Mux2xBits16_inst20_O;
	wire [15:0] Mux2xBits16_inst21_O;
	wire [15:0] Mux2xBits16_inst3_O;
	wire [15:0] Mux2xBits16_inst4_O;
	wire [15:0] Mux2xBits16_inst5_O;
	wire [15:0] Mux2xBits16_inst6_O;
	wire [15:0] Mux2xBits16_inst7_O;
	wire [15:0] Mux2xBits16_inst8_O;
	wire [15:0] Mux2xBits16_inst9_O;
	wire [15:0] Mux2xUInt16_inst0_O;
	wire [31:0] Mux2xUInt32_inst0_O;
	wire [31:0] Mux2xUInt32_inst1_O;
	wire bit_const_0_None_out;
	wire bit_const_1_None_out;
	wire [15:0] const_0_16_out;
	wire [4:0] const_0_5_out;
	wire [4:0] const_10_5_out;
	wire [4:0] const_11_5_out;
	wire [4:0] const_12_5_out;
	wire [4:0] const_13_5_out;
	wire [4:0] const_14_5_out;
	wire [4:0] const_15_5_out;
	wire [4:0] const_16_5_out;
	wire [4:0] const_17_5_out;
	wire [4:0] const_18_5_out;
	wire [4:0] const_19_5_out;
	wire [0:0] const_1_1_out;
	wire [4:0] const_1_5_out;
	wire [4:0] const_2_5_out;
	wire [4:0] const_3_5_out;
	wire [4:0] const_4_5_out;
	wire [4:0] const_5_5_out;
	wire [4:0] const_6_5_out;
	wire [4:0] const_7_5_out;
	wire [4:0] const_8_5_out;
	wire [4:0] const_9_5_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bit_and_inst1_out;
	wire magma_Bit_and_inst2_out;
	wire magma_Bit_and_inst3_out;
	wire magma_Bit_not_inst0_out;
	wire magma_Bit_not_inst1_out;
	wire magma_Bit_not_inst2_out;
	wire magma_Bit_or_inst0_out;
	wire magma_Bit_or_inst1_out;
	wire magma_Bit_or_inst10_out;
	wire magma_Bit_or_inst11_out;
	wire magma_Bit_or_inst12_out;
	wire magma_Bit_or_inst13_out;
	wire magma_Bit_or_inst2_out;
	wire magma_Bit_or_inst3_out;
	wire magma_Bit_or_inst4_out;
	wire magma_Bit_or_inst5_out;
	wire magma_Bit_or_inst6_out;
	wire magma_Bit_or_inst7_out;
	wire magma_Bit_or_inst8_out;
	wire magma_Bit_or_inst9_out;
	wire [15:0] magma_Bits_16_and_inst0_out;
	wire [15:0] magma_Bits_16_not_inst0_out;
	wire [15:0] magma_Bits_16_not_inst1_out;
	wire [15:0] magma_Bits_16_or_inst0_out;
	wire [15:0] magma_Bits_16_shl_inst0_out;
	wire [15:0] magma_Bits_16_xor_inst0_out;
	wire magma_Bits_1_eq_inst0_out;
	wire magma_Bits_1_eq_inst1_out;
	wire magma_Bits_1_eq_inst2_out;
	wire magma_Bits_1_eq_inst3_out;
	wire magma_Bits_5_eq_inst0_out;
	wire magma_Bits_5_eq_inst1_out;
	wire magma_Bits_5_eq_inst10_out;
	wire magma_Bits_5_eq_inst11_out;
	wire magma_Bits_5_eq_inst12_out;
	wire magma_Bits_5_eq_inst13_out;
	wire magma_Bits_5_eq_inst14_out;
	wire magma_Bits_5_eq_inst15_out;
	wire magma_Bits_5_eq_inst16_out;
	wire magma_Bits_5_eq_inst17_out;
	wire magma_Bits_5_eq_inst18_out;
	wire magma_Bits_5_eq_inst19_out;
	wire magma_Bits_5_eq_inst2_out;
	wire magma_Bits_5_eq_inst20_out;
	wire magma_Bits_5_eq_inst21_out;
	wire magma_Bits_5_eq_inst22_out;
	wire magma_Bits_5_eq_inst23_out;
	wire magma_Bits_5_eq_inst24_out;
	wire magma_Bits_5_eq_inst25_out;
	wire magma_Bits_5_eq_inst26_out;
	wire magma_Bits_5_eq_inst27_out;
	wire magma_Bits_5_eq_inst28_out;
	wire magma_Bits_5_eq_inst29_out;
	wire magma_Bits_5_eq_inst3_out;
	wire magma_Bits_5_eq_inst30_out;
	wire magma_Bits_5_eq_inst4_out;
	wire magma_Bits_5_eq_inst5_out;
	wire magma_Bits_5_eq_inst6_out;
	wire magma_Bits_5_eq_inst7_out;
	wire magma_Bits_5_eq_inst8_out;
	wire magma_Bits_5_eq_inst9_out;
	wire [15:0] magma_SInt_16_ashr_inst0_out;
	wire magma_SInt_16_eq_inst0_out;
	wire [15:0] magma_SInt_16_neg_inst0_out;
	wire magma_SInt_16_sge_inst0_out;
	wire magma_SInt_16_sle_inst0_out;
	wire magma_SInt_16_sle_inst1_out;
	wire [15:0] magma_UInt_16_lshr_inst0_out;
	wire magma_UInt_16_uge_inst0_out;
	wire magma_UInt_16_ule_inst0_out;
	wire [16:0] magma_UInt_17_add_inst0_out;
	wire [16:0] magma_UInt_17_add_inst1_out;
	wire [16:0] magma_UInt_17_add_inst2_out;
	wire [16:0] magma_UInt_17_add_inst3_out;
	wire [31:0] magma_UInt_32_mul_inst0_out;
	PEGEN_Mux2xBit Mux2xBit_inst0(
		.I0(magma_UInt_16_ule_inst0_out),
		.I1(magma_SInt_16_sle_inst0_out),
		.S(magma_Bits_1_eq_inst1_out),
		.O(Mux2xBit_inst0_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst1(
		.I0(magma_UInt_16_uge_inst0_out),
		.I1(magma_SInt_16_sge_inst0_out),
		.S(magma_Bits_1_eq_inst2_out),
		.O(Mux2xBit_inst1_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst10(
		.I0(Mux2xBit_inst9_O),
		.I1(bit_const_0_None_out),
		.S(magma_Bits_5_eq_inst18_out),
		.O(Mux2xBit_inst10_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst11(
		.I0(Mux2xBit_inst10_O),
		.I1(a[15]),
		.S(magma_Bits_5_eq_inst17_out),
		.O(Mux2xBit_inst11_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst12(
		.I0(bit_const_0_None_out),
		.I1(bit_const_0_None_out),
		.S(magma_Bits_5_eq_inst16_out),
		.O(Mux2xBit_inst12_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst13(
		.I0(bit_const_0_None_out),
		.I1(bit_const_0_None_out),
		.S(magma_Bits_5_eq_inst16_out),
		.O(Mux2xBit_inst13_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst14(
		.I0(Mux2xBit_inst11_O),
		.I1(bit_const_0_None_out),
		.S(magma_Bits_5_eq_inst16_out),
		.O(Mux2xBit_inst14_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst15(
		.I0(Mux2xBit_inst12_O),
		.I1(bit_const_0_None_out),
		.S(magma_Bits_5_eq_inst15_out),
		.O(Mux2xBit_inst15_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst16(
		.I0(Mux2xBit_inst13_O),
		.I1(bit_const_0_None_out),
		.S(magma_Bits_5_eq_inst15_out),
		.O(Mux2xBit_inst16_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst17(
		.I0(Mux2xBit_inst14_O),
		.I1(bit_const_0_None_out),
		.S(magma_Bits_5_eq_inst15_out),
		.O(Mux2xBit_inst17_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst18(
		.I0(Mux2xBit_inst15_O),
		.I1(bit_const_0_None_out),
		.S(magma_Bits_5_eq_inst14_out),
		.O(Mux2xBit_inst18_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst19(
		.I0(Mux2xBit_inst16_O),
		.I1(bit_const_0_None_out),
		.S(magma_Bits_5_eq_inst14_out),
		.O(Mux2xBit_inst19_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst2(
		.I0(bit_const_0_None_out),
		.I1(bit_const_1_None_out),
		.S(magma_Bit_or_inst6_out),
		.O(Mux2xBit_inst2_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst20(
		.I0(Mux2xBit_inst17_O),
		.I1(bit_const_0_None_out),
		.S(magma_Bits_5_eq_inst14_out),
		.O(Mux2xBit_inst20_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst21(
		.I0(Mux2xBit_inst18_O),
		.I1(magma_UInt_17_add_inst1_out[16]),
		.S(magma_Bit_or_inst7_out),
		.O(Mux2xBit_inst21_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst22(
		.I0(Mux2xBit_inst19_O),
		.I1(magma_Bit_or_inst8_out),
		.S(magma_Bit_or_inst7_out),
		.O(Mux2xBit_inst22_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst23(
		.I0(Mux2xBit_inst20_O),
		.I1(magma_UInt_17_add_inst1_out[16]),
		.S(magma_Bit_or_inst7_out),
		.O(Mux2xBit_inst23_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst3(
		.I0(bit_const_0_None_out),
		.I1(bit_const_0_None_out),
		.S(magma_Bits_5_eq_inst30_out),
		.O(Mux2xBit_inst3_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst4(
		.I0(Mux2xBit_inst3_O),
		.I1(bit_const_0_None_out),
		.S(magma_Bit_or_inst13_out),
		.O(Mux2xBit_inst4_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst5(
		.I0(Mux2xBit_inst4_O),
		.I1(bit_const_0_None_out),
		.S(magma_Bits_5_eq_inst23_out),
		.O(Mux2xBit_inst5_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst6(
		.I0(Mux2xBit_inst5_O),
		.I1(bit_const_0_None_out),
		.S(magma_Bits_5_eq_inst22_out),
		.O(Mux2xBit_inst6_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst7(
		.I0(Mux2xBit_inst6_O),
		.I1(bit_const_0_None_out),
		.S(magma_Bits_5_eq_inst21_out),
		.O(Mux2xBit_inst7_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst8(
		.I0(Mux2xBit_inst7_O),
		.I1(bit_const_0_None_out),
		.S(magma_Bits_5_eq_inst20_out),
		.O(Mux2xBit_inst8_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst9(
		.I0(Mux2xBit_inst8_O),
		.I1(bit_const_0_None_out),
		.S(magma_Bits_5_eq_inst19_out),
		.O(Mux2xBit_inst9_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst0(
		.I0(b),
		.I1(a),
		.S(Mux2xBit_inst0_O),
		.O(Mux2xBits16_inst0_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst1(
		.I0(b),
		.I1(Mux2xBits16_inst0_O),
		.S(magma_Bits_5_eq_inst0_out),
		.O(Mux2xBits16_inst1_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst10(
		.I0(Mux2xBits16_inst9_O),
		.I1(magma_UInt_17_add_inst3_out[15:0]),
		.S(magma_Bit_or_inst13_out),
		.O(Mux2xBits16_inst10_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst11(
		.I0(Mux2xBits16_inst10_O),
		.I1(magma_Bits_16_shl_inst0_out),
		.S(magma_Bits_5_eq_inst23_out),
		.O(Mux2xBits16_inst11_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst12(
		.I0(Mux2xBits16_inst11_O),
		.I1(Mux2xBits16_inst4_O),
		.S(magma_Bits_5_eq_inst22_out),
		.O(Mux2xBits16_inst12_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst13(
		.I0(Mux2xBits16_inst12_O),
		.I1(magma_Bits_16_xor_inst0_out),
		.S(magma_Bits_5_eq_inst21_out),
		.O(Mux2xBits16_inst13_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst14(
		.I0(Mux2xBits16_inst13_O),
		.I1(magma_Bits_16_or_inst0_out),
		.S(magma_Bits_5_eq_inst20_out),
		.O(Mux2xBits16_inst14_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst15(
		.I0(Mux2xBits16_inst14_O),
		.I1(magma_Bits_16_and_inst0_out),
		.S(magma_Bits_5_eq_inst19_out),
		.O(Mux2xBits16_inst15_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst16(
		.I0(Mux2xBits16_inst15_O),
		.I1(Mux2xBits16_inst8_O),
		.S(magma_Bits_5_eq_inst18_out),
		.O(Mux2xBits16_inst16_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst17(
		.I0(Mux2xBits16_inst16_O),
		.I1(Mux2xBits16_inst7_O),
		.S(magma_Bits_5_eq_inst17_out),
		.O(Mux2xBits16_inst17_O)
	);
	wire [15:0] Mux2xBits16_inst18_I1;
	assign Mux2xBits16_inst18_I1 = {magma_UInt_32_mul_inst0_out[31], magma_UInt_32_mul_inst0_out[30], magma_UInt_32_mul_inst0_out[29], magma_UInt_32_mul_inst0_out[28], magma_UInt_32_mul_inst0_out[27], magma_UInt_32_mul_inst0_out[26], magma_UInt_32_mul_inst0_out[25], magma_UInt_32_mul_inst0_out[24], magma_UInt_32_mul_inst0_out[23], magma_UInt_32_mul_inst0_out[22], magma_UInt_32_mul_inst0_out[21], magma_UInt_32_mul_inst0_out[20], magma_UInt_32_mul_inst0_out[19], magma_UInt_32_mul_inst0_out[18], magma_UInt_32_mul_inst0_out[17], magma_UInt_32_mul_inst0_out[16]};
	PEGEN_Mux2xBits16 Mux2xBits16_inst18(
		.I0(Mux2xBits16_inst17_O),
		.I1(Mux2xBits16_inst18_I1),
		.S(magma_Bits_5_eq_inst16_out),
		.O(Mux2xBits16_inst18_O)
	);
	wire [15:0] Mux2xBits16_inst19_I1;
	assign Mux2xBits16_inst19_I1 = {magma_UInt_32_mul_inst0_out[23], magma_UInt_32_mul_inst0_out[22], magma_UInt_32_mul_inst0_out[21], magma_UInt_32_mul_inst0_out[20], magma_UInt_32_mul_inst0_out[19], magma_UInt_32_mul_inst0_out[18], magma_UInt_32_mul_inst0_out[17], magma_UInt_32_mul_inst0_out[16], magma_UInt_32_mul_inst0_out[15], magma_UInt_32_mul_inst0_out[14], magma_UInt_32_mul_inst0_out[13], magma_UInt_32_mul_inst0_out[12], magma_UInt_32_mul_inst0_out[11], magma_UInt_32_mul_inst0_out[10], magma_UInt_32_mul_inst0_out[9], magma_UInt_32_mul_inst0_out[8]};
	PEGEN_Mux2xBits16 Mux2xBits16_inst19(
		.I0(Mux2xBits16_inst18_O),
		.I1(Mux2xBits16_inst19_I1),
		.S(magma_Bits_5_eq_inst15_out),
		.O(Mux2xBits16_inst19_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst2(
		.I0(c),
		.I1(Mux2xBits16_inst1_O),
		.S(Mux2xBit_inst1_O),
		.O(Mux2xBits16_inst2_O)
	);
	wire [15:0] Mux2xBits16_inst20_I1;
	assign Mux2xBits16_inst20_I1 = {magma_UInt_32_mul_inst0_out[15], magma_UInt_32_mul_inst0_out[14], magma_UInt_32_mul_inst0_out[13], magma_UInt_32_mul_inst0_out[12], magma_UInt_32_mul_inst0_out[11], magma_UInt_32_mul_inst0_out[10], magma_UInt_32_mul_inst0_out[9], magma_UInt_32_mul_inst0_out[8], magma_UInt_32_mul_inst0_out[7], magma_UInt_32_mul_inst0_out[6], magma_UInt_32_mul_inst0_out[5], magma_UInt_32_mul_inst0_out[4], magma_UInt_32_mul_inst0_out[3], magma_UInt_32_mul_inst0_out[2], magma_UInt_32_mul_inst0_out[1], magma_UInt_32_mul_inst0_out[0]};
	PEGEN_Mux2xBits16 Mux2xBits16_inst20(
		.I0(Mux2xBits16_inst19_O),
		.I1(Mux2xBits16_inst20_I1),
		.S(magma_Bits_5_eq_inst14_out),
		.O(Mux2xBits16_inst20_O)
	);
	wire [15:0] Mux2xBits16_inst21_I1;
	assign Mux2xBits16_inst21_I1 = {magma_UInt_17_add_inst1_out[15], magma_UInt_17_add_inst1_out[14], magma_UInt_17_add_inst1_out[13], magma_UInt_17_add_inst1_out[12], magma_UInt_17_add_inst1_out[11], magma_UInt_17_add_inst1_out[10], magma_UInt_17_add_inst1_out[9], magma_UInt_17_add_inst1_out[8], magma_UInt_17_add_inst1_out[7], magma_UInt_17_add_inst1_out[6], magma_UInt_17_add_inst1_out[5], magma_UInt_17_add_inst1_out[4], magma_UInt_17_add_inst1_out[3], magma_UInt_17_add_inst1_out[2], magma_UInt_17_add_inst1_out[1], magma_UInt_17_add_inst1_out[0]};
	PEGEN_Mux2xBits16 Mux2xBits16_inst21(
		.I0(Mux2xBits16_inst20_O),
		.I1(Mux2xBits16_inst21_I1),
		.S(magma_Bit_or_inst7_out),
		.O(Mux2xBits16_inst21_O)
	);
	wire [15:0] Mux2xBits16_inst3_I1;
	assign Mux2xBits16_inst3_I1 = {magma_UInt_32_mul_inst0_out[15], magma_UInt_32_mul_inst0_out[14], magma_UInt_32_mul_inst0_out[13], magma_UInt_32_mul_inst0_out[12], magma_UInt_32_mul_inst0_out[11], magma_UInt_32_mul_inst0_out[10], magma_UInt_32_mul_inst0_out[9], magma_UInt_32_mul_inst0_out[8], magma_UInt_32_mul_inst0_out[7], magma_UInt_32_mul_inst0_out[6], magma_UInt_32_mul_inst0_out[5], magma_UInt_32_mul_inst0_out[4], magma_UInt_32_mul_inst0_out[3], magma_UInt_32_mul_inst0_out[2], magma_UInt_32_mul_inst0_out[1], magma_UInt_32_mul_inst0_out[0]};
	PEGEN_Mux2xBits16 Mux2xBits16_inst3(
		.I0(a),
		.I1(Mux2xBits16_inst3_I1),
		.S(magma_Bits_5_eq_inst1_out),
		.O(Mux2xBits16_inst3_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst4(
		.I0(magma_UInt_16_lshr_inst0_out),
		.I1(magma_SInt_16_ashr_inst0_out),
		.S(magma_Bits_1_eq_inst3_out),
		.O(Mux2xBits16_inst4_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst5(
		.I0(b),
		.I1(magma_Bits_16_not_inst0_out),
		.S(magma_Bit_or_inst1_out),
		.O(Mux2xBits16_inst5_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst6(
		.I0(c),
		.I1(magma_Bits_16_not_inst1_out),
		.S(magma_Bit_or_inst6_out),
		.O(Mux2xBits16_inst6_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst7(
		.I0(magma_SInt_16_neg_inst0_out),
		.I1(a),
		.S(magma_SInt_16_sle_inst1_out),
		.O(Mux2xBits16_inst7_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst8(
		.I0(Mux2xBits16_inst5_O),
		.I1(a),
		.S(d),
		.O(Mux2xBits16_inst8_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst9(
		.I0(Mux2xBits16_inst4_O),
		.I1(Mux2xBits16_inst2_O),
		.S(magma_Bits_5_eq_inst30_out),
		.O(Mux2xBits16_inst9_O)
	);
	wire [15:0] Mux2xUInt16_inst0_I0;
	assign Mux2xUInt16_inst0_I0 = {magma_UInt_32_mul_inst0_out[15], magma_UInt_32_mul_inst0_out[14], magma_UInt_32_mul_inst0_out[13], magma_UInt_32_mul_inst0_out[12], magma_UInt_32_mul_inst0_out[11], magma_UInt_32_mul_inst0_out[10], magma_UInt_32_mul_inst0_out[9], magma_UInt_32_mul_inst0_out[8], magma_UInt_32_mul_inst0_out[7], magma_UInt_32_mul_inst0_out[6], magma_UInt_32_mul_inst0_out[5], magma_UInt_32_mul_inst0_out[4], magma_UInt_32_mul_inst0_out[3], magma_UInt_32_mul_inst0_out[2], magma_UInt_32_mul_inst0_out[1], magma_UInt_32_mul_inst0_out[0]};
	wire [15:0] Mux2xUInt16_inst0_I1;
	assign Mux2xUInt16_inst0_I1 = {magma_UInt_17_add_inst1_out[15], magma_UInt_17_add_inst1_out[14], magma_UInt_17_add_inst1_out[13], magma_UInt_17_add_inst1_out[12], magma_UInt_17_add_inst1_out[11], magma_UInt_17_add_inst1_out[10], magma_UInt_17_add_inst1_out[9], magma_UInt_17_add_inst1_out[8], magma_UInt_17_add_inst1_out[7], magma_UInt_17_add_inst1_out[6], magma_UInt_17_add_inst1_out[5], magma_UInt_17_add_inst1_out[4], magma_UInt_17_add_inst1_out[3], magma_UInt_17_add_inst1_out[2], magma_UInt_17_add_inst1_out[1], magma_UInt_17_add_inst1_out[0]};
	PEGEN_Mux2xUInt16 Mux2xUInt16_inst0(
		.I0(Mux2xUInt16_inst0_I0),
		.I1(Mux2xUInt16_inst0_I1),
		.S(magma_Bit_or_inst4_out),
		.O(Mux2xUInt16_inst0_O)
	);
	wire [31:0] Mux2xUInt32_inst0_I0;
	assign Mux2xUInt32_inst0_I0 = {bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, a};
	wire [31:0] Mux2xUInt32_inst0_I1;
	assign Mux2xUInt32_inst0_I1 = {a[15], a[15], a[15], a[15], a[15], a[15], a[15], a[15], a[15], a[15], a[15], a[15], a[15], a[15], a[15], a[15], a};
	PEGEN_Mux2xUInt32 Mux2xUInt32_inst0(
		.I0(Mux2xUInt32_inst0_I0),
		.I1(Mux2xUInt32_inst0_I1),
		.S(magma_Bits_1_eq_inst0_out),
		.O(Mux2xUInt32_inst0_O)
	);
	wire [31:0] Mux2xUInt32_inst1_I0;
	assign Mux2xUInt32_inst1_I0 = {bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, b};
	wire [31:0] Mux2xUInt32_inst1_I1;
	assign Mux2xUInt32_inst1_I1 = {b[15], b[15], b[15], b[15], b[15], b[15], b[15], b[15], b[15], b[15], b[15], b[15], b[15], b[15], b[15], b[15], b};
	PEGEN_Mux2xUInt32 Mux2xUInt32_inst1(
		.I0(Mux2xUInt32_inst1_I0),
		.I1(Mux2xUInt32_inst1_I1),
		.S(magma_Bits_1_eq_inst0_out),
		.O(Mux2xUInt32_inst1_O)
	);
	PEGEN_corebit_const #(.value(1'b0)) bit_const_0_None(.out(bit_const_0_None_out));
	PEGEN_corebit_const #(.value(1'b1)) bit_const_1_None(.out(bit_const_1_None_out));
	PEGEN_coreir_const #(
		.value(16'h0000),
		.width(16)
	) const_0_16(.out(const_0_16_out));
	PEGEN_coreir_const #(
		.value(5'h00),
		.width(5)
	) const_0_5(.out(const_0_5_out));
	PEGEN_coreir_const #(
		.value(5'h0a),
		.width(5)
	) const_10_5(.out(const_10_5_out));
	PEGEN_coreir_const #(
		.value(5'h0b),
		.width(5)
	) const_11_5(.out(const_11_5_out));
	PEGEN_coreir_const #(
		.value(5'h0c),
		.width(5)
	) const_12_5(.out(const_12_5_out));
	PEGEN_coreir_const #(
		.value(5'h0d),
		.width(5)
	) const_13_5(.out(const_13_5_out));
	PEGEN_coreir_const #(
		.value(5'h0e),
		.width(5)
	) const_14_5(.out(const_14_5_out));
	PEGEN_coreir_const #(
		.value(5'h0f),
		.width(5)
	) const_15_5(.out(const_15_5_out));
	PEGEN_coreir_const #(
		.value(5'h10),
		.width(5)
	) const_16_5(.out(const_16_5_out));
	PEGEN_coreir_const #(
		.value(5'h11),
		.width(5)
	) const_17_5(.out(const_17_5_out));
	PEGEN_coreir_const #(
		.value(5'h12),
		.width(5)
	) const_18_5(.out(const_18_5_out));
	PEGEN_coreir_const #(
		.value(5'h13),
		.width(5)
	) const_19_5(.out(const_19_5_out));
	PEGEN_coreir_const #(
		.value(1'h1),
		.width(1)
	) const_1_1(.out(const_1_1_out));
	PEGEN_coreir_const #(
		.value(5'h01),
		.width(5)
	) const_1_5(.out(const_1_5_out));
	PEGEN_coreir_const #(
		.value(5'h02),
		.width(5)
	) const_2_5(.out(const_2_5_out));
	PEGEN_coreir_const #(
		.value(5'h03),
		.width(5)
	) const_3_5(.out(const_3_5_out));
	PEGEN_coreir_const #(
		.value(5'h04),
		.width(5)
	) const_4_5(.out(const_4_5_out));
	PEGEN_coreir_const #(
		.value(5'h05),
		.width(5)
	) const_5_5(.out(const_5_5_out));
	PEGEN_coreir_const #(
		.value(5'h06),
		.width(5)
	) const_6_5(.out(const_6_5_out));
	PEGEN_coreir_const #(
		.value(5'h07),
		.width(5)
	) const_7_5(.out(const_7_5_out));
	PEGEN_coreir_const #(
		.value(5'h08),
		.width(5)
	) const_8_5(.out(const_8_5_out));
	PEGEN_coreir_const #(
		.value(5'h09),
		.width(5)
	) const_9_5(.out(const_9_5_out));
	PEGEN_corebit_and magma_Bit_and_inst0(
		.in0(a[15]),
		.in1(Mux2xBits16_inst5_O[15]),
		.out(magma_Bit_and_inst0_out)
	);
	PEGEN_corebit_and magma_Bit_and_inst1(
		.in0(magma_Bit_and_inst0_out),
		.in1(magma_Bit_not_inst0_out),
		.out(magma_Bit_and_inst1_out)
	);
	PEGEN_corebit_and magma_Bit_and_inst2(
		.in0(magma_Bit_not_inst1_out),
		.in1(magma_Bit_not_inst2_out),
		.out(magma_Bit_and_inst2_out)
	);
	PEGEN_corebit_and magma_Bit_and_inst3(
		.in0(magma_Bit_and_inst2_out),
		.in1(magma_UInt_17_add_inst1_out[15]),
		.out(magma_Bit_and_inst3_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst0(
		.in(magma_UInt_17_add_inst1_out[15]),
		.out(magma_Bit_not_inst0_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst1(
		.in(a[15]),
		.out(magma_Bit_not_inst1_out)
	);
	PEGEN_corebit_not magma_Bit_not_inst2(
		.in(Mux2xBits16_inst5_O[15]),
		.out(magma_Bit_not_inst2_out)
	);
	PEGEN_corebit_or magma_Bit_or_inst0(
		.in0(magma_Bits_5_eq_inst2_out),
		.in1(magma_Bits_5_eq_inst3_out),
		.out(magma_Bit_or_inst0_out)
	);
	PEGEN_corebit_or magma_Bit_or_inst1(
		.in0(magma_Bit_or_inst0_out),
		.in1(magma_Bits_5_eq_inst4_out),
		.out(magma_Bit_or_inst1_out)
	);
	PEGEN_corebit_or magma_Bit_or_inst10(
		.in0(magma_Bit_or_inst9_out),
		.in1(magma_Bits_5_eq_inst26_out),
		.out(magma_Bit_or_inst10_out)
	);
	PEGEN_corebit_or magma_Bit_or_inst11(
		.in0(magma_Bit_or_inst10_out),
		.in1(magma_Bits_5_eq_inst27_out),
		.out(magma_Bit_or_inst11_out)
	);
	PEGEN_corebit_or magma_Bit_or_inst12(
		.in0(magma_Bit_or_inst11_out),
		.in1(magma_Bits_5_eq_inst28_out),
		.out(magma_Bit_or_inst12_out)
	);
	PEGEN_corebit_or magma_Bit_or_inst13(
		.in0(magma_Bit_or_inst12_out),
		.in1(magma_Bits_5_eq_inst29_out),
		.out(magma_Bit_or_inst13_out)
	);
	PEGEN_corebit_or magma_Bit_or_inst2(
		.in0(magma_Bits_5_eq_inst5_out),
		.in1(magma_Bits_5_eq_inst6_out),
		.out(magma_Bit_or_inst2_out)
	);
	PEGEN_corebit_or magma_Bit_or_inst3(
		.in0(magma_Bit_or_inst2_out),
		.in1(magma_Bits_5_eq_inst7_out),
		.out(magma_Bit_or_inst3_out)
	);
	PEGEN_corebit_or magma_Bit_or_inst4(
		.in0(magma_Bit_or_inst3_out),
		.in1(magma_Bits_5_eq_inst8_out),
		.out(magma_Bit_or_inst4_out)
	);
	PEGEN_corebit_or magma_Bit_or_inst5(
		.in0(magma_Bits_5_eq_inst9_out),
		.in1(magma_Bits_5_eq_inst10_out),
		.out(magma_Bit_or_inst5_out)
	);
	PEGEN_corebit_or magma_Bit_or_inst6(
		.in0(magma_Bit_or_inst5_out),
		.in1(magma_Bits_5_eq_inst11_out),
		.out(magma_Bit_or_inst6_out)
	);
	PEGEN_corebit_or magma_Bit_or_inst7(
		.in0(magma_Bits_5_eq_inst12_out),
		.in1(magma_Bits_5_eq_inst13_out),
		.out(magma_Bit_or_inst7_out)
	);
	PEGEN_corebit_or magma_Bit_or_inst8(
		.in0(magma_Bit_and_inst1_out),
		.in1(magma_Bit_and_inst3_out),
		.out(magma_Bit_or_inst8_out)
	);
	PEGEN_corebit_or magma_Bit_or_inst9(
		.in0(magma_Bits_5_eq_inst24_out),
		.in1(magma_Bits_5_eq_inst25_out),
		.out(magma_Bit_or_inst9_out)
	);
	PEGEN_coreir_and #(.width(16)) magma_Bits_16_and_inst0(
		.in0(a),
		.in1(Mux2xBits16_inst5_O),
		.out(magma_Bits_16_and_inst0_out)
	);
	PEGEN_coreir_not #(.width(16)) magma_Bits_16_not_inst0(
		.in(b),
		.out(magma_Bits_16_not_inst0_out)
	);
	PEGEN_coreir_not #(.width(16)) magma_Bits_16_not_inst1(
		.in(c),
		.out(magma_Bits_16_not_inst1_out)
	);
	PEGEN_coreir_or #(.width(16)) magma_Bits_16_or_inst0(
		.in0(a),
		.in1(Mux2xBits16_inst5_O),
		.out(magma_Bits_16_or_inst0_out)
	);
	PEGEN_coreir_shl #(.width(16)) magma_Bits_16_shl_inst0(
		.in0(a),
		.in1(Mux2xBits16_inst5_O),
		.out(magma_Bits_16_shl_inst0_out)
	);
	PEGEN_coreir_xor #(.width(16)) magma_Bits_16_xor_inst0(
		.in0(a),
		.in1(Mux2xBits16_inst5_O),
		.out(magma_Bits_16_xor_inst0_out)
	);
	PEGEN_coreir_eq #(.width(1)) magma_Bits_1_eq_inst0(
		.in0(signed_),
		.in1(const_1_1_out),
		.out(magma_Bits_1_eq_inst0_out)
	);
	PEGEN_coreir_eq #(.width(1)) magma_Bits_1_eq_inst1(
		.in0(signed_),
		.in1(const_1_1_out),
		.out(magma_Bits_1_eq_inst1_out)
	);
	PEGEN_coreir_eq #(.width(1)) magma_Bits_1_eq_inst2(
		.in0(signed_),
		.in1(const_1_1_out),
		.out(magma_Bits_1_eq_inst2_out)
	);
	PEGEN_coreir_eq #(.width(1)) magma_Bits_1_eq_inst3(
		.in0(signed_),
		.in1(const_1_1_out),
		.out(magma_Bits_1_eq_inst3_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst0(
		.in0(alu),
		.in1(const_18_5_out),
		.out(magma_Bits_5_eq_inst0_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst1(
		.in0(alu),
		.in1(const_19_5_out),
		.out(magma_Bits_5_eq_inst1_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst10(
		.in0(alu),
		.in1(const_15_5_out),
		.out(magma_Bits_5_eq_inst10_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst11(
		.in0(alu),
		.in1(const_17_5_out),
		.out(magma_Bits_5_eq_inst11_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst12(
		.in0(alu),
		.in1(const_0_5_out),
		.out(magma_Bits_5_eq_inst12_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst13(
		.in0(alu),
		.in1(const_1_5_out),
		.out(magma_Bits_5_eq_inst13_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst14(
		.in0(alu),
		.in1(const_4_5_out),
		.out(magma_Bits_5_eq_inst14_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst15(
		.in0(alu),
		.in1(const_5_5_out),
		.out(magma_Bits_5_eq_inst15_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst16(
		.in0(alu),
		.in1(const_6_5_out),
		.out(magma_Bits_5_eq_inst16_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst17(
		.in0(alu),
		.in1(const_2_5_out),
		.out(magma_Bits_5_eq_inst17_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst18(
		.in0(alu),
		.in1(const_3_5_out),
		.out(magma_Bits_5_eq_inst18_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst19(
		.in0(alu),
		.in1(const_10_5_out),
		.out(magma_Bits_5_eq_inst19_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst2(
		.in0(alu),
		.in1(const_1_5_out),
		.out(magma_Bits_5_eq_inst2_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst20(
		.in0(alu),
		.in1(const_9_5_out),
		.out(magma_Bits_5_eq_inst20_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst21(
		.in0(alu),
		.in1(const_11_5_out),
		.out(magma_Bits_5_eq_inst21_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst22(
		.in0(alu),
		.in1(const_7_5_out),
		.out(magma_Bits_5_eq_inst22_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst23(
		.in0(alu),
		.in1(const_8_5_out),
		.out(magma_Bits_5_eq_inst23_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst24(
		.in0(alu),
		.in1(const_12_5_out),
		.out(magma_Bits_5_eq_inst24_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst25(
		.in0(alu),
		.in1(const_13_5_out),
		.out(magma_Bits_5_eq_inst25_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst26(
		.in0(alu),
		.in1(const_14_5_out),
		.out(magma_Bits_5_eq_inst26_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst27(
		.in0(alu),
		.in1(const_16_5_out),
		.out(magma_Bits_5_eq_inst27_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst28(
		.in0(alu),
		.in1(const_15_5_out),
		.out(magma_Bits_5_eq_inst28_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst29(
		.in0(alu),
		.in1(const_17_5_out),
		.out(magma_Bits_5_eq_inst29_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst3(
		.in0(alu),
		.in1(const_16_5_out),
		.out(magma_Bits_5_eq_inst3_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst30(
		.in0(alu),
		.in1(const_18_5_out),
		.out(magma_Bits_5_eq_inst30_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst4(
		.in0(alu),
		.in1(const_17_5_out),
		.out(magma_Bits_5_eq_inst4_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst5(
		.in0(alu),
		.in1(const_14_5_out),
		.out(magma_Bits_5_eq_inst5_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst6(
		.in0(alu),
		.in1(const_15_5_out),
		.out(magma_Bits_5_eq_inst6_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst7(
		.in0(alu),
		.in1(const_16_5_out),
		.out(magma_Bits_5_eq_inst7_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst8(
		.in0(alu),
		.in1(const_17_5_out),
		.out(magma_Bits_5_eq_inst8_out)
	);
	PEGEN_coreir_eq #(.width(5)) magma_Bits_5_eq_inst9(
		.in0(alu),
		.in1(const_13_5_out),
		.out(magma_Bits_5_eq_inst9_out)
	);
	PEGEN_coreir_ashr #(.width(16)) magma_SInt_16_ashr_inst0(
		.in0(Mux2xBits16_inst3_O),
		.in1(c),
		.out(magma_SInt_16_ashr_inst0_out)
	);
	PEGEN_coreir_eq #(.width(16)) magma_SInt_16_eq_inst0(
		.in0(const_0_16_out),
		.in1(Mux2xBits16_inst21_O),
		.out(magma_SInt_16_eq_inst0_out)
	);
	PEGEN_coreir_neg #(.width(16)) magma_SInt_16_neg_inst0(
		.in(a),
		.out(magma_SInt_16_neg_inst0_out)
	);
	PEGEN_coreir_sge #(.width(16)) magma_SInt_16_sge_inst0(
		.in0(Mux2xBits16_inst1_O),
		.in1(c),
		.out(magma_SInt_16_sge_inst0_out)
	);
	PEGEN_coreir_sle #(.width(16)) magma_SInt_16_sle_inst0(
		.in0(a),
		.in1(b),
		.out(magma_SInt_16_sle_inst0_out)
	);
	PEGEN_coreir_sle #(.width(16)) magma_SInt_16_sle_inst1(
		.in0(const_0_16_out),
		.in1(a),
		.out(magma_SInt_16_sle_inst1_out)
	);
	PEGEN_coreir_lshr #(.width(16)) magma_UInt_16_lshr_inst0(
		.in0(Mux2xBits16_inst3_O),
		.in1(c),
		.out(magma_UInt_16_lshr_inst0_out)
	);
	PEGEN_coreir_uge #(.width(16)) magma_UInt_16_uge_inst0(
		.in0(Mux2xBits16_inst1_O),
		.in1(c),
		.out(magma_UInt_16_uge_inst0_out)
	);
	PEGEN_coreir_ule #(.width(16)) magma_UInt_16_ule_inst0(
		.in0(a),
		.in1(b),
		.out(magma_UInt_16_ule_inst0_out)
	);
	wire [16:0] magma_UInt_17_add_inst0_in0;
	assign magma_UInt_17_add_inst0_in0 = {bit_const_0_None_out, a};
	wire [16:0] magma_UInt_17_add_inst0_in1;
	assign magma_UInt_17_add_inst0_in1 = {bit_const_0_None_out, Mux2xBits16_inst5_O};
	PEGEN_coreir_add #(.width(17)) magma_UInt_17_add_inst0(
		.in0(magma_UInt_17_add_inst0_in0),
		.in1(magma_UInt_17_add_inst0_in1),
		.out(magma_UInt_17_add_inst0_out)
	);
	wire [16:0] magma_UInt_17_add_inst1_in1;
	assign magma_UInt_17_add_inst1_in1 = {bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, d};
	PEGEN_coreir_add #(.width(17)) magma_UInt_17_add_inst1(
		.in0(magma_UInt_17_add_inst0_out),
		.in1(magma_UInt_17_add_inst1_in1),
		.out(magma_UInt_17_add_inst1_out)
	);
	wire [16:0] magma_UInt_17_add_inst2_in0;
	assign magma_UInt_17_add_inst2_in0 = {bit_const_0_None_out, Mux2xUInt16_inst0_O};
	wire [16:0] magma_UInt_17_add_inst2_in1;
	assign magma_UInt_17_add_inst2_in1 = {bit_const_0_None_out, Mux2xBits16_inst6_O};
	PEGEN_coreir_add #(.width(17)) magma_UInt_17_add_inst2(
		.in0(magma_UInt_17_add_inst2_in0),
		.in1(magma_UInt_17_add_inst2_in1),
		.out(magma_UInt_17_add_inst2_out)
	);
	wire [16:0] magma_UInt_17_add_inst3_in1;
	assign magma_UInt_17_add_inst3_in1 = {bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, Mux2xBit_inst2_O};
	PEGEN_coreir_add #(.width(17)) magma_UInt_17_add_inst3(
		.in0(magma_UInt_17_add_inst2_out),
		.in1(magma_UInt_17_add_inst3_in1),
		.out(magma_UInt_17_add_inst3_out)
	);
	PEGEN_coreir_mul #(.width(32)) magma_UInt_32_mul_inst0(
		.in0(Mux2xUInt32_inst0_O),
		.in1(Mux2xUInt32_inst1_O),
		.out(magma_UInt_32_mul_inst0_out)
	);
	assign res = Mux2xBits16_inst21_O;
	assign res_p = Mux2xBit_inst23_O;
	assign Z = magma_SInt_16_eq_inst0_out;
	assign N = Mux2xBits16_inst21_O[15];
	assign C = Mux2xBit_inst21_O;
	assign V = Mux2xBit_inst22_O;
endmodule
module PEGEN_PE (
	inst,
	data0,
	data1,
	data2,
	bit0,
	bit1,
	bit2,
	clk_en,
	O0,
	O1,
	O2,
	O3,
	O4,
	CLK,
	ASYNCRESET
);
	input [83:0] inst;
	input [15:0] data0;
	input [15:0] data1;
	input [15:0] data2;
	input bit0;
	input bit1;
	input bit2;
	input clk_en;
	output wire [15:0] O0;
	output wire O1;
	output wire [15:0] O2;
	output wire [15:0] O3;
	output wire [15:0] O4;
	input CLK;
	input ASYNCRESET;
	wire [15:0] ALU_inst0_res;
	wire ALU_inst0_res_p;
	wire ALU_inst0_Z;
	wire ALU_inst0_N;
	wire ALU_inst0_C;
	wire ALU_inst0_V;
	wire Cond_inst0_O;
	wire [15:0] FPCustom_inst0_res;
	wire FPCustom_inst0_res_p;
	wire FPCustom_inst0_V;
	wire [15:0] FPU_inst0_res;
	wire FPU_inst0_N;
	wire FPU_inst0_Z;
	wire LUT_inst0_O;
	wire Mux2xBit_inst0_O;
	wire Mux2xBit_inst1_O;
	wire Mux2xBit_inst2_O;
	wire Mux2xBit_inst3_O;
	wire Mux2xBit_inst4_O;
	wire Mux2xBit_inst5_O;
	wire Mux2xBit_inst6_O;
	wire Mux2xBit_inst7_O;
	wire [15:0] Mux2xBits16_inst0_O;
	wire [15:0] Mux2xBits16_inst1_O;
	wire [4:0] Mux2xMagmaADTALU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst0_O;
	wire [2:0] Mux2xMagmaADTFPCustom_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst0_O;
	wire [2:0] Mux2xMagmaADTFPCustom_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst1_O;
	wire [1:0] Mux2xMagmaADTFPU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst0_O;
	wire [1:0] Mux2xMagmaADTFPU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst1_O;
	wire [15:0] RegisterMode_inst0_O0;
	wire [15:0] RegisterMode_inst0_O1;
	wire [15:0] RegisterMode_inst1_O0;
	wire [15:0] RegisterMode_inst1_O1;
	wire [15:0] RegisterMode_inst2_O0;
	wire [15:0] RegisterMode_inst2_O1;
	wire RegisterMode_inst3_O0;
	wire RegisterMode_inst3_O1;
	wire RegisterMode_inst4_O0;
	wire RegisterMode_inst4_O1;
	wire RegisterMode_inst5_O0;
	wire RegisterMode_inst5_O1;
	wire bit_const_0_None_out;
	wire [1:0] const_0_2_out;
	wire [2:0] const_0_3_out;
	wire [4:0] const_0_5_out;
	wire [1:0] const_1_2_out;
	wire [1:0] const_2_2_out;
	wire magma_Bits_2_eq_inst0_out;
	wire magma_Bits_2_eq_inst1_out;
	wire magma_Bits_2_eq_inst2_out;
	wire magma_Bits_2_eq_inst3_out;
	wire magma_Bits_2_eq_inst4_out;
	wire magma_Bits_2_eq_inst5_out;
	wire magma_Bits_2_eq_inst6_out;
	PEGEN_ALU ALU_inst0(
		.alu(Mux2xMagmaADTALU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst0_O),
		.signed_(inst[7:7]),
		.a(RegisterMode_inst0_O0),
		.b(RegisterMode_inst1_O0),
		.c(RegisterMode_inst2_O0),
		.d(RegisterMode_inst3_O0),
		.res(ALU_inst0_res),
		.res_p(ALU_inst0_res_p),
		.Z(ALU_inst0_Z),
		.N(ALU_inst0_N),
		.C(ALU_inst0_C),
		.V(ALU_inst0_V),
		.CLK(CLK),
		.ASYNCRESET(ASYNCRESET)
	);
	PEGEN_Cond Cond_inst0(
		.code(inst[20:16]),
		.alu(Mux2xBit_inst7_O),
		.lut(LUT_inst0_O),
		.Z(Mux2xBit_inst6_O),
		.N(Mux2xBit_inst4_O),
		.C(ALU_inst0_C),
		.V(Mux2xBit_inst5_O),
		.O(Cond_inst0_O),
		.CLK(CLK),
		.ASYNCRESET(ASYNCRESET)
	);
	PEGEN_FPCustom FPCustom_inst0(
		.op(Mux2xMagmaADTFPCustom_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst1_O),
		.signed_(inst[7:7]),
		.a(RegisterMode_inst0_O0),
		.b(RegisterMode_inst1_O0),
		.res(FPCustom_inst0_res),
		.res_p(FPCustom_inst0_res_p),
		.V(FPCustom_inst0_V),
		.CLK(CLK),
		.ASYNCRESET(ASYNCRESET)
	);
	PEGEN_FPU FPU_inst0(
		.fpu_op(Mux2xMagmaADTFPU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst1_O),
		.a(RegisterMode_inst0_O0),
		.b(RegisterMode_inst1_O0),
		.res(FPU_inst0_res),
		.N(FPU_inst0_N),
		.Z(FPU_inst0_Z),
		.CLK(CLK),
		.ASYNCRESET(ASYNCRESET)
	);
	wire [7:0] LUT_inst0_lut;
	assign LUT_inst0_lut = {inst[15], inst[14], inst[13], inst[12], inst[11], inst[10], inst[9], inst[8]};
	PEGEN_LUT LUT_inst0(
		.lut(LUT_inst0_lut),
		.bit0(RegisterMode_inst3_O0),
		.bit1(RegisterMode_inst4_O0),
		.bit2(RegisterMode_inst5_O0),
		.O(LUT_inst0_O),
		.CLK(CLK),
		.ASYNCRESET(ASYNCRESET)
	);
	PEGEN_Mux2xBit Mux2xBit_inst0(
		.I0(bit_const_0_None_out),
		.I1(FPU_inst0_N),
		.S(magma_Bits_2_eq_inst6_out),
		.O(Mux2xBit_inst0_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst1(
		.I0(FPCustom_inst0_V),
		.I1(bit_const_0_None_out),
		.S(magma_Bits_2_eq_inst6_out),
		.O(Mux2xBit_inst1_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst2(
		.I0(bit_const_0_None_out),
		.I1(FPU_inst0_Z),
		.S(magma_Bits_2_eq_inst6_out),
		.O(Mux2xBit_inst2_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst3(
		.I0(FPCustom_inst0_res_p),
		.I1(bit_const_0_None_out),
		.S(magma_Bits_2_eq_inst6_out),
		.O(Mux2xBit_inst3_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst4(
		.I0(Mux2xBit_inst0_O),
		.I1(ALU_inst0_N),
		.S(magma_Bits_2_eq_inst5_out),
		.O(Mux2xBit_inst4_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst5(
		.I0(Mux2xBit_inst1_O),
		.I1(ALU_inst0_V),
		.S(magma_Bits_2_eq_inst5_out),
		.O(Mux2xBit_inst5_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst6(
		.I0(Mux2xBit_inst2_O),
		.I1(ALU_inst0_Z),
		.S(magma_Bits_2_eq_inst5_out),
		.O(Mux2xBit_inst6_O)
	);
	PEGEN_Mux2xBit Mux2xBit_inst7(
		.I0(Mux2xBit_inst3_O),
		.I1(ALU_inst0_res_p),
		.S(magma_Bits_2_eq_inst5_out),
		.O(Mux2xBit_inst7_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst0(
		.I0(FPCustom_inst0_res),
		.I1(FPU_inst0_res),
		.S(magma_Bits_2_eq_inst6_out),
		.O(Mux2xBits16_inst0_O)
	);
	PEGEN_Mux2xBits16 Mux2xBits16_inst1(
		.I0(Mux2xBits16_inst0_O),
		.I1(ALU_inst0_res),
		.S(magma_Bits_2_eq_inst5_out),
		.O(Mux2xBits16_inst1_O)
	);
	wire [4:0] Mux2xMagmaADTALU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst0_I1;
	assign Mux2xMagmaADTALU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst0_I1 = {inst[6], inst[5], inst[4], inst[3], inst[2]};
	PEGEN_Mux2xMagmaADTALU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3 Mux2xMagmaADTALU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst0(
		.I0(const_0_5_out),
		.I1(Mux2xMagmaADTALU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst0_I1),
		.S(magma_Bits_2_eq_inst0_out),
		.O(Mux2xMagmaADTALU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst0_O)
	);
	wire [2:0] Mux2xMagmaADTFPCustom_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst0_I0;
	assign Mux2xMagmaADTFPCustom_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst0_I0 = {inst[4], inst[3], inst[2]};
	PEGEN_Mux2xMagmaADTFPCustom_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3 Mux2xMagmaADTFPCustom_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst0(
		.I0(Mux2xMagmaADTFPCustom_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst0_I0),
		.I1(const_0_3_out),
		.S(magma_Bits_2_eq_inst2_out),
		.O(Mux2xMagmaADTFPCustom_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst0_O)
	);
	PEGEN_Mux2xMagmaADTFPCustom_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3 Mux2xMagmaADTFPCustom_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst1(
		.I0(Mux2xMagmaADTFPCustom_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst0_O),
		.I1(const_0_3_out),
		.S(magma_Bits_2_eq_inst0_out),
		.O(Mux2xMagmaADTFPCustom_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst1_O)
	);
	wire [1:0] Mux2xMagmaADTFPU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst0_I1;
	assign Mux2xMagmaADTFPU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst0_I1 = {inst[3], inst[2]};
	PEGEN_Mux2xMagmaADTFPU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3 Mux2xMagmaADTFPU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst0(
		.I0(const_0_2_out),
		.I1(Mux2xMagmaADTFPU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst0_I1),
		.S(magma_Bits_2_eq_inst2_out),
		.O(Mux2xMagmaADTFPU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst0_O)
	);
	PEGEN_Mux2xMagmaADTFPU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3 Mux2xMagmaADTFPU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst1(
		.I0(Mux2xMagmaADTFPU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst0_O),
		.I1(const_0_2_out),
		.S(magma_Bits_2_eq_inst0_out),
		.O(Mux2xMagmaADTFPU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst1_O)
	);
	wire [15:0] RegisterMode_inst0_const_;
	assign RegisterMode_inst0_const_ = {inst[38], inst[37], inst[36], inst[35], inst[34], inst[33], inst[32], inst[31], inst[30], inst[29], inst[28], inst[27], inst[26], inst[25], inst[24], inst[23]};
	PEGEN_RegisterMode RegisterMode_inst0(
		.mode(inst[22:21]),
		.const_(RegisterMode_inst0_const_),
		.value(data0),
		.clk_en(clk_en),
		.O0(RegisterMode_inst0_O0),
		.O1(RegisterMode_inst0_O1),
		.CLK(CLK),
		.ASYNCRESET(ASYNCRESET)
	);
	wire [15:0] RegisterMode_inst1_const_;
	assign RegisterMode_inst1_const_ = {inst[56], inst[55], inst[54], inst[53], inst[52], inst[51], inst[50], inst[49], inst[48], inst[47], inst[46], inst[45], inst[44], inst[43], inst[42], inst[41]};
	PEGEN_RegisterMode RegisterMode_inst1(
		.mode(inst[40:39]),
		.const_(RegisterMode_inst1_const_),
		.value(data1),
		.clk_en(clk_en),
		.O0(RegisterMode_inst1_O0),
		.O1(RegisterMode_inst1_O1),
		.CLK(CLK),
		.ASYNCRESET(ASYNCRESET)
	);
	wire [15:0] RegisterMode_inst2_const_;
	assign RegisterMode_inst2_const_ = {inst[74], inst[73], inst[72], inst[71], inst[70], inst[69], inst[68], inst[67], inst[66], inst[65], inst[64], inst[63], inst[62], inst[61], inst[60], inst[59]};
	PEGEN_RegisterMode RegisterMode_inst2(
		.mode(inst[58:57]),
		.const_(RegisterMode_inst2_const_),
		.value(data2),
		.clk_en(clk_en),
		.O0(RegisterMode_inst2_O0),
		.O1(RegisterMode_inst2_O1),
		.CLK(CLK),
		.ASYNCRESET(ASYNCRESET)
	);
	PEGEN_RegisterMode_unq1 RegisterMode_inst3(
		.mode(inst[76:75]),
		.const_(inst[77]),
		.value(bit0),
		.clk_en(clk_en),
		.O0(RegisterMode_inst3_O0),
		.O1(RegisterMode_inst3_O1),
		.CLK(CLK),
		.ASYNCRESET(ASYNCRESET)
	);
	PEGEN_RegisterMode_unq1 RegisterMode_inst4(
		.mode(inst[79:78]),
		.const_(inst[80]),
		.value(bit1),
		.clk_en(clk_en),
		.O0(RegisterMode_inst4_O0),
		.O1(RegisterMode_inst4_O1),
		.CLK(CLK),
		.ASYNCRESET(ASYNCRESET)
	);
	PEGEN_RegisterMode_unq1 RegisterMode_inst5(
		.mode(inst[82:81]),
		.const_(inst[83]),
		.value(bit2),
		.clk_en(clk_en),
		.O0(RegisterMode_inst5_O0),
		.O1(RegisterMode_inst5_O1),
		.CLK(CLK),
		.ASYNCRESET(ASYNCRESET)
	);
	PEGEN_corebit_const #(.value(1'b0)) bit_const_0_None(.out(bit_const_0_None_out));
	PEGEN_coreir_const #(
		.value(2'h0),
		.width(2)
	) const_0_2(.out(const_0_2_out));
	PEGEN_coreir_const #(
		.value(3'h0),
		.width(3)
	) const_0_3(.out(const_0_3_out));
	PEGEN_coreir_const #(
		.value(5'h00),
		.width(5)
	) const_0_5(.out(const_0_5_out));
	PEGEN_coreir_const #(
		.value(2'h1),
		.width(2)
	) const_1_2(.out(const_1_2_out));
	PEGEN_coreir_const #(
		.value(2'h2),
		.width(2)
	) const_2_2(.out(const_2_2_out));
	wire [1:0] magma_Bits_2_eq_inst0_in0;
	assign magma_Bits_2_eq_inst0_in0 = {inst[1], inst[0]};
	PEGEN_coreir_eq #(.width(2)) magma_Bits_2_eq_inst0(
		.in0(magma_Bits_2_eq_inst0_in0),
		.in1(const_0_2_out),
		.out(magma_Bits_2_eq_inst0_out)
	);
	wire [1:0] magma_Bits_2_eq_inst1_in0;
	assign magma_Bits_2_eq_inst1_in0 = {inst[1], inst[0]};
	PEGEN_coreir_eq #(.width(2)) magma_Bits_2_eq_inst1(
		.in0(magma_Bits_2_eq_inst1_in0),
		.in1(const_0_2_out),
		.out(magma_Bits_2_eq_inst1_out)
	);
	wire [1:0] magma_Bits_2_eq_inst2_in0;
	assign magma_Bits_2_eq_inst2_in0 = {inst[1], inst[0]};
	PEGEN_coreir_eq #(.width(2)) magma_Bits_2_eq_inst2(
		.in0(magma_Bits_2_eq_inst2_in0),
		.in1(const_2_2_out),
		.out(magma_Bits_2_eq_inst2_out)
	);
	wire [1:0] magma_Bits_2_eq_inst3_in0;
	assign magma_Bits_2_eq_inst3_in0 = {inst[1], inst[0]};
	PEGEN_coreir_eq #(.width(2)) magma_Bits_2_eq_inst3(
		.in0(magma_Bits_2_eq_inst3_in0),
		.in1(const_2_2_out),
		.out(magma_Bits_2_eq_inst3_out)
	);
	wire [1:0] magma_Bits_2_eq_inst4_in0;
	assign magma_Bits_2_eq_inst4_in0 = {inst[1], inst[0]};
	PEGEN_coreir_eq #(.width(2)) magma_Bits_2_eq_inst4(
		.in0(magma_Bits_2_eq_inst4_in0),
		.in1(const_1_2_out),
		.out(magma_Bits_2_eq_inst4_out)
	);
	wire [1:0] magma_Bits_2_eq_inst5_in0;
	assign magma_Bits_2_eq_inst5_in0 = {inst[1], inst[0]};
	PEGEN_coreir_eq #(.width(2)) magma_Bits_2_eq_inst5(
		.in0(magma_Bits_2_eq_inst5_in0),
		.in1(const_0_2_out),
		.out(magma_Bits_2_eq_inst5_out)
	);
	wire [1:0] magma_Bits_2_eq_inst6_in0;
	assign magma_Bits_2_eq_inst6_in0 = {inst[1], inst[0]};
	PEGEN_coreir_eq #(.width(2)) magma_Bits_2_eq_inst6(
		.in0(magma_Bits_2_eq_inst6_in0),
		.in1(const_2_2_out),
		.out(magma_Bits_2_eq_inst6_out)
	);
	assign O0 = Mux2xBits16_inst1_O;
	assign O1 = Cond_inst0_O;
	assign O2 = RegisterMode_inst0_O1;
	assign O3 = RegisterMode_inst1_O1;
	assign O4 = RegisterMode_inst2_O1;
endmodule
